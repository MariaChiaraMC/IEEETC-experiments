module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 ;
  output y0 ;
  wire n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 ;
  assign n23 = x1 ^ x0 ;
  assign n24 = x2 ^ x1 ;
  assign n25 = n24 ^ x2 ;
  assign n26 = x3 ^ x2 ;
  assign n27 = ~n25 & ~n26 ;
  assign n28 = n27 ^ x2 ;
  assign n29 = n23 & ~n28 ;
  assign n30 = x5 ^ x3 ;
  assign n31 = ~x4 & ~n30 ;
  assign n32 = n29 & n31 ;
  assign n237 = ~x19 & ~x20 ;
  assign n33 = x0 & ~x1 ;
  assign n34 = ~x21 & n33 ;
  assign n35 = ~x2 & n34 ;
  assign n59 = x9 & x10 ;
  assign n60 = x11 & ~x12 ;
  assign n61 = ~x2 & x4 ;
  assign n62 = n60 & n61 ;
  assign n63 = n59 & n62 ;
  assign n64 = x0 & ~x4 ;
  assign n65 = x0 & ~x13 ;
  assign n66 = n61 & ~n65 ;
  assign n67 = ~n64 & ~n66 ;
  assign n68 = x1 & ~n67 ;
  assign n69 = ~n63 & ~n68 ;
  assign n36 = ~x6 & ~x13 ;
  assign n37 = ~x4 & ~x12 ;
  assign n38 = ~x7 & n37 ;
  assign n39 = n36 & n38 ;
  assign n40 = x11 ^ x10 ;
  assign n41 = ~x8 & n40 ;
  assign n42 = ~x0 & ~x11 ;
  assign n43 = n42 ^ x2 ;
  assign n44 = x9 ^ x2 ;
  assign n45 = n44 ^ x2 ;
  assign n46 = n45 ^ n41 ;
  assign n47 = ~n43 & n46 ;
  assign n48 = n47 ^ n42 ;
  assign n49 = n41 & n48 ;
  assign n50 = n39 & n49 ;
  assign n51 = ~x2 & ~n24 ;
  assign n52 = x0 & n51 ;
  assign n53 = n52 ^ n24 ;
  assign n54 = ~n50 & n53 ;
  assign n70 = n69 ^ n54 ;
  assign n71 = n70 ^ n54 ;
  assign n55 = x2 & ~x4 ;
  assign n56 = ~x0 & n55 ;
  assign n57 = n56 ^ n54 ;
  assign n58 = n57 ^ n54 ;
  assign n72 = n71 ^ n58 ;
  assign n73 = ~x12 & x13 ;
  assign n74 = ~x2 & n73 ;
  assign n75 = ~x0 & ~n74 ;
  assign n76 = n75 ^ x4 ;
  assign n77 = n76 ^ x1 ;
  assign n78 = ~x8 & x9 ;
  assign n79 = ~x10 & x13 ;
  assign n80 = n79 ^ x12 ;
  assign n81 = ~x11 & ~n80 ;
  assign n82 = n81 ^ x12 ;
  assign n83 = n78 & ~n82 ;
  assign n84 = x7 & x11 ;
  assign n85 = n73 & n84 ;
  assign n86 = x8 & x10 ;
  assign n87 = n60 & n86 ;
  assign n88 = x12 & ~x16 ;
  assign n89 = x7 & ~n88 ;
  assign n90 = ~n87 & n89 ;
  assign n91 = ~x6 & ~n90 ;
  assign n92 = x10 ^ x8 ;
  assign n93 = n92 ^ x16 ;
  assign n94 = n93 ^ x16 ;
  assign n95 = n94 ^ x10 ;
  assign n96 = x15 ^ x10 ;
  assign n97 = n40 & n96 ;
  assign n98 = x16 ^ x10 ;
  assign n99 = ~n94 & n98 ;
  assign n100 = n99 ^ n95 ;
  assign n101 = n97 & ~n100 ;
  assign n102 = n101 ^ n99 ;
  assign n103 = ~n95 & n102 ;
  assign n104 = n103 ^ n99 ;
  assign n105 = n104 ^ n92 ;
  assign n106 = n105 ^ x12 ;
  assign n107 = n106 ^ n105 ;
  assign n108 = n107 ^ x7 ;
  assign n109 = x16 ^ x13 ;
  assign n110 = x16 & ~n109 ;
  assign n111 = n110 ^ n105 ;
  assign n112 = n111 ^ x16 ;
  assign n113 = ~n108 & n112 ;
  assign n114 = n113 ^ n110 ;
  assign n115 = n114 ^ x16 ;
  assign n116 = ~x7 & n115 ;
  assign n117 = n116 ^ x7 ;
  assign n118 = n91 & n117 ;
  assign n119 = x12 & ~x13 ;
  assign n120 = ~x8 & ~x15 ;
  assign n121 = ~x13 & ~n59 ;
  assign n122 = ~n120 & ~n121 ;
  assign n123 = x13 ^ x6 ;
  assign n124 = n123 ^ n122 ;
  assign n126 = x11 & ~x16 ;
  assign n127 = x12 ^ x10 ;
  assign n128 = x12 ^ x11 ;
  assign n129 = x12 ^ x9 ;
  assign n130 = x12 & ~n129 ;
  assign n131 = n130 ^ x12 ;
  assign n132 = ~n128 & n131 ;
  assign n133 = n132 ^ n130 ;
  assign n134 = n133 ^ x12 ;
  assign n135 = n134 ^ x9 ;
  assign n136 = n127 & ~n135 ;
  assign n137 = n136 ^ x12 ;
  assign n138 = ~n126 & ~n137 ;
  assign n125 = x9 & n84 ;
  assign n139 = n138 ^ n125 ;
  assign n140 = ~x13 & n139 ;
  assign n141 = n140 ^ n138 ;
  assign n142 = ~n124 & n141 ;
  assign n143 = n142 ^ n140 ;
  assign n144 = n143 ^ n138 ;
  assign n145 = n144 ^ x13 ;
  assign n146 = ~n122 & ~n145 ;
  assign n147 = ~n119 & ~n146 ;
  assign n148 = ~x17 & ~n147 ;
  assign n149 = ~n118 & n148 ;
  assign n150 = x2 & ~n149 ;
  assign n151 = ~n85 & ~n150 ;
  assign n152 = ~n83 & n151 ;
  assign n153 = n152 ^ x2 ;
  assign n154 = x4 & ~n153 ;
  assign n155 = n154 ^ x2 ;
  assign n156 = n77 & ~n155 ;
  assign n157 = n156 ^ n154 ;
  assign n158 = n157 ^ x2 ;
  assign n159 = n158 ^ x4 ;
  assign n160 = ~x1 & ~n159 ;
  assign n161 = n160 ^ n54 ;
  assign n162 = n161 ^ n54 ;
  assign n163 = n162 ^ n71 ;
  assign n164 = n71 & ~n163 ;
  assign n165 = n164 ^ n71 ;
  assign n166 = ~n72 & n165 ;
  assign n167 = n166 ^ n164 ;
  assign n168 = n167 ^ n54 ;
  assign n169 = n168 ^ n71 ;
  assign n170 = ~x3 & n169 ;
  assign n171 = n170 ^ n54 ;
  assign n172 = ~n35 & n171 ;
  assign n173 = x5 & ~n172 ;
  assign n174 = x4 ^ x0 ;
  assign n175 = ~x1 & ~x2 ;
  assign n176 = n175 ^ n174 ;
  assign n177 = x3 ^ x0 ;
  assign n178 = n177 ^ x3 ;
  assign n179 = n30 & n178 ;
  assign n180 = n179 ^ x3 ;
  assign n181 = n180 ^ n174 ;
  assign n182 = ~n176 & n181 ;
  assign n183 = n182 ^ n179 ;
  assign n184 = n183 ^ x3 ;
  assign n185 = n184 ^ n175 ;
  assign n186 = ~n174 & ~n185 ;
  assign n187 = n186 ^ n174 ;
  assign n193 = x3 & x4 ;
  assign n190 = x0 & ~x5 ;
  assign n191 = ~x1 & n190 ;
  assign n188 = ~x0 & x1 ;
  assign n189 = ~x5 & n188 ;
  assign n192 = n191 ^ n189 ;
  assign n194 = n193 ^ n192 ;
  assign n195 = n194 ^ n189 ;
  assign n205 = n195 ^ n192 ;
  assign n206 = n205 ^ n189 ;
  assign n207 = n206 ^ n189 ;
  assign n196 = ~x3 & n39 ;
  assign n208 = ~x10 & x11 ;
  assign n197 = x10 & ~x11 ;
  assign n209 = n208 ^ n197 ;
  assign n210 = n209 ^ n197 ;
  assign n211 = n197 ^ x9 ;
  assign n212 = n211 ^ n197 ;
  assign n213 = n210 & n212 ;
  assign n214 = n213 ^ n197 ;
  assign n215 = x8 & n214 ;
  assign n216 = n215 ^ n197 ;
  assign n217 = n196 & n216 ;
  assign n218 = n217 ^ n192 ;
  assign n219 = n218 ^ n192 ;
  assign n220 = n219 ^ n189 ;
  assign n221 = n207 & n220 ;
  assign n198 = n78 & n197 ;
  assign n199 = x2 & n198 ;
  assign n200 = n196 & n199 ;
  assign n201 = n200 ^ n192 ;
  assign n202 = n201 ^ n195 ;
  assign n203 = n202 ^ n189 ;
  assign n204 = n195 & n203 ;
  assign n222 = n221 ^ n204 ;
  assign n223 = n222 ^ n195 ;
  assign n224 = n204 ^ n189 ;
  assign n225 = n224 ^ n206 ;
  assign n226 = ~n189 & n225 ;
  assign n227 = n226 ^ n204 ;
  assign n228 = n223 & n227 ;
  assign n229 = n228 ^ n221 ;
  assign n230 = n229 ^ n226 ;
  assign n231 = n230 ^ n195 ;
  assign n232 = n231 ^ n189 ;
  assign n233 = n232 ^ n206 ;
  assign n234 = n233 ^ n191 ;
  assign n235 = n187 & ~n234 ;
  assign n236 = ~n173 & n235 ;
  assign n238 = n237 ^ n236 ;
  assign n239 = n238 ^ n236 ;
  assign n240 = n236 ^ x18 ;
  assign n241 = ~n239 & n240 ;
  assign n242 = n241 ^ n236 ;
  assign n243 = ~n32 & n242 ;
  assign n244 = x14 & ~n243 ;
  assign y0 = n244 ;
endmodule
