module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 ;
  assign n18 = x1 & ~x7 ;
  assign n19 = x5 & ~x6 ;
  assign n20 = n18 & n19 ;
  assign n21 = x3 & ~n20 ;
  assign n22 = ~x2 & ~n21 ;
  assign n17 = x3 ^ x0 ;
  assign n23 = n22 ^ n17 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ x0 ;
  assign n26 = n22 ^ x0 ;
  assign n27 = ~n25 & ~n26 ;
  assign n28 = n27 ^ n22 ;
  assign n29 = n25 ^ n22 ;
  assign n39 = ~x9 & ~x10 ;
  assign n40 = ~x14 & ~x15 ;
  assign n41 = x13 & ~n40 ;
  assign n42 = ~x8 & ~x12 ;
  assign n43 = x15 ^ x14 ;
  assign n44 = ~x13 & ~n43 ;
  assign n45 = n42 & ~n44 ;
  assign n46 = ~n41 & n45 ;
  assign n168 = ~x11 & n18 ;
  assign n169 = n46 & n168 ;
  assign n170 = ~n39 & n169 ;
  assign n36 = x6 & ~x11 ;
  assign n37 = x9 & x10 ;
  assign n38 = n36 & ~n37 ;
  assign n47 = ~n39 & n46 ;
  assign n48 = n38 & n47 ;
  assign n35 = x5 ^ x1 ;
  assign n49 = n48 ^ n35 ;
  assign n50 = n35 ^ x1 ;
  assign n51 = n49 & n50 ;
  assign n52 = n51 ^ n35 ;
  assign n59 = ~x8 & ~n37 ;
  assign n57 = ~x12 & x14 ;
  assign n53 = x12 & ~x14 ;
  assign n54 = x10 & ~x15 ;
  assign n55 = ~x9 & ~n54 ;
  assign n56 = n53 & ~n55 ;
  assign n58 = n57 ^ n56 ;
  assign n60 = n59 ^ n58 ;
  assign n70 = n60 ^ n58 ;
  assign n61 = ~x10 & x15 ;
  assign n62 = ~x8 & x9 ;
  assign n63 = n61 & n62 ;
  assign n64 = n63 ^ n60 ;
  assign n65 = n64 ^ n58 ;
  assign n66 = n60 ^ n56 ;
  assign n67 = n66 ^ n63 ;
  assign n68 = n67 ^ n65 ;
  assign n69 = ~n65 & ~n68 ;
  assign n71 = n70 ^ n69 ;
  assign n72 = n71 ^ n65 ;
  assign n73 = n58 ^ x15 ;
  assign n74 = n69 ^ n65 ;
  assign n75 = n73 & ~n74 ;
  assign n76 = n75 ^ n58 ;
  assign n77 = ~n72 & n76 ;
  assign n78 = n77 ^ n58 ;
  assign n79 = n78 ^ n57 ;
  assign n80 = n79 ^ n58 ;
  assign n81 = n36 & n80 ;
  assign n82 = ~x12 & ~x15 ;
  assign n83 = x14 & ~x15 ;
  assign n84 = ~x13 & ~n83 ;
  assign n85 = x11 & x14 ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = n82 & ~n86 ;
  assign n88 = x12 & x14 ;
  assign n89 = n38 & ~n88 ;
  assign n90 = n89 ^ x6 ;
  assign n91 = n90 ^ x6 ;
  assign n92 = x8 ^ x6 ;
  assign n93 = n92 ^ x6 ;
  assign n94 = n91 & ~n93 ;
  assign n95 = n94 ^ x6 ;
  assign n96 = n84 & n95 ;
  assign n97 = n96 ^ x6 ;
  assign n98 = ~n87 & n97 ;
  assign n99 = ~n81 & n98 ;
  assign n100 = ~x11 & n55 ;
  assign n101 = ~x8 & n100 ;
  assign n102 = ~n88 & ~n101 ;
  assign n103 = x14 ^ x12 ;
  assign n104 = n61 ^ x15 ;
  assign n105 = n43 ^ x15 ;
  assign n106 = ~n104 & ~n105 ;
  assign n107 = n106 ^ x15 ;
  assign n108 = ~n103 & n107 ;
  assign n109 = ~x13 & ~n108 ;
  assign n110 = x6 & n109 ;
  assign n111 = ~n102 & n110 ;
  assign n112 = ~x10 & ~x11 ;
  assign n113 = n41 & ~n82 ;
  assign n114 = ~n112 & n113 ;
  assign n115 = ~n111 & ~n114 ;
  assign n116 = ~n53 & ~n57 ;
  assign n117 = x15 & n116 ;
  assign n118 = n40 ^ x11 ;
  assign n119 = n118 ^ n40 ;
  assign n120 = x14 ^ x8 ;
  assign n121 = n120 ^ x14 ;
  assign n122 = n121 ^ x10 ;
  assign n123 = n122 ^ x14 ;
  assign n124 = n123 ^ n122 ;
  assign n128 = n122 ^ x12 ;
  assign n129 = n122 & ~n128 ;
  assign n125 = x10 ^ x9 ;
  assign n126 = ~n121 & ~n125 ;
  assign n132 = n129 ^ n126 ;
  assign n127 = n126 ^ n124 ;
  assign n130 = n129 ^ n122 ;
  assign n131 = ~n127 & n130 ;
  assign n133 = n132 ^ n131 ;
  assign n134 = ~n124 & n133 ;
  assign n135 = n134 ^ n129 ;
  assign n136 = n135 ^ n131 ;
  assign n137 = n136 ^ n120 ;
  assign n140 = n137 ^ x10 ;
  assign n141 = n140 ^ n137 ;
  assign n138 = n137 ^ n62 ;
  assign n139 = n138 ^ n137 ;
  assign n142 = n141 ^ n139 ;
  assign n143 = n137 ^ n116 ;
  assign n144 = n143 ^ n137 ;
  assign n145 = n144 ^ n141 ;
  assign n146 = ~n141 & n145 ;
  assign n147 = n146 ^ n141 ;
  assign n148 = n142 & ~n147 ;
  assign n149 = n148 ^ n146 ;
  assign n150 = n149 ^ n137 ;
  assign n151 = n150 ^ n141 ;
  assign n152 = x15 & ~n151 ;
  assign n153 = n152 ^ n137 ;
  assign n154 = n153 ^ n40 ;
  assign n155 = ~n119 & n154 ;
  assign n156 = n155 ^ n40 ;
  assign n157 = ~n117 & ~n156 ;
  assign n158 = x13 & ~n157 ;
  assign n159 = n115 & ~n158 ;
  assign n160 = n99 & n159 ;
  assign n161 = n35 & ~n160 ;
  assign n162 = n161 ^ x7 ;
  assign n163 = n52 & n162 ;
  assign n164 = n163 ^ n161 ;
  assign n165 = x7 & n164 ;
  assign n166 = n165 ^ x7 ;
  assign n167 = n166 ^ x7 ;
  assign n171 = n170 ^ n167 ;
  assign n172 = n167 ^ n22 ;
  assign n173 = n171 & ~n172 ;
  assign n30 = n22 ^ x1 ;
  assign n31 = n30 ^ n22 ;
  assign n32 = n31 ^ n22 ;
  assign n33 = n32 ^ n25 ;
  assign n34 = ~n25 & n33 ;
  assign n174 = n173 ^ n34 ;
  assign n175 = n174 ^ n31 ;
  assign n176 = n175 ^ n170 ;
  assign n177 = n176 ^ n22 ;
  assign n178 = n177 ^ n25 ;
  assign n179 = n29 & n178 ;
  assign n180 = n179 ^ n34 ;
  assign n181 = n180 ^ n22 ;
  assign n182 = n181 ^ x0 ;
  assign n183 = ~n28 & ~n182 ;
  assign n184 = n183 ^ n179 ;
  assign n185 = n184 ^ x0 ;
  assign n186 = n185 ^ n25 ;
  assign n187 = n186 ^ n22 ;
  assign n188 = n187 ^ n22 ;
  assign n189 = x4 & n188 ;
  assign y0 = n189 ;
endmodule
