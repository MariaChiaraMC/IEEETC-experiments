module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 ;
  assign n9 = x5 & x6 ;
  assign n10 = x3 & n9 ;
  assign n11 = ~x2 & ~n10 ;
  assign n12 = ~x5 & ~x6 ;
  assign n13 = ~x7 & n12 ;
  assign n14 = ~x3 & ~n9 ;
  assign n15 = ~n13 & n14 ;
  assign n16 = n11 & ~n15 ;
  assign n17 = x7 & n9 ;
  assign n18 = x3 & ~n17 ;
  assign n19 = x2 & ~n18 ;
  assign n20 = ~x1 & n19 ;
  assign n21 = ~n16 & ~n20 ;
  assign n22 = ~x4 & ~n21 ;
  assign n23 = x4 ^ x2 ;
  assign n24 = n23 ^ x2 ;
  assign n25 = n24 ^ x1 ;
  assign n26 = n12 ^ n9 ;
  assign n27 = n24 ^ x3 ;
  assign n28 = ~n26 & n27 ;
  assign n29 = n28 ^ n12 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n30 ^ x2 ;
  assign n32 = ~x2 & n31 ;
  assign n33 = n32 ^ x3 ;
  assign n34 = n33 ^ x2 ;
  assign n35 = n34 ^ n24 ;
  assign n36 = n35 ^ x1 ;
  assign n37 = ~n25 & n36 ;
  assign n38 = n37 ^ n32 ;
  assign n39 = n38 ^ x3 ;
  assign n40 = n39 ^ n24 ;
  assign n41 = ~x1 & n40 ;
  assign n42 = n41 ^ x1 ;
  assign n43 = n42 ^ x2 ;
  assign n44 = ~n22 & ~n43 ;
  assign y0 = ~n44 ;
endmodule
