module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 ;
  assign n15 = x11 ^ x8 ;
  assign n16 = x9 & ~x12 ;
  assign n17 = x13 ^ x10 ;
  assign n18 = x13 ^ x1 ;
  assign n19 = n18 ^ x1 ;
  assign n20 = x1 ^ x0 ;
  assign n21 = ~n19 & n20 ;
  assign n22 = n21 ^ x1 ;
  assign n23 = n17 & n22 ;
  assign n24 = n16 & n23 ;
  assign n25 = ~x9 & x12 ;
  assign n26 = ~x10 & x13 ;
  assign n27 = x3 & n26 ;
  assign n28 = x10 & ~x13 ;
  assign n29 = x2 & n28 ;
  assign n30 = ~n27 & ~n29 ;
  assign n31 = n25 & ~n30 ;
  assign n32 = ~n24 & ~n31 ;
  assign n33 = n32 ^ x11 ;
  assign n34 = n33 ^ n32 ;
  assign n35 = x12 ^ x9 ;
  assign n36 = x5 & n26 ;
  assign n37 = x4 & n28 ;
  assign n38 = ~n36 & ~n37 ;
  assign n39 = n38 ^ x12 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = x7 & n26 ;
  assign n42 = x6 & n28 ;
  assign n43 = ~n41 & ~n42 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = n40 & n44 ;
  assign n46 = n45 ^ n38 ;
  assign n47 = n35 & ~n46 ;
  assign n48 = n47 ^ n32 ;
  assign n49 = n34 & ~n48 ;
  assign n50 = n49 ^ n32 ;
  assign n51 = n15 & ~n50 ;
  assign y0 = n51 ;
endmodule
