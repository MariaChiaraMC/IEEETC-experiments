module top( x0 , x1 , x2 , x3 , x4 , y0 );
  input x0 , x1 , x2 , x3 , x4 ;
  output y0 ;
  wire n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 ;
  assign n6 = x3 ^ x2 ;
  assign n7 = n6 ^ x4 ;
  assign n8 = x4 ^ x1 ;
  assign n9 = n8 ^ x4 ;
  assign n10 = x4 ^ x3 ;
  assign n11 = n10 ^ x4 ;
  assign n12 = ~n9 & ~n11 ;
  assign n13 = n12 ^ x4 ;
  assign n14 = x0 & x4 ;
  assign n15 = n14 ^ n7 ;
  assign n16 = n13 & n15 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = n7 & n17 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = n19 ^ n7 ;
  assign y0 = n20 ;
endmodule
