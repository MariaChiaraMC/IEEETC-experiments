module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n16 = ~x1 & x8 ;
  assign n17 = x7 & x13 ;
  assign n18 = x4 & n17 ;
  assign n19 = n16 & n18 ;
  assign n20 = x6 & x11 ;
  assign n21 = ~x2 & n20 ;
  assign n22 = ~x5 & n21 ;
  assign n23 = n19 & n22 ;
  assign n24 = x0 & x12 ;
  assign n25 = x10 & x14 ;
  assign n26 = x9 & n25 ;
  assign n27 = n24 & n26 ;
  assign n28 = x3 & n27 ;
  assign n29 = n23 & n28 ;
  assign y0 = n29 ;
endmodule
