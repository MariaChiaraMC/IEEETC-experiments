module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n18 = x8 & x9 ;
  assign n19 = x0 & ~x6 ;
  assign n20 = n18 & n19 ;
  assign n21 = ~x1 & ~x3 ;
  assign n22 = ~x4 & n21 ;
  assign n23 = n20 & n22 ;
  assign n24 = ~x10 & x14 ;
  assign n25 = n23 & n24 ;
  assign n26 = x5 & ~x12 ;
  assign n27 = x11 & x15 ;
  assign n28 = x13 & n27 ;
  assign n29 = ~x2 & x7 ;
  assign n30 = x16 & ~n29 ;
  assign n31 = n28 & n30 ;
  assign n32 = n26 & n31 ;
  assign n33 = n25 & n32 ;
  assign y0 = n33 ;
endmodule
