module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 ;
  assign n17 = ~x0 & ~x2 ;
  assign n43 = x1 & ~x7 ;
  assign n19 = x4 & x5 ;
  assign n44 = x3 & n19 ;
  assign n45 = n43 & n44 ;
  assign n46 = n45 ^ x6 ;
  assign n18 = x7 ^ x1 ;
  assign n20 = n19 ^ x7 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = ~x8 & x9 ;
  assign n24 = x15 ^ x13 ;
  assign n25 = x14 & ~x15 ;
  assign n26 = ~n24 & n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n23 & n27 ;
  assign n29 = ~x13 & ~x15 ;
  assign n30 = x14 & ~n29 ;
  assign n31 = ~x11 & ~x12 ;
  assign n32 = x10 & n31 ;
  assign n33 = ~n30 & n32 ;
  assign n34 = n33 ^ n28 ;
  assign n35 = n28 & n34 ;
  assign n36 = n35 ^ n19 ;
  assign n37 = n36 ^ n28 ;
  assign n38 = ~n22 & n37 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n39 ^ n28 ;
  assign n41 = n18 & n40 ;
  assign n42 = n41 ^ x6 ;
  assign n47 = n46 ^ n42 ;
  assign n48 = n47 ^ x3 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = n47 ^ n46 ;
  assign n51 = n50 ^ x6 ;
  assign n52 = ~n49 & n51 ;
  assign n53 = n52 ^ n46 ;
  assign n54 = ~x4 & x5 ;
  assign n55 = ~n46 & ~n54 ;
  assign n56 = n55 ^ x6 ;
  assign n57 = ~n53 & ~n56 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = ~x6 & n58 ;
  assign n60 = n59 ^ n52 ;
  assign n61 = n60 ^ n45 ;
  assign n62 = n61 ^ n46 ;
  assign n63 = n17 & ~n62 ;
  assign y0 = n63 ;
endmodule
