// Benchmark "./pla/sqr6.pla_res_11NonExact" written by ABC on Fri Nov 20 10:29:18 2020

module \./pla/sqr6.pla_res_11NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = x0;
endmodule


