module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 ;
  assign n17 = ~x3 & ~x4 ;
  assign n18 = x1 ^ x0 ;
  assign n19 = ~x11 & ~x12 ;
  assign n20 = ~x9 & ~x10 ;
  assign n21 = ~x8 & n20 ;
  assign n22 = n19 & ~n21 ;
  assign n23 = x14 ^ x13 ;
  assign n24 = n23 ^ x15 ;
  assign n25 = n24 ^ x8 ;
  assign n32 = n25 ^ n24 ;
  assign n26 = n25 ^ x14 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n25 ^ x15 ;
  assign n29 = n28 ^ x14 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n27 & n30 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = x9 & x10 ;
  assign n36 = ~x15 & ~n35 ;
  assign n37 = n36 ^ n24 ;
  assign n38 = n31 ^ n27 ;
  assign n39 = n37 & n38 ;
  assign n40 = n39 ^ n24 ;
  assign n41 = ~n34 & n40 ;
  assign n42 = n41 ^ n24 ;
  assign n43 = n42 ^ n24 ;
  assign n44 = n22 & n43 ;
  assign n45 = ~x7 & ~n44 ;
  assign n46 = ~x2 & ~x5 ;
  assign n47 = ~n45 & n46 ;
  assign n48 = x1 & ~n47 ;
  assign n49 = n18 & n48 ;
  assign n50 = n49 ^ n18 ;
  assign n51 = n17 & n50 ;
  assign y0 = n51 ;
endmodule
