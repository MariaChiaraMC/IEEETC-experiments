// Benchmark "./radd.pla" written by ABC on Thu Apr 23 11:00:00 2020

module \./radd.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z0  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z0;
  assign z0 = 1'b1;
endmodule


