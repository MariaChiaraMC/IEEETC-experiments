module top( x0 , x1 , x2 , x3 , x4 , y0 );
  input x0 , x1 , x2 , x3 , x4 ;
  output y0 ;
  wire n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 ;
  assign n6 = x3 ^ x1 ;
  assign n7 = n6 ^ x4 ;
  assign n8 = x4 ^ x3 ;
  assign n9 = n8 ^ x3 ;
  assign n10 = n9 ^ n7 ;
  assign n11 = x3 ^ x0 ;
  assign n12 = n11 ^ x2 ;
  assign n13 = ~x2 & ~n12 ;
  assign n14 = n13 ^ x3 ;
  assign n15 = n14 ^ x2 ;
  assign n16 = n10 & ~n15 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n17 ^ x2 ;
  assign n19 = ~n7 & ~n18 ;
  assign y0 = n19 ;
endmodule
