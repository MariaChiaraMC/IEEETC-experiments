module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 ;
  output y0 ;
  wire n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 ;
  assign n21 = ~x0 & x1 ;
  assign n22 = n21 ^ x5 ;
  assign n23 = n22 ^ x2 ;
  assign n24 = n23 ^ n22 ;
  assign n28 = n22 ^ x3 ;
  assign n29 = n22 & n28 ;
  assign n25 = x0 & ~x1 ;
  assign n26 = x5 & ~n25 ;
  assign n32 = n29 ^ n26 ;
  assign n27 = n26 ^ n24 ;
  assign n30 = n29 ^ n22 ;
  assign n31 = n27 & n30 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = n24 & n33 ;
  assign n35 = n34 ^ n29 ;
  assign n36 = n35 ^ n31 ;
  assign n37 = n36 ^ x5 ;
  assign n38 = ~x4 & n37 ;
  assign n39 = ~x18 & ~x19 ;
  assign n40 = ~x9 & n25 ;
  assign n41 = x5 & ~x12 ;
  assign n42 = ~x16 & n41 ;
  assign n43 = ~n40 & ~n42 ;
  assign n44 = ~x8 & ~n43 ;
  assign n45 = ~x0 & ~x1 ;
  assign n46 = ~x4 & x9 ;
  assign n47 = ~n45 & n46 ;
  assign n48 = ~x0 & ~x15 ;
  assign n49 = ~x12 & ~x13 ;
  assign n50 = x8 & n49 ;
  assign n51 = ~n48 & n50 ;
  assign n52 = ~x6 & ~x7 ;
  assign n53 = n51 & n52 ;
  assign n54 = n47 & n53 ;
  assign n55 = ~n44 & ~n54 ;
  assign n56 = x11 & ~n55 ;
  assign n57 = ~x7 & ~x15 ;
  assign n58 = x11 & n57 ;
  assign n59 = ~x9 & ~x11 ;
  assign n60 = ~x7 & ~x8 ;
  assign n61 = ~n59 & n60 ;
  assign n62 = n41 & ~n61 ;
  assign n63 = ~n58 & n62 ;
  assign n64 = ~n56 & ~n63 ;
  assign n65 = ~x10 & ~n64 ;
  assign n66 = x6 & ~x11 ;
  assign n67 = ~x8 & ~x11 ;
  assign n68 = ~x9 & ~n67 ;
  assign n69 = x10 & x15 ;
  assign n70 = ~n68 & n69 ;
  assign n71 = ~n66 & ~n70 ;
  assign n72 = n59 ^ x7 ;
  assign n78 = n72 ^ n59 ;
  assign n79 = n78 ^ x8 ;
  assign n80 = n79 ^ x8 ;
  assign n81 = n72 ^ x16 ;
  assign n82 = n81 ^ x8 ;
  assign n83 = ~n80 & n82 ;
  assign n73 = n72 ^ n57 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = n74 ^ n59 ;
  assign n76 = n75 ^ x8 ;
  assign n77 = ~n59 & ~n76 ;
  assign n84 = n83 ^ n77 ;
  assign n85 = n84 ^ n59 ;
  assign n86 = n77 ^ x8 ;
  assign n87 = n86 ^ n79 ;
  assign n88 = ~x8 & ~n87 ;
  assign n89 = n88 ^ n77 ;
  assign n90 = ~n85 & n89 ;
  assign n91 = n90 ^ n83 ;
  assign n92 = n91 ^ n88 ;
  assign n93 = n92 ^ n59 ;
  assign n94 = n93 ^ x8 ;
  assign n95 = n94 ^ n79 ;
  assign n96 = n95 ^ x7 ;
  assign n97 = n71 & ~n96 ;
  assign n98 = ~x12 & ~n97 ;
  assign n99 = ~x8 & x16 ;
  assign n100 = ~x9 & ~x10 ;
  assign n101 = n58 & n100 ;
  assign n102 = n99 & n101 ;
  assign n103 = x13 & ~n102 ;
  assign n104 = x6 & ~x7 ;
  assign n105 = ~n103 & ~n104 ;
  assign n106 = ~x17 & n105 ;
  assign n107 = ~n98 & n106 ;
  assign n108 = x5 & ~n107 ;
  assign n109 = ~n65 & ~n108 ;
  assign n110 = x2 & ~x3 ;
  assign n111 = ~n109 & n110 ;
  assign n112 = x2 & x4 ;
  assign n113 = n21 & n112 ;
  assign n114 = ~x2 & ~x3 ;
  assign n115 = x2 ^ x1 ;
  assign n116 = n114 & ~n115 ;
  assign n117 = n116 ^ n115 ;
  assign n118 = x5 & ~n117 ;
  assign n119 = x3 & ~x5 ;
  assign n120 = n119 ^ x4 ;
  assign n121 = n120 ^ n119 ;
  assign n122 = ~x11 & ~x13 ;
  assign n123 = ~x12 & n122 ;
  assign n124 = n110 & n123 ;
  assign n125 = n52 & ~n100 ;
  assign n126 = n125 ^ x8 ;
  assign n127 = n126 ^ n125 ;
  assign n128 = x9 & x10 ;
  assign n129 = n128 ^ n125 ;
  assign n130 = n127 & n129 ;
  assign n131 = n130 ^ n125 ;
  assign n132 = n124 & n131 ;
  assign n133 = n132 ^ n119 ;
  assign n134 = ~n121 & n133 ;
  assign n135 = n134 ^ n119 ;
  assign n136 = ~n45 & n135 ;
  assign n137 = ~n118 & ~n136 ;
  assign n138 = ~n113 & n137 ;
  assign n139 = x11 ^ x10 ;
  assign n140 = ~x1 & x3 ;
  assign n141 = ~x2 & n140 ;
  assign n142 = ~x5 & ~n141 ;
  assign n143 = n142 ^ x11 ;
  assign n144 = n143 ^ n142 ;
  assign n145 = n144 ^ n139 ;
  assign n146 = ~x0 & ~x2 ;
  assign n147 = ~n140 & ~n146 ;
  assign n148 = n147 ^ n52 ;
  assign n149 = ~n147 & ~n148 ;
  assign n150 = n149 ^ n142 ;
  assign n151 = n150 ^ n147 ;
  assign n152 = n145 & n151 ;
  assign n153 = n152 ^ n149 ;
  assign n154 = n153 ^ n147 ;
  assign n155 = n139 & ~n154 ;
  assign n156 = x8 & n155 ;
  assign n157 = ~x2 & x5 ;
  assign n158 = ~n156 & ~n157 ;
  assign n159 = x9 & n49 ;
  assign n160 = ~n158 & n159 ;
  assign n161 = ~x12 & n52 ;
  assign n162 = ~x13 & ~n161 ;
  assign n163 = x5 & x11 ;
  assign n164 = n100 & ~n163 ;
  assign n165 = ~n162 & ~n164 ;
  assign n166 = ~x9 & ~n45 ;
  assign n167 = ~n141 & ~n146 ;
  assign n168 = ~n166 & ~n167 ;
  assign n169 = ~x5 & ~n168 ;
  assign n170 = ~n100 & ~n122 ;
  assign n171 = ~x8 & ~n170 ;
  assign n172 = ~n169 & n171 ;
  assign n173 = n165 & n172 ;
  assign n174 = ~n160 & ~n173 ;
  assign n175 = n174 ^ x3 ;
  assign n176 = n175 ^ x4 ;
  assign n232 = n176 ^ n175 ;
  assign n177 = x5 ^ x4 ;
  assign n178 = n146 ^ x5 ;
  assign n179 = n178 ^ n146 ;
  assign n180 = x12 ^ x11 ;
  assign n181 = n180 ^ x12 ;
  assign n182 = n181 ^ x12 ;
  assign n183 = n182 ^ x8 ;
  assign n184 = n181 ^ n139 ;
  assign n185 = n184 ^ n183 ;
  assign n186 = ~n183 & n185 ;
  assign n187 = n186 ^ x8 ;
  assign n188 = n181 ^ x8 ;
  assign n189 = n188 ^ n184 ;
  assign n192 = n184 ^ n182 ;
  assign n193 = x12 ^ x1 ;
  assign n194 = n192 & n193 ;
  assign n190 = x13 ^ x8 ;
  assign n191 = ~n188 & ~n190 ;
  assign n195 = n194 ^ n191 ;
  assign n196 = n195 ^ x12 ;
  assign n197 = n196 ^ n181 ;
  assign n198 = n197 ^ n184 ;
  assign n199 = n189 & n198 ;
  assign n200 = n199 ^ n191 ;
  assign n201 = n200 ^ n181 ;
  assign n202 = n201 ^ n184 ;
  assign n203 = n187 & n202 ;
  assign n204 = n203 ^ n191 ;
  assign n205 = n204 ^ n186 ;
  assign n206 = n205 ^ n199 ;
  assign n207 = n206 ^ n181 ;
  assign n208 = n207 ^ x8 ;
  assign n209 = n208 ^ n184 ;
  assign n210 = x9 & ~n209 ;
  assign n211 = x13 ^ x1 ;
  assign n212 = x13 ^ x0 ;
  assign n213 = n212 ^ x0 ;
  assign n214 = ~x2 & ~x12 ;
  assign n215 = n214 ^ x0 ;
  assign n216 = n213 & n215 ;
  assign n217 = n216 ^ x0 ;
  assign n218 = n211 & n217 ;
  assign n219 = n218 ^ x1 ;
  assign n220 = ~n210 & ~n219 ;
  assign n221 = n220 ^ n146 ;
  assign n222 = n179 & n221 ;
  assign n223 = n222 ^ n146 ;
  assign n224 = ~n177 & ~n223 ;
  assign n225 = n224 ^ x4 ;
  assign n226 = n225 ^ n176 ;
  assign n227 = n226 ^ n175 ;
  assign n228 = n176 ^ n174 ;
  assign n229 = n228 ^ n225 ;
  assign n230 = n229 ^ n227 ;
  assign n231 = ~n227 & n230 ;
  assign n233 = n232 ^ n231 ;
  assign n234 = n233 ^ n227 ;
  assign n235 = n175 ^ n25 ;
  assign n236 = n231 ^ n227 ;
  assign n237 = ~n235 & ~n236 ;
  assign n238 = n237 ^ n175 ;
  assign n239 = n234 & n238 ;
  assign n240 = n239 ^ n175 ;
  assign n241 = n240 ^ x3 ;
  assign n242 = n241 ^ n175 ;
  assign n243 = n138 & n242 ;
  assign n244 = ~n111 & n243 ;
  assign n245 = n39 & ~n244 ;
  assign n246 = x14 & ~n245 ;
  assign n247 = ~n38 & n246 ;
  assign y0 = ~n247 ;
endmodule
