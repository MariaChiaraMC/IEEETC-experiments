// Benchmark "./spla.pla" written by ABC on Thu Apr 23 11:00:01 2020

module \./spla.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15,
    z0  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15;
  output z0;
  wire new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_, new_n24_,
    new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_;
  assign new_n18_ = ~x7 & ~x10;
  assign new_n19_ = ~x2 & ~x14;
  assign new_n20_ = ~x4 & ~x6;
  assign new_n21_ = new_n19_ & new_n20_;
  assign new_n22_ = x5 & ~x11;
  assign new_n23_ = ~x9 & ~x12;
  assign new_n24_ = new_n22_ & new_n23_;
  assign new_n25_ = ~x3 & ~x15;
  assign new_n26_ = ~x8 & ~x13;
  assign new_n27_ = new_n25_ & new_n26_;
  assign new_n28_ = new_n24_ & new_n27_;
  assign new_n29_ = new_n21_ & new_n28_;
  assign new_n30_ = new_n18_ & new_n29_;
  assign z0 = ~x1 | new_n30_;
endmodule


