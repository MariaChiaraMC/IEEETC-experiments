module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 ;
  assign n11 = ~x0 & ~x2 ;
  assign n12 = x3 & n11 ;
  assign n13 = x6 & ~n12 ;
  assign n14 = ~x1 & x6 ;
  assign n15 = x3 ^ x2 ;
  assign n16 = ~x8 & ~x9 ;
  assign n17 = n16 ^ x3 ;
  assign n18 = n16 ^ x1 ;
  assign n19 = ~n16 & n18 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = ~n17 & ~n20 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = n23 ^ x1 ;
  assign n25 = n15 & n24 ;
  assign n26 = x0 & n25 ;
  assign n27 = ~n14 & ~n26 ;
  assign n28 = ~n13 & ~n27 ;
  assign n29 = ~x0 & ~x3 ;
  assign n30 = ~x2 & x6 ;
  assign n31 = x8 & ~x9 ;
  assign n32 = x1 & n31 ;
  assign n33 = n30 & n32 ;
  assign n34 = n29 & n33 ;
  assign n35 = ~n28 & ~n34 ;
  assign n57 = ~x0 & x1 ;
  assign n115 = ~x2 & ~x3 ;
  assign n116 = x8 & n115 ;
  assign n117 = x6 & ~n116 ;
  assign n118 = n57 & n117 ;
  assign n36 = x0 & ~x3 ;
  assign n37 = x1 & n36 ;
  assign n38 = x2 & ~x6 ;
  assign n39 = ~n16 & n38 ;
  assign n40 = x8 & x9 ;
  assign n41 = ~x2 & ~x6 ;
  assign n42 = ~n40 & n41 ;
  assign n43 = ~n39 & ~n42 ;
  assign n44 = n37 & ~n43 ;
  assign n45 = x1 & ~n30 ;
  assign n46 = x2 & ~x9 ;
  assign n47 = ~x8 & ~n46 ;
  assign n48 = ~n45 & n47 ;
  assign n49 = ~n30 & ~n46 ;
  assign n50 = x8 & ~n14 ;
  assign n51 = ~n49 & n50 ;
  assign n52 = ~x8 & x9 ;
  assign n53 = ~x6 & n52 ;
  assign n54 = x0 & ~n53 ;
  assign n55 = ~n51 & n54 ;
  assign n56 = ~n48 & n55 ;
  assign n58 = n30 & ~n31 ;
  assign n59 = n39 & ~n40 ;
  assign n60 = ~n58 & ~n59 ;
  assign n61 = n57 & ~n60 ;
  assign n62 = ~n56 & ~n61 ;
  assign n63 = x3 & ~n62 ;
  assign n64 = n63 ^ n44 ;
  assign n65 = x3 & x9 ;
  assign n66 = x1 & ~n41 ;
  assign n67 = x2 & ~x8 ;
  assign n68 = ~n41 & ~n67 ;
  assign n69 = ~n66 & ~n68 ;
  assign n70 = n65 & n69 ;
  assign n71 = x6 & n32 ;
  assign n72 = x2 & n71 ;
  assign n73 = ~n70 & ~n72 ;
  assign n74 = n73 ^ x0 ;
  assign n75 = n74 ^ n73 ;
  assign n80 = x9 ^ x8 ;
  assign n77 = x9 ^ x3 ;
  assign n76 = x8 ^ x1 ;
  assign n78 = n77 ^ n76 ;
  assign n79 = n78 ^ x8 ;
  assign n81 = n80 ^ n79 ;
  assign n82 = n76 ^ x9 ;
  assign n83 = n82 ^ x8 ;
  assign n84 = n83 ^ x8 ;
  assign n85 = n78 & ~n84 ;
  assign n86 = n85 ^ n78 ;
  assign n87 = ~n83 & n86 ;
  assign n88 = n87 ^ x8 ;
  assign n89 = ~n81 & n88 ;
  assign n90 = n89 ^ n85 ;
  assign n91 = n90 ^ x8 ;
  assign n92 = n91 ^ x1 ;
  assign n93 = n92 ^ n80 ;
  assign n94 = n30 & ~n93 ;
  assign n95 = n94 ^ n73 ;
  assign n96 = n75 & ~n95 ;
  assign n97 = n96 ^ n73 ;
  assign n98 = n97 ^ n44 ;
  assign n99 = n64 & ~n98 ;
  assign n100 = n99 ^ n96 ;
  assign n101 = n100 ^ n73 ;
  assign n102 = n101 ^ n63 ;
  assign n103 = ~n44 & ~n102 ;
  assign n104 = n103 ^ n44 ;
  assign n119 = n118 ^ n104 ;
  assign n120 = n119 ^ n104 ;
  assign n105 = x2 ^ x0 ;
  assign n106 = n105 ^ x2 ;
  assign n107 = x8 & n65 ;
  assign n108 = ~x6 & n107 ;
  assign n109 = n108 ^ x2 ;
  assign n110 = n106 & n109 ;
  assign n111 = n110 ^ x2 ;
  assign n112 = ~x1 & n111 ;
  assign n113 = n112 ^ n104 ;
  assign n114 = n113 ^ n104 ;
  assign n121 = n120 ^ n114 ;
  assign n122 = ~x2 & n80 ;
  assign n123 = n37 & ~n122 ;
  assign n124 = ~x3 & ~x9 ;
  assign n125 = ~n67 & ~n124 ;
  assign n126 = n57 & ~n125 ;
  assign n127 = n12 & ~n16 ;
  assign n128 = ~n126 & ~n127 ;
  assign n129 = ~n123 & n128 ;
  assign n130 = ~x6 & ~n129 ;
  assign n131 = n130 ^ n104 ;
  assign n132 = n131 ^ n104 ;
  assign n133 = n132 ^ n120 ;
  assign n134 = ~n120 & n133 ;
  assign n135 = n134 ^ n120 ;
  assign n136 = n121 & ~n135 ;
  assign n137 = n136 ^ n134 ;
  assign n138 = n137 ^ n104 ;
  assign n139 = n138 ^ n120 ;
  assign n140 = x5 & n139 ;
  assign n141 = n140 ^ n104 ;
  assign n142 = n35 & ~n141 ;
  assign n143 = ~x4 & ~n142 ;
  assign n144 = ~x2 & x4 ;
  assign n145 = ~x1 & n144 ;
  assign n146 = n145 ^ x5 ;
  assign n147 = n146 ^ n145 ;
  assign n148 = n147 ^ n29 ;
  assign n149 = n16 ^ x2 ;
  assign n150 = n149 ^ n16 ;
  assign n151 = n40 ^ n16 ;
  assign n152 = n151 ^ n16 ;
  assign n153 = n150 & ~n152 ;
  assign n154 = n153 ^ n16 ;
  assign n155 = ~x6 & n154 ;
  assign n156 = n155 ^ n16 ;
  assign n158 = n156 ^ x2 ;
  assign n157 = n156 ^ n52 ;
  assign n159 = n158 ^ n157 ;
  assign n160 = n158 ^ x6 ;
  assign n161 = n160 ^ n158 ;
  assign n162 = n159 & n161 ;
  assign n163 = n162 ^ n158 ;
  assign n164 = x1 & n163 ;
  assign n165 = n164 ^ n156 ;
  assign n166 = ~x4 & n165 ;
  assign n167 = x9 ^ x6 ;
  assign n168 = x8 & n167 ;
  assign n169 = n168 ^ x6 ;
  assign n170 = n145 & ~n169 ;
  assign n171 = n170 ^ n166 ;
  assign n172 = ~n166 & n171 ;
  assign n173 = n172 ^ n145 ;
  assign n174 = n173 ^ n166 ;
  assign n175 = ~n148 & n174 ;
  assign n176 = n175 ^ n172 ;
  assign n177 = n176 ^ n166 ;
  assign n178 = n29 & ~n177 ;
  assign n179 = n178 ^ n29 ;
  assign n180 = ~n143 & ~n179 ;
  assign n181 = ~x7 & ~n180 ;
  assign n182 = ~x4 & ~x5 ;
  assign n183 = ~x9 & n57 ;
  assign n184 = n18 ^ n16 ;
  assign n185 = x7 & n40 ;
  assign n186 = n185 ^ n16 ;
  assign n187 = n184 & n186 ;
  assign n188 = n187 ^ n16 ;
  assign n189 = x0 & n188 ;
  assign n190 = ~n183 & ~n189 ;
  assign n191 = ~x3 & n41 ;
  assign n192 = ~n190 & n191 ;
  assign n193 = n182 & n192 ;
  assign n194 = ~n181 & ~n193 ;
  assign y0 = ~n194 ;
endmodule
