module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
  assign n9 = ~x2 & x3 ;
  assign n10 = n9 ^ x1 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = ~x6 & x7 ;
  assign n13 = x4 & ~n12 ;
  assign n14 = x2 & ~x5 ;
  assign n15 = ~n13 & ~n14 ;
  assign n16 = ~x3 & ~n15 ;
  assign n17 = ~x3 & x6 ;
  assign n18 = ~x7 & n17 ;
  assign n19 = n18 ^ x5 ;
  assign n20 = n18 ^ x4 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = n9 ^ x2 ;
  assign n23 = ~x4 & ~n22 ;
  assign n24 = n23 ^ n9 ;
  assign n25 = ~n21 & n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n26 ^ n9 ;
  assign n28 = n27 ^ x4 ;
  assign n29 = ~n19 & ~n28 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = ~n16 & ~n30 ;
  assign n32 = n31 ^ n9 ;
  assign n33 = ~n11 & n32 ;
  assign n34 = n33 ^ n9 ;
  assign n35 = ~x0 & n34 ;
  assign y0 = n35 ;
endmodule
