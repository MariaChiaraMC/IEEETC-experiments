module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 ;
  assign n9 = ~x5 & x7 ;
  assign n10 = x3 & ~x6 ;
  assign n11 = ~x1 & ~x4 ;
  assign n12 = n10 & n11 ;
  assign n13 = n9 & n12 ;
  assign n19 = x5 ^ x3 ;
  assign n14 = x3 ^ x1 ;
  assign n16 = n14 ^ x6 ;
  assign n15 = n14 ^ x5 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n17 ^ n14 ;
  assign n27 = n18 ^ n16 ;
  assign n28 = n27 ^ n14 ;
  assign n20 = n19 ^ x7 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n21 ^ n19 ;
  assign n29 = n28 ^ n22 ;
  assign n30 = n29 ^ n19 ;
  assign n31 = ~n19 & n30 ;
  assign n32 = n31 ^ n18 ;
  assign n33 = n32 ^ n22 ;
  assign n34 = n33 ^ n19 ;
  assign n35 = n34 ^ n14 ;
  assign n36 = n22 ^ n19 ;
  assign n37 = n36 ^ n14 ;
  assign n38 = ~n33 & n37 ;
  assign n39 = n38 ^ n18 ;
  assign n40 = n39 ^ n22 ;
  assign n41 = n40 ^ n19 ;
  assign n42 = n41 ^ n14 ;
  assign n43 = n35 & n42 ;
  assign n23 = n22 ^ n18 ;
  assign n24 = n23 ^ n19 ;
  assign n25 = n24 ^ n14 ;
  assign n26 = n24 & n25 ;
  assign n44 = n43 ^ n26 ;
  assign n45 = n44 ^ n31 ;
  assign n46 = n45 ^ n18 ;
  assign n47 = n46 ^ n22 ;
  assign n48 = n47 ^ n19 ;
  assign n49 = n48 ^ n14 ;
  assign n50 = x4 & n49 ;
  assign n51 = ~x2 & ~n50 ;
  assign n52 = ~n13 & n51 ;
  assign n53 = ~x0 & ~n52 ;
  assign n54 = x5 ^ x4 ;
  assign n55 = x2 & ~n54 ;
  assign n56 = ~x1 & x6 ;
  assign n57 = ~x3 & n56 ;
  assign n58 = n57 ^ x1 ;
  assign n59 = x5 ^ x1 ;
  assign n60 = n59 ^ x1 ;
  assign n61 = n60 ^ n55 ;
  assign n62 = n58 & n61 ;
  assign n63 = n62 ^ n57 ;
  assign n64 = n55 & n63 ;
  assign n65 = n64 ^ x2 ;
  assign n66 = n53 & ~n65 ;
  assign y0 = n66 ;
endmodule
