module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 ;
  assign n10 = x1 ^ x0 ;
  assign n11 = ~x6 & x7 ;
  assign n12 = ~x5 & n11 ;
  assign n13 = x4 & n12 ;
  assign n14 = x6 & x7 ;
  assign n15 = x0 & x5 ;
  assign n16 = n14 & n15 ;
  assign n17 = ~n13 & ~n16 ;
  assign n18 = n17 ^ x8 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = x5 & ~x6 ;
  assign n21 = ~x7 & ~n20 ;
  assign n22 = ~x4 & ~n21 ;
  assign n23 = x6 & ~x7 ;
  assign n24 = n15 & n23 ;
  assign n25 = ~n22 & ~n24 ;
  assign n26 = n25 ^ x0 ;
  assign n27 = n25 ^ n11 ;
  assign n28 = n27 ^ n11 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = x4 & x6 ;
  assign n31 = n30 ^ x5 ;
  assign n32 = n30 & ~n31 ;
  assign n33 = n32 ^ n11 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = ~n29 & n34 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = ~n26 & n37 ;
  assign n39 = n38 ^ n25 ;
  assign n40 = n39 ^ n17 ;
  assign n41 = ~n19 & n40 ;
  assign n42 = n41 ^ n17 ;
  assign n43 = ~x2 & ~n42 ;
  assign n44 = n43 ^ n10 ;
  assign n45 = n44 ^ x1 ;
  assign n46 = n45 ^ n44 ;
  assign n47 = ~x5 & x6 ;
  assign n48 = x1 & n47 ;
  assign n49 = ~x2 & ~x6 ;
  assign n50 = ~x5 & n49 ;
  assign n51 = n50 ^ x2 ;
  assign n52 = n51 ^ n50 ;
  assign n53 = n50 ^ x1 ;
  assign n54 = n53 ^ n50 ;
  assign n55 = ~n52 & n54 ;
  assign n56 = n55 ^ n50 ;
  assign n57 = x7 & n56 ;
  assign n58 = n57 ^ n50 ;
  assign n59 = ~n48 & ~n58 ;
  assign n60 = ~x8 & ~n59 ;
  assign n61 = ~x6 & ~x8 ;
  assign n62 = ~n23 & ~n61 ;
  assign n63 = x1 & ~x5 ;
  assign n64 = ~n11 & n63 ;
  assign n65 = n62 & n64 ;
  assign n66 = x6 & x8 ;
  assign n67 = ~x7 & n66 ;
  assign n68 = x5 & n67 ;
  assign n69 = ~n65 & ~n68 ;
  assign n70 = ~n60 & n69 ;
  assign n71 = x2 & x5 ;
  assign n72 = x7 ^ x6 ;
  assign n73 = n71 & ~n72 ;
  assign n74 = n70 & ~n73 ;
  assign n75 = x4 & ~n74 ;
  assign n76 = ~x4 & ~x7 ;
  assign n77 = ~x2 & n47 ;
  assign n78 = x5 & ~x8 ;
  assign n79 = ~n77 & ~n78 ;
  assign n80 = n76 & ~n79 ;
  assign n81 = x1 & n80 ;
  assign n82 = ~x4 & n20 ;
  assign n83 = ~x2 & x7 ;
  assign n84 = n83 ^ x2 ;
  assign n85 = x8 & n84 ;
  assign n86 = n85 ^ x2 ;
  assign n87 = n82 & n86 ;
  assign n88 = ~x5 & x8 ;
  assign n89 = ~x6 & ~x7 ;
  assign n90 = x2 & n89 ;
  assign n91 = n88 & n90 ;
  assign n92 = ~x2 & x5 ;
  assign n93 = ~x8 & n14 ;
  assign n94 = n92 & n93 ;
  assign n95 = ~n91 & ~n94 ;
  assign n96 = ~n87 & n95 ;
  assign n97 = ~n81 & n96 ;
  assign n98 = ~n75 & n97 ;
  assign n99 = n98 ^ n44 ;
  assign n100 = n99 ^ n10 ;
  assign n101 = ~n46 & n100 ;
  assign n102 = n101 ^ n98 ;
  assign n103 = ~x4 & ~x8 ;
  assign n104 = n71 & n103 ;
  assign n106 = n88 ^ x7 ;
  assign n113 = n106 ^ n88 ;
  assign n105 = n88 ^ x2 ;
  assign n107 = n106 ^ n105 ;
  assign n108 = n107 ^ n88 ;
  assign n109 = n105 ^ x6 ;
  assign n110 = n109 ^ n105 ;
  assign n111 = n110 ^ n108 ;
  assign n112 = n108 & ~n111 ;
  assign n114 = n113 ^ n112 ;
  assign n115 = n114 ^ n108 ;
  assign n116 = n88 ^ x4 ;
  assign n117 = n116 ^ n88 ;
  assign n118 = n112 ^ n108 ;
  assign n119 = ~n117 & n118 ;
  assign n120 = n119 ^ n88 ;
  assign n121 = n115 & n120 ;
  assign n122 = n121 ^ n88 ;
  assign n123 = n122 ^ n88 ;
  assign n124 = n123 ^ n88 ;
  assign n125 = ~n104 & ~n124 ;
  assign n126 = x6 ^ x4 ;
  assign n127 = n126 ^ x6 ;
  assign n128 = n66 ^ x6 ;
  assign n129 = ~n127 & ~n128 ;
  assign n130 = n129 ^ x6 ;
  assign n131 = n92 & ~n130 ;
  assign n132 = n125 & ~n131 ;
  assign n133 = n98 & n132 ;
  assign n134 = n133 ^ n10 ;
  assign n135 = n102 & ~n134 ;
  assign n136 = n135 ^ n133 ;
  assign n137 = ~n10 & n136 ;
  assign n138 = n137 ^ n101 ;
  assign n139 = n138 ^ x0 ;
  assign n140 = n139 ^ n98 ;
  assign n141 = ~x3 & ~n140 ;
  assign n142 = ~x1 & x3 ;
  assign n143 = n23 & n142 ;
  assign n144 = x2 & ~n143 ;
  assign n145 = ~x5 & ~x8 ;
  assign n146 = ~n144 & n145 ;
  assign n147 = ~x2 & ~n11 ;
  assign n148 = n147 ^ n89 ;
  assign n149 = n148 ^ n89 ;
  assign n150 = n89 ^ x3 ;
  assign n151 = n150 ^ n89 ;
  assign n152 = ~n149 & n151 ;
  assign n153 = n152 ^ n89 ;
  assign n154 = ~x1 & n153 ;
  assign n155 = n154 ^ n89 ;
  assign n156 = n146 & n155 ;
  assign n157 = n77 ^ x1 ;
  assign n158 = n157 ^ n77 ;
  assign n164 = n77 ^ x8 ;
  assign n165 = ~n77 & n164 ;
  assign n159 = x8 ^ x6 ;
  assign n160 = x5 ^ x1 ;
  assign n161 = n160 ^ x8 ;
  assign n162 = n159 & ~n161 ;
  assign n168 = n165 ^ n162 ;
  assign n163 = n162 ^ n158 ;
  assign n166 = n165 ^ n77 ;
  assign n167 = n163 & ~n166 ;
  assign n169 = n168 ^ n167 ;
  assign n170 = n158 & n169 ;
  assign n171 = n170 ^ n165 ;
  assign n172 = n171 ^ n167 ;
  assign n173 = n172 ^ x1 ;
  assign n174 = x7 & ~n173 ;
  assign n175 = x1 & x8 ;
  assign n176 = ~n50 & ~n71 ;
  assign n177 = n175 & ~n176 ;
  assign n178 = ~n68 & ~n177 ;
  assign n179 = ~n174 & n178 ;
  assign n180 = x3 & ~n179 ;
  assign n181 = x8 & n83 ;
  assign n182 = ~n67 & ~n93 ;
  assign n183 = x2 & ~n182 ;
  assign n184 = ~n181 & ~n183 ;
  assign n185 = n63 & ~n184 ;
  assign n186 = ~x2 & n89 ;
  assign n187 = ~x8 & n186 ;
  assign n188 = n187 ^ n91 ;
  assign n189 = x1 & n188 ;
  assign n190 = n189 ^ n91 ;
  assign n191 = ~n185 & ~n190 ;
  assign n192 = ~n180 & n191 ;
  assign n193 = n192 ^ x4 ;
  assign n194 = n193 ^ n192 ;
  assign n195 = n194 ^ n156 ;
  assign n196 = ~n23 & ~n49 ;
  assign n197 = n142 & n196 ;
  assign n198 = ~x2 & x3 ;
  assign n199 = ~n11 & ~n198 ;
  assign n200 = x1 & ~n83 ;
  assign n201 = ~n199 & n200 ;
  assign n202 = ~n197 & ~n201 ;
  assign n203 = x5 & ~n202 ;
  assign n204 = n47 & n83 ;
  assign n205 = n12 ^ x2 ;
  assign n206 = n205 ^ n12 ;
  assign n207 = n206 ^ n204 ;
  assign n208 = n89 & n150 ;
  assign n209 = n208 ^ n12 ;
  assign n210 = n209 ^ n89 ;
  assign n211 = n207 & n210 ;
  assign n212 = n211 ^ n208 ;
  assign n213 = n212 ^ n89 ;
  assign n214 = ~n204 & n213 ;
  assign n215 = n214 ^ n204 ;
  assign n216 = ~x1 & n215 ;
  assign n217 = ~n203 & ~n216 ;
  assign n218 = x8 & n217 ;
  assign n219 = ~x7 & ~n71 ;
  assign n220 = ~x1 & ~n219 ;
  assign n221 = x6 ^ x5 ;
  assign n222 = n221 ^ x6 ;
  assign n223 = n11 ^ x6 ;
  assign n224 = n222 & ~n223 ;
  assign n225 = n224 ^ x6 ;
  assign n226 = x1 & n225 ;
  assign n227 = n226 ^ x5 ;
  assign n228 = n227 ^ x2 ;
  assign n229 = n228 ^ n227 ;
  assign n230 = x3 & ~n47 ;
  assign n231 = n230 ^ n227 ;
  assign n232 = n229 & n231 ;
  assign n233 = n232 ^ n227 ;
  assign n234 = ~n220 & n233 ;
  assign n235 = ~x8 & ~n234 ;
  assign n236 = n235 ^ n218 ;
  assign n237 = ~n218 & n236 ;
  assign n238 = n237 ^ n192 ;
  assign n239 = n238 ^ n218 ;
  assign n240 = ~n195 & n239 ;
  assign n241 = n240 ^ n237 ;
  assign n242 = n241 ^ n218 ;
  assign n243 = ~n156 & ~n242 ;
  assign n244 = n243 ^ n156 ;
  assign n245 = ~x0 & n244 ;
  assign n246 = ~n141 & ~n245 ;
  assign y0 = ~n246 ;
endmodule
