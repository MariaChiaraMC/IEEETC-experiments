module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n11 = x9 ^ x8 ;
  assign n12 = ~x2 & n11 ;
  assign n13 = n12 ^ x8 ;
  assign n15 = n13 ^ x4 ;
  assign n14 = n13 ^ x5 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n15 ^ x2 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n16 & ~n18 ;
  assign n20 = n19 ^ n15 ;
  assign n21 = x0 & n20 ;
  assign n22 = n21 ^ n13 ;
  assign n23 = ~x1 & n22 ;
  assign n24 = x3 ^ x0 ;
  assign n25 = n24 ^ x3 ;
  assign n26 = n25 ^ x1 ;
  assign n28 = x7 ^ x6 ;
  assign n29 = x6 ^ x2 ;
  assign n30 = n29 ^ x6 ;
  assign n31 = n28 & ~n30 ;
  assign n27 = x6 ^ x3 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = ~n26 & n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n34 ^ x3 ;
  assign n36 = n35 ^ n27 ;
  assign n37 = x1 & n36 ;
  assign n38 = ~n23 & ~n37 ;
  assign y0 = ~n38 ;
endmodule
