module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 ;
  assign n17 = ~x13 & ~x14 ;
  assign n18 = x10 & ~x11 ;
  assign n19 = n17 & n18 ;
  assign n20 = ~x12 & ~x15 ;
  assign n21 = x0 & x9 ;
  assign n22 = n20 & n21 ;
  assign n23 = n19 & n22 ;
  assign n24 = x5 & x6 ;
  assign n26 = ~x14 & ~x15 ;
  assign n27 = x11 ^ x2 ;
  assign n28 = n27 ^ x2 ;
  assign n29 = n24 ^ x2 ;
  assign n30 = n28 & n29 ;
  assign n31 = n30 ^ x2 ;
  assign n32 = ~x12 & ~n31 ;
  assign n33 = n32 ^ x11 ;
  assign n34 = ~n26 & ~n33 ;
  assign n25 = x11 & x12 ;
  assign n35 = n34 ^ n25 ;
  assign n36 = n24 & ~n35 ;
  assign n37 = ~x8 & x12 ;
  assign n38 = ~x1 & n37 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = x11 & ~n25 ;
  assign n41 = n40 ^ n36 ;
  assign n42 = n39 & n41 ;
  assign n43 = n42 ^ n40 ;
  assign n44 = n36 & n43 ;
  assign n45 = n44 ^ n34 ;
  assign n46 = n45 ^ x4 ;
  assign n47 = n46 ^ n45 ;
  assign n48 = n47 ^ x13 ;
  assign n49 = x3 & ~x11 ;
  assign n50 = ~x2 & n49 ;
  assign n51 = x14 ^ x5 ;
  assign n65 = n51 ^ x5 ;
  assign n55 = x6 ^ x5 ;
  assign n56 = n55 ^ n51 ;
  assign n57 = n56 ^ x5 ;
  assign n52 = x12 ^ x7 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n53 ^ x5 ;
  assign n58 = n57 ^ n54 ;
  assign n59 = x15 ^ x12 ;
  assign n60 = n51 ^ x12 ;
  assign n61 = n60 ^ x5 ;
  assign n62 = ~n59 & n61 ;
  assign n63 = n62 ^ n53 ;
  assign n64 = ~n58 & n63 ;
  assign n66 = n65 ^ n64 ;
  assign n67 = n66 ^ n57 ;
  assign n68 = n67 ^ n58 ;
  assign n69 = n58 ^ n57 ;
  assign n70 = n65 ^ n63 ;
  assign n71 = n70 ^ n57 ;
  assign n72 = n71 ^ n58 ;
  assign n73 = ~n69 & ~n72 ;
  assign n74 = n73 ^ n53 ;
  assign n75 = ~n68 & n74 ;
  assign n76 = n75 ^ n64 ;
  assign n77 = n76 ^ n65 ;
  assign n78 = n77 ^ n57 ;
  assign n79 = n78 ^ n58 ;
  assign n80 = n50 & ~n79 ;
  assign n81 = x6 & x7 ;
  assign n82 = x15 & ~n81 ;
  assign n83 = n82 ^ x14 ;
  assign n84 = n83 ^ n82 ;
  assign n85 = n84 ^ n50 ;
  assign n86 = x6 & n20 ;
  assign n87 = x0 & x6 ;
  assign n88 = ~x1 & ~n87 ;
  assign n89 = x12 & ~n88 ;
  assign n90 = n89 ^ n86 ;
  assign n91 = ~n86 & n90 ;
  assign n92 = n91 ^ n82 ;
  assign n93 = n92 ^ n86 ;
  assign n94 = n85 & n93 ;
  assign n95 = n94 ^ n91 ;
  assign n96 = n95 ^ n86 ;
  assign n97 = n50 & ~n96 ;
  assign n98 = n97 ^ n50 ;
  assign n99 = ~x5 & n98 ;
  assign n100 = ~x6 & ~x7 ;
  assign n101 = x11 & ~x12 ;
  assign n102 = ~x2 & ~n26 ;
  assign n103 = n101 & n102 ;
  assign n104 = ~x11 & x12 ;
  assign n105 = ~x8 & n104 ;
  assign n106 = ~n103 & ~n105 ;
  assign n107 = n100 & ~n106 ;
  assign n108 = ~x0 & x14 ;
  assign n109 = x3 & x6 ;
  assign n110 = ~n108 & n109 ;
  assign n111 = n102 & n104 ;
  assign n112 = ~n110 & n111 ;
  assign n113 = ~n107 & ~n112 ;
  assign n114 = ~x1 & ~x5 ;
  assign n115 = ~n113 & n114 ;
  assign n116 = ~n99 & ~n115 ;
  assign n117 = ~x3 & ~n114 ;
  assign n118 = x5 & ~x7 ;
  assign n119 = x6 & n118 ;
  assign n120 = ~n117 & ~n119 ;
  assign n121 = x12 & ~n120 ;
  assign n122 = n100 & n114 ;
  assign n123 = n122 ^ x2 ;
  assign n124 = n122 ^ n37 ;
  assign n125 = n124 ^ n37 ;
  assign n126 = n101 ^ n37 ;
  assign n127 = ~n125 & n126 ;
  assign n128 = n127 ^ n37 ;
  assign n129 = ~n123 & n128 ;
  assign n130 = n129 ^ x2 ;
  assign n131 = ~n121 & ~n130 ;
  assign n132 = ~n25 & ~n26 ;
  assign n133 = ~n131 & n132 ;
  assign n134 = n116 & ~n133 ;
  assign n135 = n134 ^ n80 ;
  assign n136 = ~n80 & ~n135 ;
  assign n137 = n136 ^ n45 ;
  assign n138 = n137 ^ n80 ;
  assign n139 = n48 & n138 ;
  assign n140 = n139 ^ n136 ;
  assign n141 = n140 ^ n80 ;
  assign n142 = x13 & ~n141 ;
  assign n143 = n142 ^ x13 ;
  assign n144 = ~n23 & ~n143 ;
  assign y0 = ~n144 ;
endmodule
