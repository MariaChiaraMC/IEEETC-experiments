module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 ;
  assign n8 = ~x5 & ~x6 ;
  assign n9 = ~x4 & n8 ;
  assign n10 = x2 & ~x6 ;
  assign n11 = x4 & ~n10 ;
  assign n12 = x2 & ~x5 ;
  assign n13 = n12 ^ x6 ;
  assign n14 = n13 ^ x3 ;
  assign n15 = x2 ^ x0 ;
  assign n16 = ~x6 & ~n15 ;
  assign n17 = n16 ^ x0 ;
  assign n18 = ~n14 & ~n17 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n19 ^ x0 ;
  assign n21 = n20 ^ x6 ;
  assign n22 = x3 & n21 ;
  assign n23 = ~n11 & n22 ;
  assign n24 = n10 ^ x0 ;
  assign n25 = n24 ^ x0 ;
  assign n26 = ~x0 & x4 ;
  assign n27 = n26 ^ x0 ;
  assign n28 = n25 & n27 ;
  assign n29 = n28 ^ x0 ;
  assign n30 = x5 & n29 ;
  assign n31 = x5 ^ x2 ;
  assign n40 = n31 ^ x2 ;
  assign n32 = n31 ^ n15 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = n33 ^ x2 ;
  assign n35 = x4 & ~x6 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ n32 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = ~n34 & n38 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = n41 ^ n34 ;
  assign n43 = x6 ^ x2 ;
  assign n44 = n39 ^ n34 ;
  assign n45 = n43 & ~n44 ;
  assign n46 = n45 ^ x2 ;
  assign n47 = n42 & ~n46 ;
  assign n48 = n47 ^ x2 ;
  assign n49 = n48 ^ x5 ;
  assign n50 = n49 ^ x2 ;
  assign n51 = n50 ^ x2 ;
  assign n52 = n51 ^ n50 ;
  assign n53 = x4 & ~n8 ;
  assign n54 = n53 ^ n50 ;
  assign n55 = n54 ^ n50 ;
  assign n56 = ~n52 & ~n55 ;
  assign n57 = n56 ^ n50 ;
  assign n58 = ~x3 & ~n57 ;
  assign n59 = n58 ^ n50 ;
  assign n60 = ~n30 & n59 ;
  assign n61 = n60 ^ x1 ;
  assign n62 = n61 ^ n60 ;
  assign n63 = x0 & x3 ;
  assign n64 = n8 & n63 ;
  assign n65 = ~x3 & ~x5 ;
  assign n66 = x4 ^ x2 ;
  assign n67 = n66 ^ x2 ;
  assign n68 = n67 ^ n65 ;
  assign n69 = x0 & x6 ;
  assign n70 = n69 ^ x2 ;
  assign n71 = n68 & n70 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = n65 & n72 ;
  assign n74 = ~x0 & x6 ;
  assign n75 = n74 ^ x5 ;
  assign n76 = ~x2 & ~x3 ;
  assign n77 = n76 ^ n74 ;
  assign n78 = n77 ^ n76 ;
  assign n79 = n78 ^ n75 ;
  assign n80 = ~x2 & ~x6 ;
  assign n81 = n80 ^ x4 ;
  assign n82 = x4 & n81 ;
  assign n83 = n82 ^ n76 ;
  assign n84 = n83 ^ x4 ;
  assign n85 = ~n79 & ~n84 ;
  assign n86 = n85 ^ n82 ;
  assign n87 = n86 ^ x4 ;
  assign n88 = n75 & n87 ;
  assign n89 = n88 ^ n74 ;
  assign n90 = ~n73 & ~n89 ;
  assign n91 = ~n64 & n90 ;
  assign n92 = n91 ^ n60 ;
  assign n93 = n62 & n92 ;
  assign n94 = n93 ^ n60 ;
  assign n95 = ~n23 & n94 ;
  assign n96 = ~n9 & n95 ;
  assign y0 = ~n96 ;
endmodule
