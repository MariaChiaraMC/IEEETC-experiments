module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 ;
  assign n30 = ~x4 & x5 ;
  assign n50 = ~x1 & x6 ;
  assign n51 = n30 & ~n50 ;
  assign n20 = x2 & x5 ;
  assign n21 = x4 & x6 ;
  assign n22 = ~n20 & n21 ;
  assign n8 = x0 & x2 ;
  assign n24 = x4 & ~n8 ;
  assign n25 = x1 & ~n24 ;
  assign n23 = x6 ^ x5 ;
  assign n26 = n25 ^ n23 ;
  assign n31 = ~x0 & ~x2 ;
  assign n32 = n30 & ~n31 ;
  assign n33 = n32 ^ x6 ;
  assign n27 = x2 & ~x4 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = n28 ^ n25 ;
  assign n34 = n33 ^ n29 ;
  assign n35 = n33 ^ n32 ;
  assign n36 = n35 ^ n26 ;
  assign n37 = n34 & ~n36 ;
  assign n38 = n37 ^ n32 ;
  assign n39 = ~n25 & ~n32 ;
  assign n40 = n39 ^ n26 ;
  assign n41 = ~n38 & ~n40 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = ~n26 & n42 ;
  assign n44 = n43 ^ n37 ;
  assign n45 = n44 ^ x6 ;
  assign n46 = n45 ^ n32 ;
  assign n47 = ~n22 & ~n46 ;
  assign n52 = n51 ^ n47 ;
  assign n53 = n52 ^ n47 ;
  assign n9 = n8 ^ x1 ;
  assign n10 = n9 ^ x5 ;
  assign n11 = x6 ^ x2 ;
  assign n12 = ~x1 & n11 ;
  assign n13 = n12 ^ x2 ;
  assign n14 = ~n10 & ~n13 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n15 ^ x2 ;
  assign n17 = n16 ^ x1 ;
  assign n18 = ~x5 & n17 ;
  assign n19 = x4 & n18 ;
  assign n48 = n47 ^ n19 ;
  assign n49 = n48 ^ n47 ;
  assign n54 = n53 ^ n49 ;
  assign n55 = n20 & ~n21 ;
  assign n56 = n55 ^ n47 ;
  assign n57 = n56 ^ n47 ;
  assign n58 = n57 ^ n53 ;
  assign n59 = ~n53 & n58 ;
  assign n60 = n59 ^ n53 ;
  assign n61 = n54 & ~n60 ;
  assign n62 = n61 ^ n59 ;
  assign n63 = n62 ^ n47 ;
  assign n64 = n63 ^ n53 ;
  assign n65 = ~x3 & n64 ;
  assign n66 = n65 ^ n47 ;
  assign y0 = n66 ;
endmodule
