module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 ;
  assign n16 = x9 & x13 ;
  assign n17 = n16 ^ x11 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = n18 ^ x10 ;
  assign n20 = ~x3 & x14 ;
  assign n21 = ~x9 & ~n20 ;
  assign n22 = x6 & ~x14 ;
  assign n23 = ~x4 & ~x13 ;
  assign n24 = ~x7 & ~x8 ;
  assign n25 = ~x5 & ~n24 ;
  assign n26 = n23 & n25 ;
  assign n27 = n22 & n26 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = ~n21 & n28 ;
  assign n30 = n29 ^ n16 ;
  assign n31 = n30 ^ n21 ;
  assign n32 = n19 & n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ n21 ;
  assign n35 = ~x10 & ~n34 ;
  assign n36 = n35 ^ x10 ;
  assign n106 = x9 & ~x14 ;
  assign n107 = x10 & n106 ;
  assign n67 = ~x5 & x7 ;
  assign n108 = x10 & ~x14 ;
  assign n109 = x1 & n108 ;
  assign n110 = ~n16 & ~n109 ;
  assign n111 = n67 & ~n110 ;
  assign n112 = ~n107 & ~n111 ;
  assign n113 = ~x11 & ~n112 ;
  assign n90 = ~x11 & x13 ;
  assign n91 = ~x3 & n90 ;
  assign n114 = ~x9 & n91 ;
  assign n115 = x9 & ~x13 ;
  assign n116 = ~x3 & ~x14 ;
  assign n117 = ~n115 & ~n116 ;
  assign n118 = ~x11 & ~n117 ;
  assign n119 = ~n114 & ~n118 ;
  assign n120 = ~x7 & x10 ;
  assign n121 = x5 & n120 ;
  assign n122 = n121 ^ x10 ;
  assign n123 = ~n119 & n122 ;
  assign n124 = x5 & x14 ;
  assign n94 = ~x9 & ~x13 ;
  assign n62 = ~x1 & ~x6 ;
  assign n125 = ~x11 & n62 ;
  assign n126 = n94 & ~n125 ;
  assign n127 = n124 & n126 ;
  assign n128 = ~n123 & ~n127 ;
  assign n129 = ~n113 & n128 ;
  assign n130 = x4 & ~n129 ;
  assign n131 = x8 & x11 ;
  assign n132 = ~x3 & n131 ;
  assign n42 = x6 & x11 ;
  assign n133 = ~n22 & ~n42 ;
  assign n134 = ~n132 & n133 ;
  assign n135 = x4 & x11 ;
  assign n136 = n115 & ~n135 ;
  assign n137 = n120 & n136 ;
  assign n138 = ~n134 & n137 ;
  assign n139 = x10 ^ x6 ;
  assign n140 = n139 ^ n24 ;
  assign n141 = n23 ^ x6 ;
  assign n142 = n141 ^ n23 ;
  assign n143 = n106 ^ n23 ;
  assign n144 = ~n142 & n143 ;
  assign n145 = n144 ^ n23 ;
  assign n146 = n145 ^ n139 ;
  assign n147 = ~n140 & n146 ;
  assign n148 = n147 ^ n144 ;
  assign n149 = n148 ^ n23 ;
  assign n150 = n149 ^ n24 ;
  assign n151 = n139 & ~n150 ;
  assign n152 = n151 ^ n139 ;
  assign n153 = ~x11 & n152 ;
  assign n154 = ~n138 & ~n153 ;
  assign n155 = ~x5 & ~n154 ;
  assign n156 = ~x10 & n16 ;
  assign n157 = ~x10 & x11 ;
  assign n158 = x14 & n157 ;
  assign n159 = ~n156 & ~n158 ;
  assign n160 = ~n155 & n159 ;
  assign n161 = ~n130 & n160 ;
  assign n162 = ~x0 & ~n161 ;
  assign n163 = x14 ^ x3 ;
  assign n164 = x7 & x10 ;
  assign n165 = x4 & x6 ;
  assign n166 = x5 & n165 ;
  assign n167 = n164 & n166 ;
  assign n168 = n167 ^ x14 ;
  assign n169 = n168 ^ n167 ;
  assign n68 = x4 & n67 ;
  assign n170 = n167 ^ n68 ;
  assign n171 = ~n169 & n170 ;
  assign n172 = n171 ^ n167 ;
  assign n173 = n163 & ~n172 ;
  assign n174 = n173 ^ x3 ;
  assign n175 = n90 & ~n174 ;
  assign n176 = x13 ^ x1 ;
  assign n177 = n176 ^ x10 ;
  assign n178 = n177 ^ x13 ;
  assign n185 = n178 ^ n176 ;
  assign n186 = n185 ^ x13 ;
  assign n187 = n186 ^ x13 ;
  assign n38 = x7 & ~x14 ;
  assign n87 = ~x4 & ~x6 ;
  assign n88 = ~x5 & n87 ;
  assign n188 = n38 & n88 ;
  assign n189 = n131 & n188 ;
  assign n190 = n189 ^ n176 ;
  assign n191 = n190 ^ n176 ;
  assign n192 = n191 ^ x13 ;
  assign n193 = n187 & ~n192 ;
  assign n179 = x13 & ~x14 ;
  assign n180 = ~x11 & n179 ;
  assign n181 = n180 ^ n176 ;
  assign n182 = n181 ^ n178 ;
  assign n183 = n182 ^ x13 ;
  assign n184 = n178 & ~n183 ;
  assign n194 = n193 ^ n184 ;
  assign n195 = n194 ^ n178 ;
  assign n196 = n184 ^ x13 ;
  assign n197 = n196 ^ n186 ;
  assign n198 = x13 & n197 ;
  assign n199 = n198 ^ n184 ;
  assign n200 = n195 & n199 ;
  assign n201 = n200 ^ n193 ;
  assign n202 = n201 ^ n198 ;
  assign n203 = n202 ^ n178 ;
  assign n204 = n203 ^ x13 ;
  assign n205 = n204 ^ n186 ;
  assign n206 = n205 ^ x1 ;
  assign n207 = ~n175 & n206 ;
  assign n208 = ~x9 & ~n207 ;
  assign n209 = x7 & ~n117 ;
  assign n210 = ~n106 & ~n209 ;
  assign n211 = ~x11 & n166 ;
  assign n212 = ~n210 & n211 ;
  assign n213 = n212 ^ x10 ;
  assign n214 = n213 ^ n212 ;
  assign n215 = n214 ^ n208 ;
  assign n216 = ~x13 & ~x14 ;
  assign n217 = x0 & n216 ;
  assign n218 = n217 ^ x13 ;
  assign n219 = n218 ^ x11 ;
  assign n220 = n218 & n219 ;
  assign n221 = n220 ^ n212 ;
  assign n222 = n221 ^ n218 ;
  assign n223 = n215 & n222 ;
  assign n224 = n223 ^ n220 ;
  assign n225 = n224 ^ n218 ;
  assign n226 = ~n208 & n225 ;
  assign n227 = n226 ^ n208 ;
  assign n228 = ~n162 & ~n227 ;
  assign n37 = ~x10 & ~x11 ;
  assign n39 = x4 & ~x9 ;
  assign n40 = ~n38 & ~n39 ;
  assign n41 = n37 & ~n40 ;
  assign n43 = x7 & ~x8 ;
  assign n44 = ~x7 & x8 ;
  assign n45 = ~x5 & n44 ;
  assign n46 = ~n43 & ~n45 ;
  assign n47 = ~x3 & n46 ;
  assign n48 = x11 & ~n47 ;
  assign n49 = ~n42 & ~n48 ;
  assign n50 = n44 ^ x14 ;
  assign n51 = n50 ^ x14 ;
  assign n52 = x14 ^ x6 ;
  assign n53 = n52 ^ x14 ;
  assign n54 = n51 & n53 ;
  assign n55 = n54 ^ x14 ;
  assign n56 = x13 & ~n55 ;
  assign n57 = n56 ^ x14 ;
  assign n58 = n49 & n57 ;
  assign n59 = x9 & ~n58 ;
  assign n60 = n59 ^ x10 ;
  assign n61 = n60 ^ n59 ;
  assign n63 = ~x0 & ~n62 ;
  assign n64 = ~x2 & x5 ;
  assign n69 = n68 ^ n64 ;
  assign n70 = n69 ^ n64 ;
  assign n65 = n64 ^ x14 ;
  assign n66 = n65 ^ n64 ;
  assign n71 = n70 ^ n66 ;
  assign n72 = n64 ^ x1 ;
  assign n73 = n72 ^ n64 ;
  assign n74 = n73 ^ n70 ;
  assign n75 = n70 & n74 ;
  assign n76 = n75 ^ n70 ;
  assign n77 = ~n71 & n76 ;
  assign n78 = n77 ^ n75 ;
  assign n79 = n78 ^ n64 ;
  assign n80 = n79 ^ n70 ;
  assign n81 = x13 & n80 ;
  assign n82 = n81 ^ n64 ;
  assign n83 = n63 & n82 ;
  assign n84 = ~n23 & ~n83 ;
  assign n85 = ~x9 & x11 ;
  assign n86 = ~n84 & n85 ;
  assign n89 = x8 ^ x7 ;
  assign n92 = n91 ^ x8 ;
  assign n93 = n92 ^ n91 ;
  assign n95 = n94 ^ n91 ;
  assign n96 = ~n93 & n95 ;
  assign n97 = n96 ^ n91 ;
  assign n98 = n89 & n97 ;
  assign n99 = n88 & n98 ;
  assign n100 = x14 & n99 ;
  assign n101 = ~n86 & ~n100 ;
  assign n102 = n101 ^ n59 ;
  assign n103 = n61 & ~n102 ;
  assign n104 = n103 ^ n59 ;
  assign n105 = ~n41 & ~n104 ;
  assign n229 = n228 ^ n105 ;
  assign n230 = x12 & n229 ;
  assign n231 = n230 ^ n228 ;
  assign n232 = n36 & n231 ;
  assign y0 = ~n232 ;
endmodule
