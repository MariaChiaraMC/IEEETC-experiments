module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n13 = ~x0 & ~x3 ;
  assign n14 = ~x6 & n13 ;
  assign n15 = ~x4 & n14 ;
  assign n16 = x10 ^ x9 ;
  assign n17 = n16 ^ x11 ;
  assign n18 = n17 ^ x8 ;
  assign n19 = ~x1 & ~x2 ;
  assign n20 = x5 & x7 ;
  assign n21 = n19 & n20 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = x11 ^ x10 ;
  assign n24 = x10 ^ x8 ;
  assign n25 = n23 & n24 ;
  assign n26 = n25 ^ x10 ;
  assign n27 = n26 ^ n18 ;
  assign n28 = n22 & ~n27 ;
  assign n29 = n28 ^ n25 ;
  assign n30 = n29 ^ x10 ;
  assign n31 = n30 ^ n21 ;
  assign n32 = n18 & ~n31 ;
  assign n33 = n32 ^ n18 ;
  assign n34 = n15 & n33 ;
  assign y0 = n34 ;
endmodule
