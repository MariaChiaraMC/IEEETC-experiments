module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 ;
  assign n13 = x5 & x10 ;
  assign n14 = x7 & ~n13 ;
  assign n15 = ~x4 & x7 ;
  assign n16 = ~x6 & ~x11 ;
  assign n17 = ~n15 & ~n16 ;
  assign n18 = ~n14 & n17 ;
  assign n19 = x9 ^ x8 ;
  assign n20 = x6 & x11 ;
  assign n21 = x4 & n20 ;
  assign n22 = n21 ^ x9 ;
  assign n23 = x8 ^ x5 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n21 & ~n24 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = n22 & n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n28 ^ n21 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = ~n19 & ~n30 ;
  assign n32 = n31 ^ x8 ;
  assign n33 = ~n18 & ~n32 ;
  assign n34 = x5 & x9 ;
  assign n35 = x4 & ~n34 ;
  assign n36 = ~x8 & ~n35 ;
  assign n37 = x0 & ~n36 ;
  assign n43 = x7 ^ x2 ;
  assign n44 = x4 ^ x2 ;
  assign n45 = ~n43 & n44 ;
  assign n38 = x6 ^ x2 ;
  assign n47 = n45 ^ n38 ;
  assign n39 = n38 ^ x2 ;
  assign n40 = x8 ^ x2 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = ~n39 & ~n41 ;
  assign n48 = n42 ^ n38 ;
  assign n49 = n48 ^ n39 ;
  assign n50 = n49 ^ x1 ;
  assign n51 = ~n47 & n50 ;
  assign n46 = n45 ^ n42 ;
  assign n52 = n51 ^ n46 ;
  assign n53 = x1 & n52 ;
  assign n54 = n53 ^ n42 ;
  assign n55 = n54 ^ n45 ;
  assign n56 = n55 ^ n51 ;
  assign n57 = n56 ^ x1 ;
  assign n58 = n57 ^ x1 ;
  assign n59 = n37 & n58 ;
  assign n60 = x4 & x7 ;
  assign n61 = x2 & ~n60 ;
  assign n62 = ~x3 & ~n61 ;
  assign n63 = n59 & ~n62 ;
  assign n64 = n33 & n63 ;
  assign y0 = n64 ;
endmodule
