module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 ;
  assign n12 = ~x4 & x10 ;
  assign n13 = x6 ^ x3 ;
  assign n14 = n13 ^ x6 ;
  assign n15 = x7 ^ x6 ;
  assign n16 = ~n14 & n15 ;
  assign n17 = n16 ^ x6 ;
  assign n18 = ~x2 & ~x6 ;
  assign n19 = n18 ^ n12 ;
  assign n20 = ~n17 & n19 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n12 & n21 ;
  assign n23 = n22 ^ n12 ;
  assign n24 = n23 ^ x0 ;
  assign n25 = x3 & x7 ;
  assign n26 = x1 & x6 ;
  assign n27 = ~x8 & x9 ;
  assign n28 = ~n26 & n27 ;
  assign n29 = ~n25 & n28 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = x3 & ~n27 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = ~n31 & n33 ;
  assign n35 = n34 ^ n29 ;
  assign n36 = n35 ^ n23 ;
  assign n37 = ~n24 & n36 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = n38 ^ n29 ;
  assign n40 = n39 ^ x0 ;
  assign n41 = n23 & ~n40 ;
  assign n42 = n41 ^ n23 ;
  assign y0 = n42 ;
endmodule
