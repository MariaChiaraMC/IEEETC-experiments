// Benchmark "./apla.pla" written by ABC on Thu Apr 23 10:59:47 2020

module \./apla.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9,
    z5  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
  output z5;
  assign z5 = 1'b1;
endmodule


