module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 ;
  assign n25 = x0 & ~x1 ;
  assign n26 = ~x2 & ~x3 ;
  assign n27 = ~x0 & n26 ;
  assign n28 = ~n25 & ~n27 ;
  assign n29 = ~x1 & n26 ;
  assign n30 = ~x4 & x5 ;
  assign n31 = ~n29 & n30 ;
  assign n32 = ~n28 & n31 ;
  assign n33 = x20 ^ x18 ;
  assign n34 = n33 ^ x18 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = x0 & x2 ;
  assign n37 = x3 & ~x5 ;
  assign n38 = x4 & n37 ;
  assign n39 = x23 & n38 ;
  assign n40 = n36 & n39 ;
  assign n47 = ~x11 & ~x15 ;
  assign n48 = x12 & x13 ;
  assign n49 = n47 & n48 ;
  assign n50 = ~x10 & x11 ;
  assign n42 = x9 & x10 ;
  assign n51 = ~x6 & ~x7 ;
  assign n52 = ~n42 & n51 ;
  assign n53 = ~n50 & n52 ;
  assign n54 = n53 ^ x13 ;
  assign n55 = n54 ^ n53 ;
  assign n56 = ~x9 & ~x10 ;
  assign n57 = x7 & x16 ;
  assign n58 = n56 & n57 ;
  assign n59 = n58 ^ n53 ;
  assign n60 = n55 & n59 ;
  assign n61 = n60 ^ n53 ;
  assign n62 = ~x12 & n61 ;
  assign n63 = n62 ^ x11 ;
  assign n64 = ~x9 & x15 ;
  assign n65 = ~x13 & ~n56 ;
  assign n66 = ~n64 & n65 ;
  assign n67 = n66 ^ n62 ;
  assign n68 = n67 ^ n66 ;
  assign n69 = n68 ^ n63 ;
  assign n70 = x6 & x7 ;
  assign n71 = n70 ^ x9 ;
  assign n72 = x9 & n71 ;
  assign n73 = n72 ^ n66 ;
  assign n74 = n73 ^ x9 ;
  assign n75 = ~n69 & ~n74 ;
  assign n76 = n75 ^ n72 ;
  assign n77 = n76 ^ x9 ;
  assign n78 = n63 & n77 ;
  assign n79 = n78 ^ n62 ;
  assign n80 = ~n49 & ~n79 ;
  assign n81 = ~x8 & ~n80 ;
  assign n82 = x8 & n42 ;
  assign n83 = n70 & n82 ;
  assign n84 = ~x17 & ~n83 ;
  assign n85 = ~x1 & n84 ;
  assign n43 = x11 & n42 ;
  assign n86 = ~n43 & ~n82 ;
  assign n87 = ~x15 & ~n86 ;
  assign n88 = x8 & n51 ;
  assign n89 = x11 & ~x15 ;
  assign n90 = ~x9 & x10 ;
  assign n91 = x16 & n90 ;
  assign n92 = ~x13 & n91 ;
  assign n93 = ~n89 & ~n92 ;
  assign n94 = n88 & ~n93 ;
  assign n95 = ~n87 & ~n94 ;
  assign n96 = ~x12 & ~n95 ;
  assign n97 = n96 ^ n85 ;
  assign n98 = ~x12 & ~n89 ;
  assign n99 = ~x6 & ~x16 ;
  assign n100 = ~n98 & n99 ;
  assign n101 = n100 ^ x12 ;
  assign n102 = n101 ^ x7 ;
  assign n109 = n102 ^ n101 ;
  assign n103 = n102 ^ x9 ;
  assign n104 = n103 ^ n101 ;
  assign n105 = n102 ^ n100 ;
  assign n106 = n105 ^ x9 ;
  assign n107 = n106 ^ n104 ;
  assign n108 = n104 & n107 ;
  assign n110 = n109 ^ n108 ;
  assign n111 = n110 ^ n104 ;
  assign n112 = x8 & x10 ;
  assign n113 = x11 & n112 ;
  assign n114 = n113 ^ n101 ;
  assign n115 = n108 ^ n104 ;
  assign n116 = n114 & n115 ;
  assign n117 = n116 ^ n101 ;
  assign n118 = ~n111 & n117 ;
  assign n119 = n118 ^ n101 ;
  assign n120 = n119 ^ x12 ;
  assign n121 = n120 ^ n101 ;
  assign n122 = n121 ^ x13 ;
  assign n123 = n122 ^ n121 ;
  assign n124 = ~x8 & x11 ;
  assign n125 = n56 & n124 ;
  assign n126 = x16 & n125 ;
  assign n127 = x15 ^ x12 ;
  assign n128 = x9 & ~x10 ;
  assign n129 = n128 ^ n47 ;
  assign n130 = ~n127 & n129 ;
  assign n131 = n130 ^ n128 ;
  assign n132 = n47 & n131 ;
  assign n133 = n132 ^ x15 ;
  assign n134 = ~n126 & ~n133 ;
  assign n135 = ~x6 & ~n134 ;
  assign n136 = n135 ^ n121 ;
  assign n137 = n123 & ~n136 ;
  assign n138 = n137 ^ n121 ;
  assign n139 = n138 ^ n85 ;
  assign n140 = ~n97 & ~n139 ;
  assign n141 = n140 ^ n137 ;
  assign n142 = n141 ^ n121 ;
  assign n143 = n142 ^ n96 ;
  assign n144 = n85 & n143 ;
  assign n145 = n144 ^ n85 ;
  assign n146 = ~n81 & n145 ;
  assign n41 = x0 & x15 ;
  assign n44 = ~x12 & n43 ;
  assign n45 = ~x13 & ~n44 ;
  assign n46 = n41 & ~n45 ;
  assign n147 = n146 ^ n46 ;
  assign n148 = n147 ^ n46 ;
  assign n149 = x0 & x16 ;
  assign n150 = ~n25 & ~n149 ;
  assign n151 = n150 ^ n46 ;
  assign n152 = n151 ^ n46 ;
  assign n153 = ~n148 & n152 ;
  assign n154 = n153 ^ n46 ;
  assign n155 = x2 & n154 ;
  assign n156 = n155 ^ n46 ;
  assign n157 = n156 ^ x4 ;
  assign n158 = n157 ^ n156 ;
  assign n159 = n158 ^ x3 ;
  assign n160 = n36 ^ x22 ;
  assign n161 = n36 & ~n160 ;
  assign n162 = n161 ^ n156 ;
  assign n163 = n162 ^ n36 ;
  assign n164 = n159 & n163 ;
  assign n165 = n164 ^ n161 ;
  assign n166 = n165 ^ n36 ;
  assign n167 = ~x3 & n166 ;
  assign n168 = n167 ^ x3 ;
  assign n169 = n168 ^ x2 ;
  assign n170 = ~x1 & ~x4 ;
  assign n171 = ~x8 & n51 ;
  assign n172 = ~n82 & ~n171 ;
  assign n173 = ~x12 & ~x13 ;
  assign n174 = ~x11 & n173 ;
  assign n175 = ~n56 & n174 ;
  assign n176 = ~n172 & n175 ;
  assign n177 = ~x12 & n51 ;
  assign n178 = ~x13 & ~n177 ;
  assign n179 = n125 & ~n178 ;
  assign n180 = ~n176 & ~n179 ;
  assign n181 = n170 & ~n180 ;
  assign n182 = x3 & ~n181 ;
  assign n183 = n182 ^ n169 ;
  assign n184 = n183 ^ n168 ;
  assign n185 = n184 ^ n183 ;
  assign n186 = ~x0 & n170 ;
  assign n187 = n186 ^ n183 ;
  assign n188 = n187 ^ n169 ;
  assign n189 = n185 & n188 ;
  assign n190 = n189 ^ n186 ;
  assign n191 = n125 & n177 ;
  assign n192 = ~x4 & n41 ;
  assign n193 = ~x13 & n192 ;
  assign n194 = n191 & n193 ;
  assign n195 = x15 ^ x0 ;
  assign n196 = n195 ^ x15 ;
  assign n197 = x21 ^ x15 ;
  assign n198 = n196 & ~n197 ;
  assign n199 = n198 ^ x15 ;
  assign n200 = ~x1 & ~n199 ;
  assign n201 = ~n194 & ~n200 ;
  assign n202 = ~n186 & n201 ;
  assign n203 = n202 ^ n169 ;
  assign n204 = ~n190 & n203 ;
  assign n205 = n204 ^ n202 ;
  assign n206 = n169 & n205 ;
  assign n207 = n206 ^ n189 ;
  assign n208 = n207 ^ x2 ;
  assign n209 = n208 ^ n186 ;
  assign n210 = x5 & n209 ;
  assign n213 = n174 ^ n37 ;
  assign n214 = n213 ^ n37 ;
  assign n211 = n171 ^ n37 ;
  assign n212 = n211 ^ n37 ;
  assign n215 = n214 ^ n212 ;
  assign n216 = ~x3 & n90 ;
  assign n217 = n216 ^ n37 ;
  assign n218 = n217 ^ n37 ;
  assign n219 = n218 ^ n214 ;
  assign n220 = n214 & n219 ;
  assign n221 = n220 ^ n214 ;
  assign n222 = n215 & n221 ;
  assign n223 = n222 ^ n220 ;
  assign n224 = n223 ^ n37 ;
  assign n225 = n224 ^ n214 ;
  assign n226 = ~x4 & n225 ;
  assign n227 = n226 ^ n37 ;
  assign n230 = n227 ^ x3 ;
  assign n231 = n230 ^ n227 ;
  assign n228 = n227 ^ x4 ;
  assign n229 = n228 ^ n227 ;
  assign n232 = n231 ^ n229 ;
  assign n233 = x5 & ~x15 ;
  assign n234 = n233 ^ n227 ;
  assign n235 = n234 ^ n227 ;
  assign n236 = n235 ^ n231 ;
  assign n237 = ~n231 & n236 ;
  assign n238 = n237 ^ n231 ;
  assign n239 = ~n232 & ~n238 ;
  assign n240 = n239 ^ n237 ;
  assign n241 = n240 ^ n227 ;
  assign n242 = n241 ^ n231 ;
  assign n243 = ~x2 & ~n242 ;
  assign n244 = n243 ^ n227 ;
  assign n245 = n25 & n244 ;
  assign n246 = ~x4 & ~x22 ;
  assign n247 = x23 & n246 ;
  assign n248 = n29 & n247 ;
  assign n249 = ~n112 & ~n171 ;
  assign n250 = ~x3 & ~x5 ;
  assign n251 = x1 & x2 ;
  assign n252 = n250 & n251 ;
  assign n253 = ~x1 & x3 ;
  assign n254 = ~x2 & n253 ;
  assign n255 = ~n252 & ~n254 ;
  assign n256 = ~x11 & ~n255 ;
  assign n257 = ~n249 & n256 ;
  assign n258 = ~x15 & n252 ;
  assign n259 = ~n253 & ~n258 ;
  assign n260 = n88 & ~n259 ;
  assign n261 = n50 & n260 ;
  assign n262 = ~n257 & ~n261 ;
  assign n263 = x9 & n173 ;
  assign n264 = ~x4 & n263 ;
  assign n265 = ~n262 & n264 ;
  assign n266 = x1 & n38 ;
  assign n267 = ~x2 & n266 ;
  assign n268 = ~n265 & ~n267 ;
  assign n269 = ~n248 & n268 ;
  assign n270 = ~x0 & ~n269 ;
  assign n271 = ~n245 & ~n270 ;
  assign n272 = ~n210 & n271 ;
  assign n273 = ~n40 & n272 ;
  assign n274 = n273 ^ x19 ;
  assign n275 = ~n273 & n274 ;
  assign n276 = n275 ^ x18 ;
  assign n277 = n276 ^ n273 ;
  assign n278 = n35 & n277 ;
  assign n279 = n278 ^ n275 ;
  assign n280 = n279 ^ n273 ;
  assign n281 = ~n32 & ~n280 ;
  assign n282 = n281 ^ n32 ;
  assign n283 = x14 & n282 ;
  assign y0 = n283 ;
endmodule
