module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 ;
  assign n13 = ~x7 & ~x8 ;
  assign n14 = ~x4 & n13 ;
  assign n10 = x7 & x8 ;
  assign n11 = ~x6 & x7 ;
  assign n12 = ~n10 & ~n11 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = x3 & ~n15 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = x2 & n17 ;
  assign n19 = ~x2 & ~x3 ;
  assign n20 = ~x4 & x7 ;
  assign n21 = n19 & n20 ;
  assign n22 = ~x8 & n21 ;
  assign n23 = ~n18 & ~n22 ;
  assign n24 = ~x5 & ~n23 ;
  assign n25 = x2 & x7 ;
  assign n26 = x5 & x6 ;
  assign n27 = x4 & n26 ;
  assign n28 = n27 ^ x4 ;
  assign n29 = ~x3 & ~n28 ;
  assign n30 = n29 ^ x4 ;
  assign n31 = n25 & ~n30 ;
  assign n32 = ~n24 & ~n31 ;
  assign n33 = ~x8 & n25 ;
  assign n34 = ~x4 & ~n26 ;
  assign n35 = ~n33 & n34 ;
  assign n36 = x8 ^ x3 ;
  assign n38 = x7 ^ x2 ;
  assign n37 = n36 ^ x8 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = n38 ^ x2 ;
  assign n41 = n40 ^ n36 ;
  assign n42 = n39 & n41 ;
  assign n43 = n42 ^ x2 ;
  assign n44 = x2 & ~x4 ;
  assign n45 = n44 ^ n36 ;
  assign n46 = n43 & ~n45 ;
  assign n47 = n46 ^ n44 ;
  assign n48 = ~n36 & n47 ;
  assign n49 = n48 ^ n42 ;
  assign n50 = n49 ^ x2 ;
  assign n51 = ~n35 & n50 ;
  assign n52 = ~x2 & x3 ;
  assign n53 = ~x5 & ~x6 ;
  assign n54 = ~x8 & n53 ;
  assign n55 = n52 & ~n54 ;
  assign n56 = ~x7 & n55 ;
  assign n57 = ~n51 & ~n56 ;
  assign n58 = n57 ^ x1 ;
  assign n59 = n58 ^ n57 ;
  assign n60 = n11 & n52 ;
  assign n61 = x8 ^ x2 ;
  assign n62 = n61 ^ n53 ;
  assign n63 = x7 ^ x3 ;
  assign n64 = n38 ^ x7 ;
  assign n65 = ~n63 & ~n64 ;
  assign n66 = n65 ^ x7 ;
  assign n67 = n66 ^ n61 ;
  assign n68 = n62 & n67 ;
  assign n69 = n68 ^ n65 ;
  assign n70 = n69 ^ x7 ;
  assign n71 = n70 ^ n53 ;
  assign n72 = ~n61 & n71 ;
  assign n73 = n72 ^ n61 ;
  assign n74 = ~n60 & n73 ;
  assign n75 = x4 & ~n74 ;
  assign n76 = x3 & ~x4 ;
  assign n77 = x5 & x7 ;
  assign n78 = n76 & n77 ;
  assign n79 = x3 & x8 ;
  assign n80 = ~x3 & n14 ;
  assign n81 = ~n79 & ~n80 ;
  assign n82 = ~n52 & ~n81 ;
  assign n83 = ~n78 & ~n82 ;
  assign n84 = ~n75 & n83 ;
  assign n85 = n10 & n27 ;
  assign n86 = x2 & n13 ;
  assign n87 = ~n85 & ~n86 ;
  assign n88 = n87 ^ x5 ;
  assign n89 = n88 ^ x3 ;
  assign n98 = n89 ^ n88 ;
  assign n90 = ~x6 & ~x8 ;
  assign n91 = n44 & n90 ;
  assign n92 = n91 ^ n89 ;
  assign n93 = n92 ^ n88 ;
  assign n94 = n89 ^ n87 ;
  assign n95 = n94 ^ n91 ;
  assign n96 = n95 ^ n93 ;
  assign n97 = n93 & n96 ;
  assign n99 = n98 ^ n97 ;
  assign n100 = n99 ^ n93 ;
  assign n101 = n88 ^ n10 ;
  assign n102 = n97 ^ n93 ;
  assign n103 = ~n101 & n102 ;
  assign n104 = n103 ^ n88 ;
  assign n105 = ~n100 & n104 ;
  assign n106 = n105 ^ n88 ;
  assign n107 = n106 ^ x5 ;
  assign n108 = n107 ^ n88 ;
  assign n109 = n84 & n108 ;
  assign n110 = n109 ^ n57 ;
  assign n111 = n59 & n110 ;
  assign n112 = n111 ^ n57 ;
  assign n113 = n32 & n112 ;
  assign n114 = ~x0 & ~n113 ;
  assign n115 = n19 & ~n20 ;
  assign n116 = ~n10 & ~n13 ;
  assign n117 = n115 & n116 ;
  assign n118 = n117 ^ n22 ;
  assign n119 = n117 ^ x0 ;
  assign n120 = n119 ^ n118 ;
  assign n121 = x7 ^ x4 ;
  assign n122 = x5 & ~n121 ;
  assign n123 = n122 ^ x4 ;
  assign n124 = n123 ^ n26 ;
  assign n125 = x0 & n124 ;
  assign n126 = n125 ^ n123 ;
  assign n127 = n120 & n126 ;
  assign n128 = n127 ^ n125 ;
  assign n129 = n128 ^ n123 ;
  assign n130 = n129 ^ x0 ;
  assign n131 = n118 & n130 ;
  assign n132 = n131 ^ n22 ;
  assign n133 = ~x1 & n132 ;
  assign n134 = ~n114 & ~n133 ;
  assign y0 = ~n134 ;
endmodule
