// Benchmark "./pla/mish.pla_dbb_orig_0NonExact" written by ABC on Fri Nov 20 10:25:31 2020

module \./pla/mish.pla_dbb_orig_0NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = ~x0;
endmodule


