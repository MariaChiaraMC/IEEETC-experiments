module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 ;
  assign n9 = ~x0 & ~x1 ;
  assign n10 = ~x3 & ~x4 ;
  assign n11 = ~x2 & ~n10 ;
  assign n12 = n9 & ~n11 ;
  assign n13 = x6 & ~n12 ;
  assign n14 = x5 & ~x7 ;
  assign n15 = n9 ^ x4 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = x3 ^ x2 ;
  assign n18 = ~x4 & n17 ;
  assign n19 = n18 ^ x3 ;
  assign n20 = ~n16 & ~n19 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n21 ^ x3 ;
  assign n23 = n22 ^ x4 ;
  assign n24 = n14 & n23 ;
  assign n25 = n13 & n24 ;
  assign y0 = n25 ;
endmodule
