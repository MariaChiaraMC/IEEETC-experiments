module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n9 = x2 ^ x1 ;
  assign n10 = n9 ^ x2 ;
  assign n11 = x5 & x6 ;
  assign n12 = ~x4 & ~n11 ;
  assign n13 = ~x2 & ~n12 ;
  assign n14 = n13 ^ x4 ;
  assign n15 = ~x3 & ~n14 ;
  assign n16 = ~x5 & ~x6 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = ~x2 & ~x7 ;
  assign n19 = ~n13 & ~n18 ;
  assign n20 = n19 ^ n15 ;
  assign n21 = ~n17 & n20 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n15 & n22 ;
  assign n24 = n23 ^ n13 ;
  assign n25 = n24 ^ x2 ;
  assign n26 = ~n10 & n25 ;
  assign n27 = n26 ^ x2 ;
  assign n28 = ~x0 & ~n27 ;
  assign y0 = n28 ;
endmodule
