module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n9 = ~x2 & x7 ;
  assign n10 = ~x5 & n9 ;
  assign n11 = ~x4 & ~n10 ;
  assign n12 = ~x3 & ~n11 ;
  assign n13 = ~x0 & ~x1 ;
  assign n14 = x3 ^ x2 ;
  assign n15 = x5 ^ x3 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = ~x6 & ~x7 ;
  assign n18 = ~x4 & n17 ;
  assign n19 = n18 ^ x6 ;
  assign n20 = ~x3 & n19 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n16 & n21 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n23 ^ n18 ;
  assign n25 = n24 ^ x3 ;
  assign n26 = n14 & ~n25 ;
  assign n27 = n26 ^ x2 ;
  assign n28 = n13 & ~n27 ;
  assign n29 = ~n12 & n28 ;
  assign y0 = n29 ;
endmodule
