module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 ;
  assign n17 = ~x6 & ~x7 ;
  assign n18 = ~x0 & x5 ;
  assign n19 = x4 & n18 ;
  assign n20 = ~n17 & n19 ;
  assign n21 = x3 & ~n20 ;
  assign n22 = x1 ^ x0 ;
  assign n23 = x7 ^ x1 ;
  assign n24 = n23 ^ x7 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = x7 ^ x6 ;
  assign n27 = x7 ^ x4 ;
  assign n28 = x7 ^ x5 ;
  assign n29 = ~x7 & ~n28 ;
  assign n30 = n29 ^ x7 ;
  assign n31 = ~n27 & ~n30 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = n32 ^ x7 ;
  assign n34 = n33 ^ x5 ;
  assign n35 = ~n26 & ~n34 ;
  assign n36 = n35 ^ x7 ;
  assign n37 = x14 & x15 ;
  assign n38 = x9 & ~n37 ;
  assign n39 = ~x10 & ~x11 ;
  assign n40 = ~x8 & ~x12 ;
  assign n41 = n39 & n40 ;
  assign n42 = n38 & n41 ;
  assign n43 = ~x14 & ~x15 ;
  assign n44 = n43 ^ x13 ;
  assign n45 = n42 & ~n44 ;
  assign n46 = ~n36 & n45 ;
  assign n47 = ~x3 & ~n46 ;
  assign n48 = n47 ^ x2 ;
  assign n49 = ~x2 & n48 ;
  assign n50 = n49 ^ x7 ;
  assign n51 = n50 ^ x2 ;
  assign n52 = n25 & ~n51 ;
  assign n53 = n52 ^ n49 ;
  assign n54 = n53 ^ x2 ;
  assign n55 = n22 & ~n54 ;
  assign n56 = ~n21 & n55 ;
  assign y0 = n56 ;
endmodule
