module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 ;
  assign n15 = ~x11 & ~x12 ;
  assign n16 = ~x10 & n15 ;
  assign n17 = ~x9 & n16 ;
  assign n18 = ~x8 & n17 ;
  assign n19 = ~x7 & n18 ;
  assign n20 = ~x6 & n19 ;
  assign n58 = ~x5 & n20 ;
  assign n59 = ~x4 & n58 ;
  assign n60 = n59 ^ x3 ;
  assign n21 = n16 ^ x7 ;
  assign n22 = n16 ^ x9 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = x11 & x12 ;
  assign n26 = n25 ^ x8 ;
  assign n27 = ~n16 & n26 ;
  assign n28 = n27 ^ x8 ;
  assign n29 = n24 & ~n28 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n30 ^ x8 ;
  assign n32 = n31 ^ n16 ;
  assign n33 = ~n21 & n32 ;
  assign n34 = n33 ^ x7 ;
  assign n35 = ~x5 & ~n34 ;
  assign n36 = ~n20 & ~n35 ;
  assign n37 = ~x0 & ~n36 ;
  assign n38 = n19 ^ x4 ;
  assign n39 = n19 ^ x6 ;
  assign n40 = n39 ^ n19 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = x10 & ~n15 ;
  assign n43 = ~x8 & ~n42 ;
  assign n44 = ~n17 & ~n43 ;
  assign n45 = n44 ^ x5 ;
  assign n46 = ~n19 & n45 ;
  assign n47 = n46 ^ x5 ;
  assign n48 = n41 & ~n47 ;
  assign n49 = n48 ^ n46 ;
  assign n50 = n49 ^ x5 ;
  assign n51 = n50 ^ n19 ;
  assign n52 = ~n38 & n51 ;
  assign n53 = n52 ^ x4 ;
  assign n54 = n37 & ~n53 ;
  assign n55 = n54 ^ x2 ;
  assign n56 = n55 ^ x1 ;
  assign n57 = n56 ^ x3 ;
  assign n61 = n60 ^ n57 ;
  assign n64 = n56 ^ x1 ;
  assign n62 = x2 ^ x1 ;
  assign n63 = n62 ^ n57 ;
  assign n65 = n64 ^ n63 ;
  assign n66 = n61 & n65 ;
  assign n67 = n66 ^ n56 ;
  assign n68 = n67 ^ n62 ;
  assign n69 = n68 ^ n64 ;
  assign n70 = n63 ^ n60 ;
  assign n71 = n67 & n70 ;
  assign n72 = n71 ^ n56 ;
  assign n73 = n72 ^ n57 ;
  assign n74 = n73 ^ n60 ;
  assign n75 = ~n69 & n74 ;
  assign y0 = n75 ;
endmodule
