module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 ;
  assign n17 = ~x1 & ~x3 ;
  assign n18 = ~x4 & x6 ;
  assign n19 = n17 & n18 ;
  assign n20 = ~x10 & n19 ;
  assign n21 = x7 ^ x2 ;
  assign n22 = x8 ^ x7 ;
  assign n23 = x15 ^ x8 ;
  assign n24 = ~n22 & ~n23 ;
  assign n25 = n21 & n24 ;
  assign n26 = n20 & n25 ;
  assign n27 = x3 & x4 ;
  assign n28 = x1 & n27 ;
  assign n29 = x2 & ~x8 ;
  assign n30 = x7 & x10 ;
  assign n31 = x6 & ~n30 ;
  assign n32 = n29 & ~n31 ;
  assign n33 = n28 & n32 ;
  assign n34 = x15 & n33 ;
  assign n35 = ~n26 & ~n34 ;
  assign n36 = ~x14 & ~n35 ;
  assign n37 = x8 & x11 ;
  assign n38 = x10 & ~x15 ;
  assign n39 = x14 & n38 ;
  assign n40 = ~x2 & ~x7 ;
  assign n41 = n39 & n40 ;
  assign n42 = n37 & n41 ;
  assign n43 = n19 & n42 ;
  assign n44 = ~n36 & ~n43 ;
  assign n45 = ~x5 & ~n44 ;
  assign n46 = x6 & x10 ;
  assign n47 = ~x7 & ~n46 ;
  assign n48 = ~x14 & n29 ;
  assign n49 = n47 & n48 ;
  assign n50 = n28 & n49 ;
  assign n51 = x15 & n50 ;
  assign n52 = ~n45 & ~n51 ;
  assign n53 = x9 & ~n52 ;
  assign n54 = ~x1 & ~x7 ;
  assign n55 = n27 & n54 ;
  assign n56 = ~x6 & ~x9 ;
  assign n57 = x5 & n38 ;
  assign n58 = n56 & n57 ;
  assign n59 = n55 & n58 ;
  assign n60 = n48 & n59 ;
  assign n61 = ~n53 & ~n60 ;
  assign n62 = ~x12 & ~x13 ;
  assign n63 = ~x0 & n62 ;
  assign n64 = ~n61 & n63 ;
  assign y0 = n64 ;
endmodule
