module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 ;
  assign n9 = x2 ^ x1 ;
  assign n10 = n9 ^ x2 ;
  assign n11 = x4 ^ x3 ;
  assign n12 = n11 ^ x3 ;
  assign n13 = x5 ^ x3 ;
  assign n14 = n13 ^ n11 ;
  assign n15 = ~n12 & n14 ;
  assign n16 = n15 ^ n11 ;
  assign n17 = n16 ^ x2 ;
  assign n18 = x6 ^ x3 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = x7 & n19 ;
  assign n21 = n20 ^ x7 ;
  assign n22 = n21 ^ n13 ;
  assign n23 = n22 ^ n18 ;
  assign n24 = n23 ^ n12 ;
  assign n25 = n24 ^ x2 ;
  assign n26 = n19 ^ x2 ;
  assign n27 = n18 ^ n14 ;
  assign n28 = n27 ^ n12 ;
  assign n29 = n28 ^ x2 ;
  assign n30 = ~n26 & ~n29 ;
  assign n31 = n30 ^ n13 ;
  assign n32 = n31 ^ n18 ;
  assign n33 = n25 & n32 ;
  assign n34 = n33 ^ x2 ;
  assign n35 = n17 & ~n34 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = n36 ^ x2 ;
  assign n38 = n37 ^ x2 ;
  assign n39 = n38 ^ x2 ;
  assign n40 = ~n10 & n39 ;
  assign n41 = n40 ^ x2 ;
  assign n42 = ~x0 & ~n41 ;
  assign y0 = n42 ;
endmodule
