module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 ;
  assign n18 = ~x3 & ~x9 ;
  assign n19 = x2 & ~n18 ;
  assign n20 = x0 & x1 ;
  assign n21 = n20 ^ x15 ;
  assign n22 = n19 & n21 ;
  assign n23 = n22 ^ x15 ;
  assign n24 = x14 & n23 ;
  assign n134 = ~x6 & x15 ;
  assign n25 = ~x4 & ~x5 ;
  assign n26 = ~x16 & n25 ;
  assign n27 = n26 ^ x4 ;
  assign n28 = n27 ^ x8 ;
  assign n73 = n28 ^ n27 ;
  assign n29 = x2 & x5 ;
  assign n30 = x11 ^ x3 ;
  assign n31 = n30 ^ x10 ;
  assign n32 = n31 ^ x10 ;
  assign n33 = n32 ^ x11 ;
  assign n34 = x11 ^ x8 ;
  assign n35 = n33 & n34 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = n36 ^ x8 ;
  assign n38 = x11 ^ x9 ;
  assign n39 = n38 ^ n31 ;
  assign n40 = n39 ^ x10 ;
  assign n41 = n40 ^ n33 ;
  assign n42 = x10 ^ x8 ;
  assign n48 = n42 ^ x11 ;
  assign n49 = n41 ^ x8 ;
  assign n50 = n48 & n49 ;
  assign n43 = x12 ^ x11 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = n44 ^ x11 ;
  assign n46 = n45 ^ n40 ;
  assign n47 = n45 & ~n46 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = n51 ^ n43 ;
  assign n53 = n52 ^ n42 ;
  assign n54 = n53 ^ x11 ;
  assign n55 = n54 ^ n33 ;
  assign n56 = n55 ^ x8 ;
  assign n57 = ~n41 & ~n56 ;
  assign n58 = n57 ^ n50 ;
  assign n59 = n58 ^ n42 ;
  assign n60 = n59 ^ n33 ;
  assign n61 = n60 ^ n40 ;
  assign n62 = ~n37 & n61 ;
  assign n63 = n62 ^ n35 ;
  assign n64 = n63 ^ n33 ;
  assign n65 = n64 ^ x8 ;
  assign n66 = n29 & ~n65 ;
  assign n67 = n66 ^ n28 ;
  assign n68 = n67 ^ n27 ;
  assign n69 = n28 ^ n26 ;
  assign n70 = n69 ^ n66 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = ~n68 & ~n71 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = n74 ^ n68 ;
  assign n76 = x5 ^ x2 ;
  assign n77 = n76 ^ n18 ;
  assign n78 = n20 ^ x2 ;
  assign n79 = n78 ^ n20 ;
  assign n80 = x12 & x13 ;
  assign n81 = n80 ^ n20 ;
  assign n82 = ~n79 & n81 ;
  assign n83 = n82 ^ n20 ;
  assign n84 = n83 ^ n76 ;
  assign n85 = ~n77 & n84 ;
  assign n86 = n85 ^ n82 ;
  assign n87 = n86 ^ n20 ;
  assign n88 = n87 ^ n18 ;
  assign n89 = n76 & ~n88 ;
  assign n90 = n89 ^ n76 ;
  assign n91 = n90 ^ n27 ;
  assign n92 = n72 ^ n68 ;
  assign n93 = ~n91 & ~n92 ;
  assign n94 = n93 ^ n27 ;
  assign n95 = ~n75 & n94 ;
  assign n96 = n95 ^ n27 ;
  assign n97 = n96 ^ x4 ;
  assign n98 = n97 ^ n27 ;
  assign n99 = n98 ^ x6 ;
  assign n112 = n99 ^ x5 ;
  assign n100 = ~x8 & x15 ;
  assign n101 = n100 ^ n98 ;
  assign n102 = n101 ^ n99 ;
  assign n103 = n102 ^ n99 ;
  assign n111 = n103 ^ x5 ;
  assign n113 = n112 ^ n111 ;
  assign n105 = n102 ^ x4 ;
  assign n106 = n105 ^ n102 ;
  assign n104 = n103 ^ n98 ;
  assign n107 = n106 ^ n104 ;
  assign n108 = n104 ^ x5 ;
  assign n109 = n107 & n108 ;
  assign n110 = n109 ^ x5 ;
  assign n114 = n113 ^ n110 ;
  assign n115 = n114 ^ n106 ;
  assign n116 = n113 ^ n112 ;
  assign n117 = n116 ^ n104 ;
  assign n118 = n112 & ~n117 ;
  assign n119 = n112 ^ n106 ;
  assign n120 = ~n19 & n119 ;
  assign n121 = n120 ^ n19 ;
  assign n122 = n121 ^ n106 ;
  assign n123 = n122 ^ n104 ;
  assign n124 = n118 & ~n123 ;
  assign n125 = n124 ^ x5 ;
  assign n126 = ~n115 & n125 ;
  assign n127 = n126 ^ n118 ;
  assign n128 = n127 ^ n124 ;
  assign n129 = n128 ^ x5 ;
  assign n130 = n129 ^ n112 ;
  assign n131 = n130 ^ n113 ;
  assign n132 = n131 ^ x6 ;
  assign n133 = n132 ^ n103 ;
  assign n135 = n134 ^ n133 ;
  assign n136 = n135 ^ n133 ;
  assign n137 = n133 ^ n25 ;
  assign n138 = n137 ^ n133 ;
  assign n139 = n136 & n138 ;
  assign n140 = n139 ^ n133 ;
  assign n141 = ~x7 & n140 ;
  assign n142 = n141 ^ n133 ;
  assign n143 = ~n24 & ~n142 ;
  assign y0 = ~n143 ;
endmodule
