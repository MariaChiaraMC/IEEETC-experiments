module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 ;
  assign n13 = x0 & x9 ;
  assign n14 = x8 ^ x5 ;
  assign n16 = x2 & x3 ;
  assign n19 = x6 & x7 ;
  assign n20 = n16 & n19 ;
  assign n15 = ~x7 & ~x11 ;
  assign n17 = ~x6 & ~n16 ;
  assign n18 = n15 & n17 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n20 ^ x8 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n21 & n23 ;
  assign n25 = n24 ^ n20 ;
  assign n26 = x10 & ~x11 ;
  assign n27 = n20 & n26 ;
  assign n28 = n27 ^ n14 ;
  assign n29 = n25 & ~n28 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = ~n14 & n30 ;
  assign n32 = n31 ^ n14 ;
  assign n33 = n32 ^ n14 ;
  assign n36 = n33 ^ x3 ;
  assign n37 = n36 ^ n33 ;
  assign n34 = n33 ^ x2 ;
  assign n35 = n34 ^ n33 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = x5 & x8 ;
  assign n40 = n19 & n39 ;
  assign n41 = n40 ^ n33 ;
  assign n42 = n41 ^ n33 ;
  assign n43 = n42 ^ n37 ;
  assign n44 = ~n37 & ~n43 ;
  assign n45 = n44 ^ n37 ;
  assign n46 = ~n38 & ~n45 ;
  assign n47 = n46 ^ n44 ;
  assign n48 = n47 ^ n33 ;
  assign n49 = n48 ^ n37 ;
  assign n50 = ~x4 & ~n49 ;
  assign n51 = n50 ^ n33 ;
  assign n52 = n13 & n51 ;
  assign n53 = ~x1 & n52 ;
  assign y0 = n53 ;
endmodule
