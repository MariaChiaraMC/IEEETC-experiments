module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;
  assign n11 = ~x4 & ~x6 ;
  assign n17 = x8 & x9 ;
  assign n18 = x7 & n17 ;
  assign n12 = ~x8 & ~x9 ;
  assign n13 = x0 & x1 ;
  assign n14 = n12 & n13 ;
  assign n15 = ~x2 & x3 ;
  assign n16 = n14 & n15 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = n18 ^ x7 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = n20 & ~n22 ;
  assign n24 = n23 ^ n18 ;
  assign n25 = ~x5 & n24 ;
  assign n26 = n25 ^ n18 ;
  assign n27 = n11 & n26 ;
  assign n28 = n18 ^ x6 ;
  assign n29 = ~x5 & ~x7 ;
  assign n30 = ~n17 & n29 ;
  assign n31 = n30 ^ x4 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = n30 ^ x5 ;
  assign n34 = ~n32 & n33 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n35 ^ n18 ;
  assign n37 = ~n28 & ~n36 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = n38 ^ n30 ;
  assign n40 = n39 ^ x6 ;
  assign n41 = ~n18 & n40 ;
  assign n42 = n41 ^ n18 ;
  assign n43 = ~n27 & n42 ;
  assign y0 = ~n43 ;
endmodule
