module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n9 = x3 ^ x1 ;
  assign n10 = n9 ^ x1 ;
  assign n11 = x5 ^ x4 ;
  assign n12 = n11 ^ x6 ;
  assign n13 = x6 ^ x5 ;
  assign n14 = n13 ^ x6 ;
  assign n15 = x7 ^ x6 ;
  assign n16 = n14 & ~n15 ;
  assign n17 = n16 ^ x6 ;
  assign n18 = n12 & n17 ;
  assign n19 = ~x1 & n18 ;
  assign n20 = n19 ^ x1 ;
  assign n21 = ~n10 & ~n20 ;
  assign n22 = n21 ^ x1 ;
  assign n23 = ~x2 & n22 ;
  assign n24 = n23 ^ x3 ;
  assign y0 = ~n24 ;
endmodule
