// Benchmark "./pla/m1.pla_9" written by ABC on Mon Apr 20 15:44:07 2020

module \./pla/m1.pla_9  ( 
    x0, x1, x2, x3, x4, x5,
    z0  );
  input  x0, x1, x2, x3, x4, x5;
  output z0;
  wire new_n8_, new_n9_, new_n10_, new_n11_, new_n12_, new_n13_, new_n14_;
  assign new_n8_ = x4 & x5;
  assign new_n9_ = ~x2 & new_n8_;
  assign new_n10_ = ~x4 & ~x5;
  assign new_n11_ = x2 & ~x3;
  assign new_n12_ = ~new_n10_ & ~new_n11_;
  assign new_n13_ = ~new_n9_ & new_n12_;
  assign new_n14_ = ~x0 & ~x1;
  assign z0 = ~new_n13_ & new_n14_;
endmodule


