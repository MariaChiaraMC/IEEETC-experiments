module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n8 = x3 ^ x0 ;
  assign n9 = x4 ^ x1 ;
  assign n10 = n9 ^ x3 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = n9 ^ x2 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = n11 & ~n13 ;
  assign n15 = n14 ^ n9 ;
  assign n16 = n8 & ~n15 ;
  assign n17 = n16 ^ n9 ;
  assign n18 = x6 ^ x1 ;
  assign n19 = n18 ^ x0 ;
  assign n20 = n19 ^ x0 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = x0 & ~x3 ;
  assign n23 = x2 & n22 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = ~n23 & ~n24 ;
  assign n26 = n25 ^ x0 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = ~n21 & n27 ;
  assign n29 = n28 ^ n25 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = n17 & ~n30 ;
  assign n32 = n31 ^ n17 ;
  assign y0 = n32 ;
endmodule
