module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n18 = ~x4 & ~x5 ;
  assign n19 = ~x1 & n18 ;
  assign n20 = ~x8 & x9 ;
  assign n21 = ~n19 & n20 ;
  assign n11 = x8 ^ x1 ;
  assign n12 = x8 ^ x4 ;
  assign n13 = n12 ^ x8 ;
  assign n14 = ~n11 & ~n13 ;
  assign n15 = n14 ^ x8 ;
  assign n16 = ~x9 & ~n15 ;
  assign n17 = n16 ^ x8 ;
  assign n22 = n21 ^ n17 ;
  assign n23 = ~x7 & n22 ;
  assign n24 = n23 ^ n17 ;
  assign y0 = n24 ;
endmodule
