module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 ;
  assign n16 = x13 ^ x11 ;
  assign n17 = ~x3 & x8 ;
  assign n18 = ~x5 & x7 ;
  assign n19 = ~x6 & n18 ;
  assign n20 = ~x4 & n19 ;
  assign n21 = ~x9 & ~x14 ;
  assign n22 = n20 & n21 ;
  assign n23 = n17 & n22 ;
  assign n24 = x10 ^ x0 ;
  assign n25 = n24 ^ x14 ;
  assign n26 = ~x1 & ~x6 ;
  assign n27 = x4 & x5 ;
  assign n28 = n26 & n27 ;
  assign n29 = ~x9 & n28 ;
  assign n30 = n29 ^ x1 ;
  assign n31 = ~x10 & n30 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = n25 & n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n34 ^ n29 ;
  assign n36 = n35 ^ x10 ;
  assign n37 = x14 & ~n36 ;
  assign n38 = ~n23 & ~n37 ;
  assign n39 = n38 ^ x13 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = ~x3 & n21 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = n40 & ~n42 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = n16 & ~n44 ;
  assign n46 = ~x12 & n45 ;
  assign n47 = ~x7 & ~x8 ;
  assign n48 = ~x11 & ~x14 ;
  assign n49 = ~x6 & n48 ;
  assign n50 = ~n47 & n49 ;
  assign n51 = ~x7 & ~x13 ;
  assign n52 = ~x4 & x11 ;
  assign n53 = x3 & ~x8 ;
  assign n54 = n52 & ~n53 ;
  assign n55 = n54 ^ x6 ;
  assign n56 = n55 ^ n51 ;
  assign n57 = n48 ^ n17 ;
  assign n58 = n54 & ~n57 ;
  assign n59 = n58 ^ n48 ;
  assign n60 = n56 & n59 ;
  assign n61 = n60 ^ n58 ;
  assign n62 = n61 ^ n48 ;
  assign n63 = n62 ^ n54 ;
  assign n64 = n51 & n63 ;
  assign n65 = ~n50 & ~n64 ;
  assign n66 = ~x5 & ~x12 ;
  assign n67 = ~n65 & n66 ;
  assign n68 = n67 ^ x4 ;
  assign n69 = n68 ^ x9 ;
  assign n97 = n69 ^ n68 ;
  assign n70 = ~x11 & ~x12 ;
  assign n71 = x9 & ~x13 ;
  assign n72 = x14 & ~n71 ;
  assign n73 = n72 ^ x7 ;
  assign n74 = x7 ^ x5 ;
  assign n75 = n74 ^ n73 ;
  assign n76 = n72 ^ x13 ;
  assign n77 = n76 ^ x13 ;
  assign n78 = x9 & ~x14 ;
  assign n79 = n78 ^ x13 ;
  assign n80 = ~n77 & ~n79 ;
  assign n81 = n80 ^ x13 ;
  assign n82 = n81 ^ n73 ;
  assign n83 = ~n75 & ~n82 ;
  assign n84 = n83 ^ n80 ;
  assign n85 = n84 ^ x13 ;
  assign n86 = n85 ^ n74 ;
  assign n87 = ~n73 & n86 ;
  assign n88 = n87 ^ n73 ;
  assign n89 = n88 ^ n72 ;
  assign n90 = n70 & n89 ;
  assign n91 = n90 ^ n69 ;
  assign n92 = n91 ^ n68 ;
  assign n93 = n69 ^ n67 ;
  assign n94 = n93 ^ n90 ;
  assign n95 = n94 ^ n92 ;
  assign n96 = ~n92 & ~n95 ;
  assign n98 = n97 ^ n96 ;
  assign n99 = n98 ^ n92 ;
  assign n100 = x1 & n18 ;
  assign n101 = x12 & ~x14 ;
  assign n102 = x13 & n101 ;
  assign n103 = n100 & n102 ;
  assign n104 = ~x12 & ~x14 ;
  assign n105 = x5 & ~x13 ;
  assign n106 = ~n104 & n105 ;
  assign n107 = ~n26 & n106 ;
  assign n108 = ~n103 & ~n107 ;
  assign n109 = x11 & x13 ;
  assign n110 = ~x2 & x11 ;
  assign n111 = ~n109 & ~n110 ;
  assign n112 = x12 & n111 ;
  assign n113 = ~x3 & ~n112 ;
  assign n114 = ~n108 & n113 ;
  assign n115 = x5 & ~x7 ;
  assign n116 = n70 & ~n115 ;
  assign n117 = x13 & n116 ;
  assign n118 = ~n114 & ~n117 ;
  assign n119 = n118 ^ n68 ;
  assign n120 = n96 ^ n92 ;
  assign n121 = n119 & ~n120 ;
  assign n122 = n121 ^ n68 ;
  assign n123 = ~n99 & n122 ;
  assign n124 = n123 ^ n68 ;
  assign n125 = n124 ^ x4 ;
  assign n126 = n125 ^ n68 ;
  assign n127 = ~x0 & n126 ;
  assign n128 = x6 & n27 ;
  assign n129 = ~x12 & n128 ;
  assign n130 = x7 & n129 ;
  assign n131 = x4 & n100 ;
  assign n132 = n104 & ~n131 ;
  assign n133 = ~n130 & ~n132 ;
  assign n139 = n133 ^ x9 ;
  assign n148 = n139 ^ n133 ;
  assign n134 = ~x6 & ~x7 ;
  assign n135 = x8 & x12 ;
  assign n136 = n134 & n135 ;
  assign n137 = ~x5 & n136 ;
  assign n138 = n137 ^ n133 ;
  assign n140 = n139 ^ n138 ;
  assign n141 = n140 ^ n139 ;
  assign n142 = n141 ^ n133 ;
  assign n143 = ~x4 & x14 ;
  assign n144 = n143 ^ n140 ;
  assign n145 = n144 ^ n140 ;
  assign n146 = n145 ^ n142 ;
  assign n147 = n142 & n146 ;
  assign n149 = n148 ^ n147 ;
  assign n150 = n149 ^ n142 ;
  assign n151 = n133 ^ x3 ;
  assign n152 = n147 ^ n142 ;
  assign n153 = ~n151 & n152 ;
  assign n154 = n153 ^ n133 ;
  assign n155 = ~n150 & n154 ;
  assign n156 = n155 ^ n133 ;
  assign n157 = n156 ^ x9 ;
  assign n158 = n157 ^ n133 ;
  assign n159 = x13 & ~n158 ;
  assign n160 = n78 & n129 ;
  assign n161 = ~n130 & ~n160 ;
  assign n162 = ~n72 & ~n161 ;
  assign n163 = ~x9 & x12 ;
  assign n164 = x14 & n163 ;
  assign n165 = ~x8 & ~x13 ;
  assign n166 = n20 & n165 ;
  assign n167 = n164 & n166 ;
  assign n168 = ~n162 & ~n167 ;
  assign n169 = ~n159 & n168 ;
  assign n172 = n169 ^ x4 ;
  assign n173 = n172 ^ n169 ;
  assign n170 = n169 ^ n101 ;
  assign n171 = n170 ^ n169 ;
  assign n174 = n173 ^ n171 ;
  assign n175 = ~x9 & ~x13 ;
  assign n176 = n175 ^ n169 ;
  assign n177 = n176 ^ n169 ;
  assign n178 = n177 ^ n173 ;
  assign n179 = ~n173 & ~n178 ;
  assign n180 = n179 ^ n173 ;
  assign n181 = ~n174 & ~n180 ;
  assign n182 = n181 ^ n179 ;
  assign n183 = n182 ^ n169 ;
  assign n184 = n183 ^ n173 ;
  assign n185 = x11 & n184 ;
  assign n186 = n185 ^ n169 ;
  assign n187 = ~n127 & n186 ;
  assign n188 = n187 ^ x10 ;
  assign n189 = n188 ^ n187 ;
  assign n190 = ~x3 & ~x4 ;
  assign n191 = ~x11 & ~n190 ;
  assign n192 = ~x12 & n175 ;
  assign n193 = ~n191 & n192 ;
  assign n194 = ~x8 & x12 ;
  assign n195 = x7 & n194 ;
  assign n196 = ~n137 & ~n195 ;
  assign n197 = ~x3 & ~n196 ;
  assign n198 = x12 ^ x11 ;
  assign n199 = x14 ^ x12 ;
  assign n200 = n199 ^ x14 ;
  assign n201 = x0 & x14 ;
  assign n202 = ~x5 & x6 ;
  assign n203 = ~n201 & n202 ;
  assign n204 = ~n47 & n203 ;
  assign n205 = ~x4 & n204 ;
  assign n206 = n205 ^ x14 ;
  assign n207 = ~n200 & n206 ;
  assign n208 = n207 ^ x14 ;
  assign n209 = ~n198 & ~n208 ;
  assign n210 = n209 ^ x11 ;
  assign n211 = ~n197 & n210 ;
  assign n212 = n71 & ~n211 ;
  assign n213 = x3 & ~x11 ;
  assign n214 = n164 & n213 ;
  assign n215 = n109 & ~n163 ;
  assign n216 = n215 ^ x9 ;
  assign n217 = n216 ^ n215 ;
  assign n218 = n215 ^ x3 ;
  assign n219 = ~n217 & ~n218 ;
  assign n220 = n219 ^ n215 ;
  assign n221 = ~n48 & ~n215 ;
  assign n222 = n221 ^ n214 ;
  assign n223 = ~n220 & ~n222 ;
  assign n224 = n223 ^ n221 ;
  assign n225 = ~n214 & n224 ;
  assign n226 = n225 ^ n214 ;
  assign n227 = n226 ^ n214 ;
  assign n228 = ~n212 & n227 ;
  assign n229 = ~n193 & n228 ;
  assign n230 = n229 ^ n187 ;
  assign n231 = ~n189 & n230 ;
  assign n232 = n231 ^ n187 ;
  assign n233 = ~n46 & n232 ;
  assign y0 = ~n233 ;
endmodule
