module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 ;
  assign n21 = ~x4 & ~x5 ;
  assign n22 = x0 & ~n21 ;
  assign n24 = n22 ^ x7 ;
  assign n23 = n22 ^ x5 ;
  assign n25 = n24 ^ n23 ;
  assign n31 = n25 ^ n24 ;
  assign n27 = ~x1 & ~x4 ;
  assign n26 = n25 ^ x2 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = n28 ^ n22 ;
  assign n30 = n29 ^ n24 ;
  assign n32 = n31 ^ n30 ;
  assign n35 = n29 ^ n22 ;
  assign n33 = n27 ^ n22 ;
  assign n34 = n33 ^ n30 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = ~n32 & ~n36 ;
  assign n38 = n37 ^ n29 ;
  assign n39 = n38 ^ n33 ;
  assign n40 = n39 ^ n35 ;
  assign n41 = n34 ^ n31 ;
  assign n42 = ~n38 & ~n41 ;
  assign n43 = n42 ^ n29 ;
  assign n44 = n43 ^ n30 ;
  assign n45 = n44 ^ n31 ;
  assign n46 = n40 & n45 ;
  assign n9 = x4 ^ x1 ;
  assign n10 = x4 ^ x0 ;
  assign n11 = n10 ^ x4 ;
  assign n12 = n9 & n11 ;
  assign n13 = n12 ^ x4 ;
  assign n14 = x2 & x4 ;
  assign n15 = n14 ^ x5 ;
  assign n16 = n13 & n15 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = x5 & n17 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = n19 ^ x5 ;
  assign n47 = n46 ^ n20 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = n46 ^ x7 ;
  assign n50 = n49 ^ n46 ;
  assign n51 = ~n48 & n50 ;
  assign n52 = n51 ^ n46 ;
  assign n53 = ~x6 & n52 ;
  assign n54 = n53 ^ n46 ;
  assign y0 = n54 ;
endmodule
