module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 ;
  assign n16 = x13 & ~x14 ;
  assign n17 = ~x10 & ~x12 ;
  assign n18 = n16 & n17 ;
  assign n19 = x7 & x10 ;
  assign n20 = ~x8 & n19 ;
  assign n21 = x1 & x4 ;
  assign n22 = ~x5 & x12 ;
  assign n23 = ~x0 & x3 ;
  assign n24 = n22 & n23 ;
  assign n25 = n16 & n24 ;
  assign n26 = n21 & n25 ;
  assign n27 = n20 & n26 ;
  assign n28 = ~x0 & ~x3 ;
  assign n29 = n28 ^ x10 ;
  assign n30 = n29 ^ x10 ;
  assign n31 = x10 ^ x4 ;
  assign n32 = n31 ^ x10 ;
  assign n33 = n30 & n32 ;
  assign n34 = n33 ^ x10 ;
  assign n35 = x5 & ~n34 ;
  assign n36 = n35 ^ x10 ;
  assign n37 = x14 & ~n36 ;
  assign n38 = n37 ^ x10 ;
  assign n39 = n38 ^ x12 ;
  assign n52 = n39 ^ n38 ;
  assign n40 = x7 & ~x12 ;
  assign n41 = x8 & ~x14 ;
  assign n42 = ~x4 & ~x5 ;
  assign n43 = ~x6 & n42 ;
  assign n44 = n41 & n43 ;
  assign n45 = n40 & n44 ;
  assign n46 = n45 ^ n39 ;
  assign n47 = n46 ^ n38 ;
  assign n48 = n39 ^ n37 ;
  assign n49 = n48 ^ n45 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = n47 & ~n50 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n53 ^ n47 ;
  assign n55 = ~x4 & x14 ;
  assign n56 = ~x0 & ~x2 ;
  assign n57 = x4 & x5 ;
  assign n58 = x3 & x8 ;
  assign n59 = ~x1 & ~x6 ;
  assign n60 = ~n58 & ~n59 ;
  assign n61 = n57 & n60 ;
  assign n62 = n56 & n61 ;
  assign n63 = ~n55 & ~n62 ;
  assign n64 = n63 ^ n38 ;
  assign n65 = n51 ^ n47 ;
  assign n66 = n64 & n65 ;
  assign n67 = n66 ^ n38 ;
  assign n68 = ~n54 & n67 ;
  assign n69 = n68 ^ n38 ;
  assign n70 = n69 ^ x10 ;
  assign n71 = n70 ^ n38 ;
  assign n72 = ~x13 & n71 ;
  assign n73 = ~x3 & n17 ;
  assign n74 = ~n72 & ~n73 ;
  assign n75 = ~n27 & n74 ;
  assign n76 = n75 ^ x9 ;
  assign n77 = n76 ^ n75 ;
  assign n78 = x3 & ~x8 ;
  assign n79 = ~x7 & ~n78 ;
  assign n80 = n42 & n79 ;
  assign n81 = ~x3 & x8 ;
  assign n82 = ~x6 & ~n81 ;
  assign n83 = ~x0 & ~x13 ;
  assign n84 = x10 & n83 ;
  assign n85 = ~x12 & n84 ;
  assign n86 = ~n82 & n85 ;
  assign n87 = n80 & n86 ;
  assign n88 = ~x1 & ~x12 ;
  assign n89 = ~x13 & x14 ;
  assign n90 = ~n88 & n89 ;
  assign n91 = ~n83 & ~n90 ;
  assign n92 = ~x10 & n91 ;
  assign n93 = ~n87 & ~n92 ;
  assign n94 = n93 ^ n75 ;
  assign n95 = n77 & n94 ;
  assign n96 = n95 ^ n75 ;
  assign n97 = ~n18 & n96 ;
  assign n98 = x11 & ~n97 ;
  assign n99 = x9 & x12 ;
  assign n100 = n99 ^ x6 ;
  assign n101 = x11 & x14 ;
  assign n102 = n101 ^ n100 ;
  assign n103 = n102 ^ n99 ;
  assign n104 = n103 ^ n102 ;
  assign n105 = ~x11 & n42 ;
  assign n106 = n28 & n40 ;
  assign n107 = ~x7 & x8 ;
  assign n108 = x9 & n107 ;
  assign n109 = n108 ^ x14 ;
  assign n110 = n109 ^ n106 ;
  assign n111 = ~x3 & x7 ;
  assign n112 = n111 ^ x0 ;
  assign n113 = x14 & n112 ;
  assign n114 = n113 ^ n111 ;
  assign n115 = n110 & ~n114 ;
  assign n116 = n115 ^ n113 ;
  assign n117 = n116 ^ n111 ;
  assign n118 = n117 ^ x14 ;
  assign n119 = ~n106 & ~n118 ;
  assign n120 = n105 & ~n119 ;
  assign n121 = n120 ^ n102 ;
  assign n122 = n121 ^ n100 ;
  assign n123 = n104 & n122 ;
  assign n124 = n123 ^ n120 ;
  assign n125 = ~x8 & n111 ;
  assign n126 = ~n120 & ~n125 ;
  assign n127 = n126 ^ n100 ;
  assign n128 = ~n124 & ~n127 ;
  assign n129 = n128 ^ n126 ;
  assign n130 = ~n100 & n129 ;
  assign n131 = n130 ^ n123 ;
  assign n132 = n131 ^ x6 ;
  assign n133 = n132 ^ n120 ;
  assign n134 = ~x10 & ~n133 ;
  assign n135 = x5 & x10 ;
  assign n136 = x14 & n135 ;
  assign n137 = n60 & n136 ;
  assign n138 = x5 & ~x7 ;
  assign n139 = ~x11 & ~x14 ;
  assign n140 = ~x3 & n139 ;
  assign n141 = ~n138 & n140 ;
  assign n142 = ~n137 & ~n141 ;
  assign n143 = ~x0 & ~n142 ;
  assign n144 = x5 & x6 ;
  assign n145 = n139 & n144 ;
  assign n146 = n111 & n145 ;
  assign n147 = ~n143 & ~n146 ;
  assign n148 = ~x12 & ~n147 ;
  assign n149 = n148 ^ x4 ;
  assign n150 = n149 ^ n148 ;
  assign n151 = ~x6 & n20 ;
  assign n152 = ~x3 & n22 ;
  assign n153 = n151 & n152 ;
  assign n154 = x14 & n153 ;
  assign n155 = ~n73 & ~n154 ;
  assign n156 = n155 ^ n148 ;
  assign n157 = ~n150 & ~n156 ;
  assign n158 = n157 ^ n148 ;
  assign n159 = ~x9 & n158 ;
  assign n160 = ~n134 & ~n159 ;
  assign n161 = ~x13 & ~n160 ;
  assign n162 = ~x14 & ~n17 ;
  assign n163 = ~x3 & ~n162 ;
  assign n164 = n43 & n107 ;
  assign n165 = n164 ^ x9 ;
  assign n166 = x12 & ~n165 ;
  assign n167 = n166 ^ x9 ;
  assign n168 = n163 & ~n167 ;
  assign n169 = n168 ^ x14 ;
  assign n170 = x0 & ~n144 ;
  assign n171 = x4 & ~n138 ;
  assign n172 = ~n170 & n171 ;
  assign n173 = ~x12 & ~n172 ;
  assign n174 = ~x11 & x13 ;
  assign n175 = ~n173 & n174 ;
  assign n176 = x10 & n175 ;
  assign n177 = n176 ^ n168 ;
  assign n178 = n177 ^ n176 ;
  assign n179 = n178 ^ n169 ;
  assign n180 = ~x9 & x12 ;
  assign n181 = ~x10 & n180 ;
  assign n182 = n181 ^ x11 ;
  assign n183 = ~x11 & ~n182 ;
  assign n184 = n183 ^ n176 ;
  assign n185 = n184 ^ x11 ;
  assign n186 = n179 & n185 ;
  assign n187 = n186 ^ n183 ;
  assign n188 = n187 ^ x11 ;
  assign n189 = ~n169 & ~n188 ;
  assign n190 = n189 ^ n168 ;
  assign n191 = ~n161 & ~n190 ;
  assign n192 = ~n98 & n191 ;
  assign y0 = ~n192 ;
endmodule
