module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 ;
  output y0 ;
  wire n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 ;
  assign n26 = x1 ^ x0 ;
  assign n27 = x2 ^ x1 ;
  assign n28 = n27 ^ x5 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = x5 ^ x3 ;
  assign n31 = x5 ^ x1 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = ~n30 & ~n32 ;
  assign n34 = n33 ^ x5 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n29 & ~n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ n30 ;
  assign n39 = n26 & ~n38 ;
  assign n40 = ~x4 & n39 ;
  assign n41 = x14 & ~n40 ;
  assign n236 = ~x19 & ~x20 ;
  assign n42 = ~x12 & ~x13 ;
  assign n43 = x9 ^ x1 ;
  assign n44 = ~x6 & ~x7 ;
  assign n45 = x8 & x11 ;
  assign n46 = n44 & n45 ;
  assign n47 = ~x10 & n46 ;
  assign n48 = x3 & ~x4 ;
  assign n49 = ~x0 & ~x2 ;
  assign n50 = n48 & n49 ;
  assign n51 = n47 & n50 ;
  assign n52 = n51 ^ n43 ;
  assign n53 = n52 ^ x9 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = ~x8 & n44 ;
  assign n56 = ~x11 & n55 ;
  assign n57 = x10 & n56 ;
  assign n58 = x0 & x2 ;
  assign n59 = ~x3 & n58 ;
  assign n60 = n57 & n59 ;
  assign n61 = n60 ^ n52 ;
  assign n62 = n61 ^ n43 ;
  assign n63 = n54 & ~n62 ;
  assign n64 = n63 ^ n60 ;
  assign n65 = ~x2 & x3 ;
  assign n66 = ~x10 & n65 ;
  assign n67 = ~x4 & n66 ;
  assign n68 = ~n59 & ~n67 ;
  assign n69 = n56 & ~n68 ;
  assign n70 = n48 ^ x3 ;
  assign n71 = ~n58 & ~n70 ;
  assign n72 = n71 ^ x3 ;
  assign n73 = n47 & ~n72 ;
  assign n74 = x8 & x10 ;
  assign n75 = ~x11 & n74 ;
  assign n76 = ~n50 & ~n59 ;
  assign n77 = n75 & ~n76 ;
  assign n78 = ~n73 & ~n77 ;
  assign n79 = ~n69 & n78 ;
  assign n80 = ~n60 & n79 ;
  assign n81 = n80 ^ n43 ;
  assign n82 = ~n64 & n81 ;
  assign n83 = n82 ^ n80 ;
  assign n84 = n43 & n83 ;
  assign n85 = n84 ^ n63 ;
  assign n86 = n85 ^ x1 ;
  assign n87 = n86 ^ n60 ;
  assign n88 = n42 & n87 ;
  assign n89 = x1 & x2 ;
  assign n90 = ~x6 & ~x13 ;
  assign n91 = ~x9 & x11 ;
  assign n92 = n74 & n91 ;
  assign n93 = ~x12 & ~n92 ;
  assign n94 = ~x7 & x16 ;
  assign n95 = x4 & n94 ;
  assign n96 = ~x0 & n95 ;
  assign n97 = ~n93 & n96 ;
  assign n98 = n90 & n97 ;
  assign n99 = n89 & n98 ;
  assign n100 = x0 & ~x21 ;
  assign n101 = ~x1 & ~n100 ;
  assign n102 = x9 & n42 ;
  assign n103 = ~x4 & n102 ;
  assign n104 = ~n101 & ~n103 ;
  assign n105 = n65 & ~n104 ;
  assign n106 = x5 & ~n105 ;
  assign n107 = ~n99 & n106 ;
  assign n108 = ~x4 & ~x22 ;
  assign n109 = ~x0 & ~n108 ;
  assign n110 = ~n49 & ~n109 ;
  assign n111 = ~x1 & n110 ;
  assign n112 = x6 & ~n45 ;
  assign n113 = x15 ^ x12 ;
  assign n114 = x13 & n113 ;
  assign n115 = n114 ^ x12 ;
  assign n116 = ~n112 & ~n115 ;
  assign n117 = n91 & ~n94 ;
  assign n118 = n116 & ~n117 ;
  assign n119 = ~x6 & x9 ;
  assign n120 = x7 & x10 ;
  assign n121 = ~n119 & ~n120 ;
  assign n122 = x10 ^ x8 ;
  assign n123 = n122 ^ x10 ;
  assign n124 = x13 ^ x10 ;
  assign n125 = n123 & n124 ;
  assign n126 = n125 ^ x10 ;
  assign n127 = ~x17 & ~n126 ;
  assign n128 = n121 & n127 ;
  assign n129 = ~x10 & n42 ;
  assign n130 = n129 ^ x12 ;
  assign n131 = n130 ^ x8 ;
  assign n132 = n131 ^ n130 ;
  assign n133 = n130 ^ x7 ;
  assign n134 = n133 ^ n130 ;
  assign n135 = n132 & ~n134 ;
  assign n136 = n135 ^ n130 ;
  assign n137 = x11 & n136 ;
  assign n138 = n137 ^ n130 ;
  assign n139 = n128 & ~n138 ;
  assign n140 = n118 & n139 ;
  assign n141 = n140 ^ x2 ;
  assign n142 = n141 ^ n140 ;
  assign n143 = ~x0 & x15 ;
  assign n144 = n143 ^ n140 ;
  assign n145 = ~n142 & n144 ;
  assign n146 = n145 ^ n140 ;
  assign n147 = n27 & ~n146 ;
  assign n148 = n147 ^ x1 ;
  assign n149 = x4 & n148 ;
  assign n150 = x2 & x23 ;
  assign n151 = n150 ^ x4 ;
  assign n152 = n151 ^ n150 ;
  assign n153 = n152 ^ x0 ;
  assign n154 = x10 & x11 ;
  assign n155 = x9 & n154 ;
  assign n156 = ~x12 & n155 ;
  assign n157 = n156 ^ x13 ;
  assign n158 = ~n156 & n157 ;
  assign n159 = n158 ^ n150 ;
  assign n160 = n159 ^ n156 ;
  assign n161 = n153 & ~n160 ;
  assign n162 = n161 ^ n158 ;
  assign n163 = n162 ^ n156 ;
  assign n164 = x0 & ~n163 ;
  assign n165 = n164 ^ x0 ;
  assign n166 = ~n149 & ~n165 ;
  assign n167 = ~n111 & n166 ;
  assign n168 = n167 ^ x3 ;
  assign n169 = n168 ^ n167 ;
  assign n170 = n169 ^ n107 ;
  assign n171 = ~x12 & n44 ;
  assign n172 = ~x13 & ~n171 ;
  assign n173 = ~x8 & ~x10 ;
  assign n174 = n91 & n173 ;
  assign n175 = ~n172 & n174 ;
  assign n176 = ~n55 & ~n74 ;
  assign n177 = ~x8 & x10 ;
  assign n178 = ~x9 & ~n177 ;
  assign n179 = ~x11 & n42 ;
  assign n180 = ~n178 & n179 ;
  assign n181 = ~n176 & n180 ;
  assign n182 = ~n175 & ~n181 ;
  assign n183 = ~n89 & n182 ;
  assign n184 = n183 ^ x4 ;
  assign n185 = ~x4 & n184 ;
  assign n186 = n185 ^ n167 ;
  assign n187 = n186 ^ x4 ;
  assign n188 = n170 & n187 ;
  assign n189 = n188 ^ n185 ;
  assign n190 = n189 ^ x4 ;
  assign n191 = n107 & ~n190 ;
  assign n192 = n191 ^ n107 ;
  assign n193 = x4 ^ x3 ;
  assign n194 = x0 & ~x1 ;
  assign n195 = n56 & n65 ;
  assign n196 = n102 & n195 ;
  assign n197 = ~x4 & ~n196 ;
  assign n198 = n194 & ~n197 ;
  assign n199 = ~x5 & ~n198 ;
  assign n200 = n199 ^ n193 ;
  assign n201 = x1 & n49 ;
  assign n202 = ~n58 & ~n201 ;
  assign n203 = n202 ^ x3 ;
  assign n204 = n203 ^ n202 ;
  assign n205 = ~x15 & x23 ;
  assign n206 = x24 & ~n205 ;
  assign n207 = n49 & ~n206 ;
  assign n208 = n42 & n89 ;
  assign n209 = n56 ^ x9 ;
  assign n210 = n56 ^ x10 ;
  assign n211 = n210 ^ x10 ;
  assign n212 = n75 ^ x10 ;
  assign n213 = ~n211 & ~n212 ;
  assign n214 = n213 ^ x10 ;
  assign n215 = n209 ^ n47 ;
  assign n216 = ~n214 & n215 ;
  assign n217 = n216 ^ n47 ;
  assign n218 = n209 & n217 ;
  assign n219 = n218 ^ x9 ;
  assign n220 = n219 ^ n209 ;
  assign n221 = n208 & n220 ;
  assign n222 = ~n207 & ~n221 ;
  assign n223 = n222 ^ n202 ;
  assign n224 = ~n204 & n223 ;
  assign n225 = n224 ^ n202 ;
  assign n226 = n225 ^ n193 ;
  assign n227 = ~n200 & n226 ;
  assign n228 = n227 ^ n224 ;
  assign n229 = n228 ^ n202 ;
  assign n230 = n229 ^ n199 ;
  assign n231 = ~n193 & ~n230 ;
  assign n232 = n231 ^ n193 ;
  assign n233 = n232 ^ n199 ;
  assign n234 = ~n192 & n233 ;
  assign n235 = ~n88 & ~n234 ;
  assign n237 = n236 ^ n235 ;
  assign n238 = n237 ^ n235 ;
  assign n239 = n235 ^ x18 ;
  assign n240 = ~n238 & n239 ;
  assign n241 = n240 ^ n235 ;
  assign n242 = n41 & n241 ;
  assign y0 = ~n242 ;
endmodule
