module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 ;
  assign n17 = ~x0 & ~x1 ;
  assign n18 = x2 & ~x15 ;
  assign n19 = n17 & n18 ;
  assign n20 = ~x8 & x9 ;
  assign n21 = ~x3 & x11 ;
  assign n22 = x14 & n21 ;
  assign n23 = x4 & x5 ;
  assign n24 = ~x6 & x10 ;
  assign n25 = n23 & n24 ;
  assign n26 = n22 & n25 ;
  assign n27 = n20 & n26 ;
  assign n28 = n19 & n27 ;
  assign n29 = ~x4 & ~x10 ;
  assign n30 = ~x9 & n29 ;
  assign n31 = ~x6 & ~x7 ;
  assign n32 = ~x1 & n31 ;
  assign n33 = n30 & n32 ;
  assign n34 = ~x2 & ~x5 ;
  assign n35 = ~x0 & ~x8 ;
  assign n36 = ~x3 & n35 ;
  assign n37 = n34 & n36 ;
  assign n38 = n33 & n37 ;
  assign n39 = ~x5 & x6 ;
  assign n40 = x7 & n39 ;
  assign n41 = x0 & x1 ;
  assign n42 = x3 & x4 ;
  assign n43 = ~x2 & n42 ;
  assign n44 = n41 & n43 ;
  assign n45 = n40 & n44 ;
  assign n46 = ~n38 & ~n45 ;
  assign n47 = x15 & ~n46 ;
  assign n48 = x5 & n19 ;
  assign n49 = x4 & x9 ;
  assign n50 = n24 & n49 ;
  assign n51 = n50 ^ n30 ;
  assign n52 = n51 ^ n50 ;
  assign n53 = x6 & x7 ;
  assign n54 = n53 ^ n50 ;
  assign n55 = n54 ^ n50 ;
  assign n56 = n52 & n55 ;
  assign n57 = n56 ^ n50 ;
  assign n58 = x3 & n57 ;
  assign n59 = n58 ^ n50 ;
  assign n60 = n48 & n59 ;
  assign n61 = ~x8 & n60 ;
  assign n62 = ~n47 & ~n61 ;
  assign n63 = n62 ^ x14 ;
  assign n64 = n63 ^ n62 ;
  assign n65 = n64 ^ x13 ;
  assign n66 = x1 & x15 ;
  assign n67 = n35 & n66 ;
  assign n68 = x2 & x9 ;
  assign n69 = x5 & n68 ;
  assign n70 = n31 & n69 ;
  assign n71 = n67 & n70 ;
  assign n72 = ~x1 & x10 ;
  assign n73 = n40 & n72 ;
  assign n74 = ~x2 & ~x8 ;
  assign n75 = x15 & n74 ;
  assign n76 = ~x9 & n75 ;
  assign n77 = n76 ^ x0 ;
  assign n78 = n77 ^ n76 ;
  assign n79 = x9 ^ x8 ;
  assign n80 = n18 & ~n79 ;
  assign n81 = n80 ^ n76 ;
  assign n82 = n78 & n81 ;
  assign n83 = n82 ^ n76 ;
  assign n84 = n73 & n83 ;
  assign n85 = ~n71 & ~n84 ;
  assign n86 = n42 & ~n85 ;
  assign n87 = ~x4 & ~x15 ;
  assign n90 = x0 & ~x9 ;
  assign n91 = x7 & n90 ;
  assign n88 = ~x7 & x9 ;
  assign n89 = n41 & n88 ;
  assign n92 = n91 ^ n89 ;
  assign n93 = n92 ^ x8 ;
  assign n100 = n93 ^ n92 ;
  assign n94 = n93 ^ x1 ;
  assign n95 = n94 ^ n92 ;
  assign n96 = n93 ^ n89 ;
  assign n97 = n96 ^ x1 ;
  assign n98 = n97 ^ n95 ;
  assign n99 = ~n95 & ~n98 ;
  assign n101 = n100 ^ n99 ;
  assign n102 = n101 ^ n95 ;
  assign n103 = n92 ^ x2 ;
  assign n104 = n99 ^ n95 ;
  assign n105 = n103 & ~n104 ;
  assign n106 = n105 ^ n92 ;
  assign n107 = ~n102 & n106 ;
  assign n108 = n107 ^ n92 ;
  assign n109 = n108 ^ n91 ;
  assign n110 = n109 ^ n92 ;
  assign n111 = n39 & n110 ;
  assign n112 = x5 & n17 ;
  assign n113 = ~x6 & n112 ;
  assign n114 = n113 ^ x2 ;
  assign n122 = n114 ^ n113 ;
  assign n115 = n114 ^ x5 ;
  assign n116 = n115 ^ n113 ;
  assign n117 = x6 & n41 ;
  assign n118 = n117 ^ x5 ;
  assign n119 = n118 ^ x5 ;
  assign n120 = n119 ^ n116 ;
  assign n121 = ~n116 & ~n120 ;
  assign n123 = n122 ^ n121 ;
  assign n124 = n123 ^ n116 ;
  assign n125 = n113 ^ x9 ;
  assign n126 = n121 ^ n116 ;
  assign n127 = ~n125 & ~n126 ;
  assign n128 = n127 ^ n113 ;
  assign n129 = n124 & ~n128 ;
  assign n130 = n129 ^ n113 ;
  assign n131 = n130 ^ x2 ;
  assign n132 = n131 ^ n113 ;
  assign n133 = x8 & ~n132 ;
  assign n134 = x7 & n133 ;
  assign n135 = ~n111 & ~n134 ;
  assign n136 = n87 & ~n135 ;
  assign n137 = n136 ^ x3 ;
  assign n138 = n137 ^ n136 ;
  assign n139 = n23 & n88 ;
  assign n140 = n139 ^ n40 ;
  assign n141 = n140 ^ n139 ;
  assign n142 = n139 ^ n49 ;
  assign n143 = n142 ^ n139 ;
  assign n144 = n141 & n143 ;
  assign n145 = n144 ^ n139 ;
  assign n146 = ~x2 & n145 ;
  assign n147 = n146 ^ n139 ;
  assign n148 = n67 & n147 ;
  assign n149 = x1 & ~x2 ;
  assign n150 = n39 & ~n149 ;
  assign n151 = ~n74 & n90 ;
  assign n152 = n150 & n151 ;
  assign n153 = n152 ^ x9 ;
  assign n154 = n153 ^ n152 ;
  assign n155 = x0 & x8 ;
  assign n156 = n150 & n155 ;
  assign n157 = n74 & n113 ;
  assign n158 = ~n156 & ~n157 ;
  assign n159 = n158 ^ n152 ;
  assign n160 = n159 ^ n152 ;
  assign n161 = n154 & ~n160 ;
  assign n162 = n161 ^ n152 ;
  assign n163 = ~x7 & n162 ;
  assign n164 = n163 ^ n152 ;
  assign n165 = n87 & n164 ;
  assign n166 = ~n148 & ~n165 ;
  assign n167 = n166 ^ n136 ;
  assign n168 = n138 & ~n167 ;
  assign n169 = n168 ^ n136 ;
  assign n170 = ~x10 & n169 ;
  assign n171 = n170 ^ n86 ;
  assign n172 = ~n86 & n171 ;
  assign n173 = n172 ^ n62 ;
  assign n174 = n173 ^ n86 ;
  assign n175 = n65 & ~n174 ;
  assign n176 = n175 ^ n172 ;
  assign n177 = n176 ^ n86 ;
  assign n178 = ~x13 & ~n177 ;
  assign n179 = n178 ^ x13 ;
  assign n180 = ~n28 & n179 ;
  assign n181 = ~x12 & ~n180 ;
  assign y0 = n181 ;
endmodule
