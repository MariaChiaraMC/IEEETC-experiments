module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 ;
  assign n13 = ~x6 & ~x11 ;
  assign n14 = x5 & x10 ;
  assign n15 = x4 & n14 ;
  assign n16 = x7 & ~n15 ;
  assign n17 = ~n13 & ~n16 ;
  assign n18 = x5 & x9 ;
  assign n19 = x4 & x6 ;
  assign n20 = ~n18 & n19 ;
  assign n21 = ~x8 & ~n20 ;
  assign n22 = x0 & ~n21 ;
  assign n23 = ~n17 & n22 ;
  assign n24 = n23 ^ x1 ;
  assign n25 = x3 & x4 ;
  assign n26 = ~x7 & n25 ;
  assign n27 = n26 ^ n18 ;
  assign n28 = n27 ^ n18 ;
  assign n29 = x9 ^ x8 ;
  assign n30 = x11 & n19 ;
  assign n31 = n30 ^ x9 ;
  assign n32 = x8 ^ x5 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n30 & ~n33 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n31 & n35 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = n37 ^ n30 ;
  assign n39 = n38 ^ n32 ;
  assign n40 = ~n29 & ~n39 ;
  assign n41 = n40 ^ x8 ;
  assign n42 = x2 & ~n41 ;
  assign n43 = x6 ^ x4 ;
  assign n44 = n43 ^ x6 ;
  assign n45 = x6 ^ x3 ;
  assign n46 = n44 & n45 ;
  assign n47 = n46 ^ x6 ;
  assign n48 = x7 & ~n47 ;
  assign n49 = n42 & ~n48 ;
  assign n50 = n49 ^ n18 ;
  assign n51 = ~n28 & n50 ;
  assign n52 = n51 ^ n18 ;
  assign n53 = n52 ^ n23 ;
  assign n54 = ~n24 & n53 ;
  assign n55 = n54 ^ n51 ;
  assign n56 = n55 ^ n18 ;
  assign n57 = n56 ^ x1 ;
  assign n58 = n23 & ~n57 ;
  assign n59 = n58 ^ n23 ;
  assign y0 = n59 ;
endmodule
