module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 ;
  assign n7 = x5 ^ x4 ;
  assign n8 = x3 ^ x2 ;
  assign n9 = x1 ^ x0 ;
  assign n10 = n9 ^ n8 ;
  assign n11 = x4 ^ x1 ;
  assign n12 = x3 ^ x1 ;
  assign n13 = n11 & ~n12 ;
  assign n14 = n13 ^ x1 ;
  assign n15 = n14 ^ n8 ;
  assign n16 = ~n10 & ~n15 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n17 ^ x1 ;
  assign n19 = n18 ^ n9 ;
  assign n20 = ~n8 & n19 ;
  assign n21 = n20 ^ n8 ;
  assign n22 = n7 & ~n21 ;
  assign y0 = n22 ;
endmodule
