module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 ;
  assign n9 = ~x0 & ~x2 ;
  assign n10 = ~x1 & n9 ;
  assign n13 = x4 ^ x3 ;
  assign n19 = x7 ^ x5 ;
  assign n11 = x5 ^ x3 ;
  assign n20 = n19 ^ n11 ;
  assign n21 = n20 ^ x5 ;
  assign n12 = n11 ^ x6 ;
  assign n14 = n13 ^ n12 ;
  assign n22 = n21 ^ n14 ;
  assign n23 = n22 ^ n13 ;
  assign n24 = ~n13 & n23 ;
  assign n25 = n24 ^ n11 ;
  assign n26 = n25 ^ n14 ;
  assign n27 = n26 ^ n13 ;
  assign n28 = n27 ^ x5 ;
  assign n29 = n14 ^ n13 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = ~n26 & ~n30 ;
  assign n32 = n31 ^ n11 ;
  assign n33 = n32 ^ n14 ;
  assign n34 = n33 ^ n13 ;
  assign n35 = n34 ^ x5 ;
  assign n36 = ~n28 & ~n35 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = n16 & ~n17 ;
  assign n37 = n36 ^ n18 ;
  assign n38 = n37 ^ n24 ;
  assign n39 = n38 ^ n11 ;
  assign n40 = n39 ^ n14 ;
  assign n41 = n40 ^ n13 ;
  assign n42 = n41 ^ x5 ;
  assign n43 = n42 ^ x3 ;
  assign n44 = n10 & ~n43 ;
  assign y0 = n44 ;
endmodule
