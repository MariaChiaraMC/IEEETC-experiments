module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 ;
  assign n8 = x6 ^ x1 ;
  assign n9 = ~x4 & ~x5 ;
  assign n10 = ~x3 & n9 ;
  assign n11 = ~x2 & n10 ;
  assign n12 = n11 ^ x6 ;
  assign n13 = n11 ^ x0 ;
  assign n14 = n11 & ~n13 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = ~n12 & n15 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = n17 ^ n11 ;
  assign n19 = n18 ^ x0 ;
  assign n20 = n8 & ~n19 ;
  assign n21 = n20 ^ x0 ;
  assign y0 = ~n21 ;
endmodule
