module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n7 = x4 ^ x2 ;
  assign n8 = n7 ^ x0 ;
  assign n9 = n8 ^ x4 ;
  assign n10 = n9 ^ n7 ;
  assign n11 = n9 ^ x4 ;
  assign n12 = ~n10 & n11 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = n13 ^ x3 ;
  assign n15 = n7 ^ x1 ;
  assign n16 = n15 ^ x4 ;
  assign n17 = ~x5 & ~n16 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = n19 ^ n15 ;
  assign n21 = n20 ^ n10 ;
  assign n22 = n21 ^ x3 ;
  assign n23 = n16 ^ x3 ;
  assign n24 = n15 ^ n11 ;
  assign n25 = n24 ^ n10 ;
  assign n26 = n25 ^ x3 ;
  assign n27 = ~n23 & n26 ;
  assign n28 = n27 ^ x4 ;
  assign n29 = n28 ^ n15 ;
  assign n30 = ~n22 & ~n29 ;
  assign n31 = n30 ^ x3 ;
  assign n32 = n14 & n31 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ x3 ;
  assign y0 = n34 ;
endmodule
