module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 ;
  assign n9 = x3 ^ x2 ;
  assign n10 = x1 & n9 ;
  assign n11 = ~x0 & ~n10 ;
  assign n14 = x5 ^ x2 ;
  assign n15 = n14 ^ x7 ;
  assign n12 = x7 ^ x6 ;
  assign n13 = n12 ^ x2 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n17 ^ n12 ;
  assign n19 = x5 ^ x4 ;
  assign n20 = n19 ^ x7 ;
  assign n21 = n20 ^ n12 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n23 ^ n15 ;
  assign n25 = n24 ^ n12 ;
  assign n26 = n25 ^ n19 ;
  assign n32 = n26 ^ n19 ;
  assign n33 = n32 ^ n18 ;
  assign n34 = n33 ^ n23 ;
  assign n35 = ~n18 & n34 ;
  assign n27 = n26 ^ n18 ;
  assign n28 = n18 ^ n12 ;
  assign n29 = n28 ^ n18 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = ~n27 & ~n30 ;
  assign n36 = n35 ^ n31 ;
  assign n37 = n36 ^ n18 ;
  assign n38 = n37 ^ n26 ;
  assign n39 = n32 ^ n26 ;
  assign n40 = n31 ^ n28 ;
  assign n41 = n40 ^ n26 ;
  assign n42 = ~n39 & n41 ;
  assign n43 = n42 ^ n31 ;
  assign n44 = n43 ^ n18 ;
  assign n45 = n44 ^ n32 ;
  assign n46 = n45 ^ n23 ;
  assign n47 = ~n38 & n46 ;
  assign n48 = n47 ^ n42 ;
  assign n49 = ~x3 & ~n48 ;
  assign n50 = x2 & x3 ;
  assign n51 = x4 & ~x5 ;
  assign n52 = n50 & n51 ;
  assign n53 = ~x1 & ~n52 ;
  assign n54 = ~n49 & n53 ;
  assign n55 = n11 & ~n54 ;
  assign y0 = n55 ;
endmodule
