module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 ;
  assign n16 = ~x12 & ~x14 ;
  assign n17 = x10 ^ x8 ;
  assign n18 = x4 ^ x3 ;
  assign n19 = n18 ^ x10 ;
  assign n20 = ~x10 & n19 ;
  assign n21 = n20 ^ x10 ;
  assign n22 = n17 & ~n21 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n23 ^ x10 ;
  assign n25 = n24 ^ n18 ;
  assign n26 = ~x4 & n25 ;
  assign n27 = n26 ^ n18 ;
  assign n28 = n16 & ~n27 ;
  assign n29 = x6 ^ x5 ;
  assign n30 = x8 & x10 ;
  assign n31 = n30 ^ x5 ;
  assign n32 = n30 ^ x11 ;
  assign n33 = ~n30 & n32 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = ~n31 & ~n34 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = n37 ^ x11 ;
  assign n39 = n29 & n38 ;
  assign n40 = n28 & n39 ;
  assign n41 = x3 & ~x5 ;
  assign n42 = n41 ^ x2 ;
  assign n43 = x2 ^ x0 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = x1 & x13 ;
  assign n46 = x7 & n45 ;
  assign n47 = n46 ^ n41 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = ~x9 & ~x13 ;
  assign n50 = ~x1 & ~x7 ;
  assign n51 = n49 & n50 ;
  assign n52 = n51 ^ n46 ;
  assign n53 = ~n48 & n52 ;
  assign n54 = n53 ^ n46 ;
  assign n55 = n54 ^ n42 ;
  assign n56 = n44 & n55 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n57 ^ n46 ;
  assign n59 = n58 ^ n43 ;
  assign n60 = n42 & n59 ;
  assign n61 = n60 ^ n42 ;
  assign n62 = n40 & n61 ;
  assign y0 = n62 ;
endmodule
