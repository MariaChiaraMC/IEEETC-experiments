module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 ;
  assign n17 = x1 ^ x0 ;
  assign n18 = n17 ^ x0 ;
  assign n19 = ~x5 & x7 ;
  assign n20 = x4 & ~x7 ;
  assign n21 = x5 & ~n20 ;
  assign n22 = ~x6 & n21 ;
  assign n23 = x10 ^ x9 ;
  assign n24 = ~x12 & n23 ;
  assign n25 = ~n22 & n24 ;
  assign n26 = ~x8 & ~x11 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = x15 ^ x14 ;
  assign n29 = n28 ^ x13 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = ~x14 & ~x15 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = n30 & n32 ;
  assign n34 = n33 ^ n28 ;
  assign n35 = n34 ^ n25 ;
  assign n36 = n27 & n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ n28 ;
  assign n39 = n38 ^ n26 ;
  assign n40 = n25 & n39 ;
  assign n41 = n40 ^ n25 ;
  assign n42 = ~n19 & ~n41 ;
  assign n43 = ~x0 & ~x2 ;
  assign n44 = ~n42 & n43 ;
  assign n45 = n44 ^ x0 ;
  assign n46 = n18 & n45 ;
  assign n47 = n46 ^ x0 ;
  assign n48 = ~x3 & n47 ;
  assign y0 = n48 ;
endmodule
