module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ;
  assign n11 = ~x2 & ~x3 ;
  assign n12 = ~x5 & n11 ;
  assign n13 = ~x6 & x8 ;
  assign n14 = n12 & n13 ;
  assign n15 = x4 & ~n14 ;
  assign n16 = ~x0 & ~n15 ;
  assign n17 = ~x1 & n16 ;
  assign n18 = x6 & n12 ;
  assign n19 = ~x4 & ~n18 ;
  assign n20 = x3 ^ x2 ;
  assign n21 = x8 ^ x7 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = x9 ^ x3 ;
  assign n24 = ~x7 & ~n23 ;
  assign n25 = n24 ^ x9 ;
  assign n26 = n22 & n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n27 ^ x9 ;
  assign n29 = n28 ^ x7 ;
  assign n30 = n20 & ~n29 ;
  assign n31 = n30 ^ x2 ;
  assign n32 = ~x7 & ~x8 ;
  assign n33 = ~x2 & n32 ;
  assign n34 = ~x6 & ~n33 ;
  assign n35 = n11 ^ x5 ;
  assign n36 = n34 & ~n35 ;
  assign n37 = ~n31 & n36 ;
  assign n38 = n19 & ~n37 ;
  assign n39 = n17 & ~n38 ;
  assign y0 = n39 ;
endmodule
