module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 ;
  assign n16 = ~x3 & ~x6 ;
  assign n17 = x10 & n16 ;
  assign n18 = ~x0 & ~x1 ;
  assign n19 = ~x8 & n18 ;
  assign n20 = x2 & x5 ;
  assign n21 = x9 & n20 ;
  assign n22 = n19 & n21 ;
  assign n23 = n17 & n22 ;
  assign n24 = x6 & x7 ;
  assign n25 = x3 & n24 ;
  assign n26 = ~x5 & n25 ;
  assign n27 = x0 & x1 ;
  assign n28 = ~x2 & n27 ;
  assign n29 = n26 & n28 ;
  assign n30 = ~n23 & ~n29 ;
  assign n31 = x4 & x13 ;
  assign n32 = ~n30 & n31 ;
  assign n33 = n32 ^ x14 ;
  assign n34 = n33 ^ n32 ;
  assign n35 = n34 ^ x11 ;
  assign n36 = ~x10 & ~x13 ;
  assign n37 = x2 & x4 ;
  assign n38 = n36 & n37 ;
  assign n39 = n26 & n38 ;
  assign n40 = x0 & ~x1 ;
  assign n41 = x9 ^ x8 ;
  assign n42 = n40 & ~n41 ;
  assign n43 = n39 & n42 ;
  assign n44 = ~x8 & ~x9 ;
  assign n45 = x13 & n44 ;
  assign n46 = x3 & n18 ;
  assign n47 = n45 & n46 ;
  assign n48 = n27 & n36 ;
  assign n49 = x8 & x9 ;
  assign n50 = ~x3 & n49 ;
  assign n51 = n48 & n50 ;
  assign n52 = ~n47 & ~n51 ;
  assign n53 = n20 & n24 ;
  assign n54 = ~n52 & n53 ;
  assign n55 = ~x10 & x13 ;
  assign n56 = ~x2 & ~x3 ;
  assign n57 = ~x9 & n56 ;
  assign n58 = n55 & n57 ;
  assign n59 = n58 ^ x7 ;
  assign n60 = n59 ^ n58 ;
  assign n61 = x3 & x10 ;
  assign n62 = x2 & n61 ;
  assign n63 = ~x13 & n62 ;
  assign n64 = n63 ^ n58 ;
  assign n65 = n60 & n64 ;
  assign n66 = n65 ^ n58 ;
  assign n67 = n19 & n66 ;
  assign n68 = n67 ^ x6 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = n49 ^ x3 ;
  assign n71 = n70 ^ n49 ;
  assign n77 = n71 ^ n70 ;
  assign n74 = n70 ^ x7 ;
  assign n78 = n77 ^ n74 ;
  assign n79 = n78 ^ n74 ;
  assign n80 = n70 ^ x2 ;
  assign n81 = n80 ^ n74 ;
  assign n82 = n79 & ~n81 ;
  assign n72 = n70 ^ x9 ;
  assign n73 = n72 ^ n71 ;
  assign n75 = n74 ^ n73 ;
  assign n76 = ~n71 & n75 ;
  assign n83 = n82 ^ n76 ;
  assign n84 = n83 ^ n71 ;
  assign n85 = n76 ^ n74 ;
  assign n86 = n85 ^ n78 ;
  assign n87 = n74 & n86 ;
  assign n88 = n87 ^ n76 ;
  assign n89 = ~n84 & n88 ;
  assign n90 = n89 ^ n82 ;
  assign n91 = n90 ^ n87 ;
  assign n92 = n91 ^ n71 ;
  assign n93 = n92 ^ n74 ;
  assign n94 = n93 ^ n78 ;
  assign n95 = n94 ^ x3 ;
  assign n96 = n48 & n95 ;
  assign n97 = n96 ^ n67 ;
  assign n98 = n69 & n97 ;
  assign n99 = n98 ^ n67 ;
  assign n100 = ~x5 & n99 ;
  assign n101 = ~n54 & ~n100 ;
  assign n102 = ~x4 & ~n101 ;
  assign n103 = n102 ^ n43 ;
  assign n104 = ~n43 & n103 ;
  assign n105 = n104 ^ n32 ;
  assign n106 = n105 ^ n43 ;
  assign n107 = n35 & n106 ;
  assign n108 = n107 ^ n104 ;
  assign n109 = n108 ^ n43 ;
  assign n110 = ~x11 & ~n109 ;
  assign n111 = n110 ^ x11 ;
  assign n112 = ~x12 & ~n111 ;
  assign y0 = n112 ;
endmodule
