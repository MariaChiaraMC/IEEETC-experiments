module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 ;
  assign n25 = ~x0 & x1 ;
  assign n26 = ~x4 & n25 ;
  assign n27 = ~x2 & n26 ;
  assign n28 = x3 & ~x5 ;
  assign n29 = n27 & ~n28 ;
  assign n30 = ~x4 & x5 ;
  assign n31 = x0 & ~x1 ;
  assign n32 = ~x2 & ~x3 ;
  assign n33 = n31 & ~n32 ;
  assign n34 = n30 & n33 ;
  assign n35 = x1 ^ x0 ;
  assign n36 = x4 ^ x1 ;
  assign n37 = n36 ^ x4 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = ~x9 & ~x10 ;
  assign n40 = ~x8 & x11 ;
  assign n41 = n39 & n40 ;
  assign n42 = x10 & ~x11 ;
  assign n43 = x8 & n42 ;
  assign n44 = ~x12 & ~x13 ;
  assign n45 = x9 & n44 ;
  assign n46 = n43 & n45 ;
  assign n47 = ~n41 & ~n46 ;
  assign n48 = n47 ^ x3 ;
  assign n49 = ~x3 & n48 ;
  assign n50 = n49 ^ x4 ;
  assign n51 = n50 ^ x3 ;
  assign n52 = ~n38 & ~n51 ;
  assign n53 = n52 ^ n49 ;
  assign n54 = n53 ^ x3 ;
  assign n55 = n35 & ~n54 ;
  assign n56 = x2 & n55 ;
  assign n58 = ~x6 & ~x7 ;
  assign n59 = ~x8 & n58 ;
  assign n60 = ~x11 & n59 ;
  assign n57 = n27 & n45 ;
  assign n61 = n60 ^ n57 ;
  assign n62 = ~x10 & x11 ;
  assign n63 = x8 & n58 ;
  assign n64 = n62 & n63 ;
  assign n65 = n64 ^ n57 ;
  assign n66 = n65 ^ n64 ;
  assign n67 = ~x3 & n44 ;
  assign n68 = x2 & n31 ;
  assign n69 = n68 ^ x10 ;
  assign n70 = n68 ^ x9 ;
  assign n71 = n70 ^ x9 ;
  assign n72 = n26 ^ x9 ;
  assign n73 = ~n71 & ~n72 ;
  assign n74 = n73 ^ x9 ;
  assign n75 = n69 & n74 ;
  assign n76 = n75 ^ x10 ;
  assign n77 = n67 & n76 ;
  assign n78 = n77 ^ n64 ;
  assign n79 = ~n66 & ~n78 ;
  assign n80 = n79 ^ n64 ;
  assign n81 = n61 & n80 ;
  assign n82 = n81 ^ n60 ;
  assign n83 = ~n56 & ~n82 ;
  assign n84 = ~x3 & ~x4 ;
  assign n85 = x2 & ~n84 ;
  assign n86 = x13 & n41 ;
  assign n87 = n41 & n58 ;
  assign n88 = ~n43 & ~n60 ;
  assign n89 = ~x13 & ~n39 ;
  assign n90 = ~n88 & n89 ;
  assign n91 = ~n87 & ~n90 ;
  assign n92 = ~x9 & ~n59 ;
  assign n93 = ~x12 & ~n92 ;
  assign n94 = ~n91 & n93 ;
  assign n95 = ~n86 & ~n94 ;
  assign n96 = ~x4 & ~n95 ;
  assign n97 = x15 ^ x6 ;
  assign n98 = ~x9 & ~n97 ;
  assign n99 = n98 ^ x6 ;
  assign n100 = ~x12 & ~n99 ;
  assign n101 = ~x13 & ~n100 ;
  assign n102 = x8 & ~n101 ;
  assign n103 = x9 & x13 ;
  assign n104 = ~x17 & ~n103 ;
  assign n105 = x18 ^ x6 ;
  assign n106 = n105 ^ x6 ;
  assign n107 = x12 ^ x6 ;
  assign n108 = n107 ^ x6 ;
  assign n109 = n106 & ~n108 ;
  assign n110 = n109 ^ x6 ;
  assign n111 = x7 & ~n110 ;
  assign n112 = n111 ^ x6 ;
  assign n113 = n104 & ~n112 ;
  assign n114 = ~n102 & n113 ;
  assign n115 = x12 ^ x10 ;
  assign n116 = n115 ^ x7 ;
  assign n117 = x16 ^ x15 ;
  assign n118 = x10 & ~n117 ;
  assign n119 = n118 ^ x16 ;
  assign n120 = ~n116 & ~n119 ;
  assign n121 = n120 ^ n118 ;
  assign n122 = n121 ^ x16 ;
  assign n123 = n122 ^ x10 ;
  assign n124 = ~x7 & ~n123 ;
  assign n125 = ~x11 & ~n124 ;
  assign n126 = x10 & ~x12 ;
  assign n127 = ~x7 & ~n126 ;
  assign n128 = ~x9 & ~n127 ;
  assign n129 = ~n125 & ~n128 ;
  assign n130 = n114 & n129 ;
  assign n133 = ~x12 & n40 ;
  assign n134 = ~x13 & ~n133 ;
  assign n131 = ~x10 & x13 ;
  assign n132 = ~x15 & n131 ;
  assign n135 = n134 ^ n132 ;
  assign n136 = n135 ^ n134 ;
  assign n137 = n134 ^ n44 ;
  assign n138 = n137 ^ n134 ;
  assign n139 = ~n136 & ~n138 ;
  assign n140 = n139 ^ n134 ;
  assign n141 = x16 & ~n140 ;
  assign n142 = n141 ^ n134 ;
  assign n143 = n130 & n142 ;
  assign n144 = ~x3 & ~n143 ;
  assign n145 = ~n96 & ~n144 ;
  assign n146 = ~x1 & n145 ;
  assign n147 = n85 & ~n146 ;
  assign n149 = x1 & x13 ;
  assign n150 = x9 & x11 ;
  assign n151 = n126 & n150 ;
  assign n152 = ~n149 & ~n151 ;
  assign n148 = x2 & ~x22 ;
  assign n153 = n152 ^ n148 ;
  assign n154 = ~x4 & n153 ;
  assign n155 = n154 ^ n152 ;
  assign n156 = ~n25 & n155 ;
  assign n157 = ~x3 & ~n156 ;
  assign n158 = ~x10 & ~x11 ;
  assign n159 = x9 & n158 ;
  assign n160 = ~x8 & n159 ;
  assign n161 = x12 & ~n160 ;
  assign n162 = x13 & ~n161 ;
  assign n163 = n32 & n162 ;
  assign n164 = ~n157 & ~n163 ;
  assign n165 = ~x0 & ~x2 ;
  assign n166 = n165 ^ x4 ;
  assign n167 = n166 ^ n165 ;
  assign n168 = x2 & n45 ;
  assign n169 = n64 & n168 ;
  assign n170 = n169 ^ n165 ;
  assign n171 = ~n167 & ~n170 ;
  assign n172 = n171 ^ n165 ;
  assign n173 = x3 & n172 ;
  assign n174 = n173 ^ x4 ;
  assign n175 = x3 ^ x0 ;
  assign n176 = x9 & n133 ;
  assign n177 = n176 ^ x3 ;
  assign n178 = n177 ^ n176 ;
  assign n179 = n178 ^ n175 ;
  assign n180 = x21 ^ x2 ;
  assign n181 = ~x21 & n180 ;
  assign n182 = n181 ^ n176 ;
  assign n183 = n182 ^ x21 ;
  assign n184 = ~n179 & n183 ;
  assign n185 = n184 ^ n181 ;
  assign n186 = n185 ^ x21 ;
  assign n187 = ~n175 & ~n186 ;
  assign n188 = n187 ^ x3 ;
  assign n189 = n174 & n188 ;
  assign n190 = n189 ^ x1 ;
  assign n191 = n190 ^ n189 ;
  assign n192 = x3 & ~x4 ;
  assign n193 = x11 ^ x10 ;
  assign n194 = n44 & n193 ;
  assign n195 = n59 & n194 ;
  assign n196 = ~n45 & ~n195 ;
  assign n197 = ~n86 & n196 ;
  assign n198 = n192 & ~n197 ;
  assign n199 = n198 ^ n189 ;
  assign n200 = n191 & ~n199 ;
  assign n201 = n200 ^ n189 ;
  assign n202 = n164 & n201 ;
  assign n203 = ~n147 & n202 ;
  assign n204 = n203 ^ x5 ;
  assign n205 = n204 ^ n203 ;
  assign n206 = ~x4 & ~n169 ;
  assign n207 = n31 & ~n206 ;
  assign n213 = ~n60 & ~n64 ;
  assign n214 = ~n43 & n213 ;
  assign n225 = x2 & ~n64 ;
  assign n226 = x9 & ~n225 ;
  assign n227 = ~n214 & n226 ;
  assign n228 = n59 & n165 ;
  assign n229 = n42 & n228 ;
  assign n230 = ~n227 & ~n229 ;
  assign n208 = x4 ^ x3 ;
  assign n209 = x2 & x23 ;
  assign n210 = n209 ^ x4 ;
  assign n211 = n210 ^ n209 ;
  assign n212 = n211 ^ n208 ;
  assign n215 = n214 ^ n168 ;
  assign n216 = ~n214 & ~n215 ;
  assign n217 = n216 ^ n209 ;
  assign n218 = n217 ^ n214 ;
  assign n219 = n212 & n218 ;
  assign n220 = n219 ^ n216 ;
  assign n221 = n220 ^ n214 ;
  assign n222 = ~n208 & ~n221 ;
  assign n231 = n230 ^ n222 ;
  assign n232 = n231 ^ n222 ;
  assign n223 = n222 ^ n192 ;
  assign n224 = n223 ^ n222 ;
  assign n233 = n232 ^ n224 ;
  assign n234 = n222 ^ n44 ;
  assign n235 = n234 ^ n222 ;
  assign n236 = n235 ^ n232 ;
  assign n237 = ~n232 & ~n236 ;
  assign n238 = n237 ^ n232 ;
  assign n239 = ~n233 & ~n238 ;
  assign n240 = n239 ^ n237 ;
  assign n241 = n240 ^ n222 ;
  assign n242 = n241 ^ n232 ;
  assign n243 = ~x1 & ~n242 ;
  assign n244 = n243 ^ n222 ;
  assign n245 = ~n207 & ~n244 ;
  assign n246 = n245 ^ n203 ;
  assign n247 = ~n205 & n246 ;
  assign n248 = n247 ^ n203 ;
  assign n249 = n83 & n248 ;
  assign n250 = ~x20 & ~n249 ;
  assign n251 = ~x19 & n250 ;
  assign n252 = ~n34 & ~n251 ;
  assign n253 = ~n29 & n252 ;
  assign n254 = x14 & ~n253 ;
  assign y0 = n254 ;
endmodule
