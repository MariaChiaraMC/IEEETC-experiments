module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n16 = x0 & x8 ;
  assign n17 = ~x7 & ~n16 ;
  assign n18 = ~x10 & n17 ;
  assign n19 = ~x0 & x2 ;
  assign n20 = x14 & n19 ;
  assign n21 = n20 ^ x1 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n22 ^ n18 ;
  assign n24 = x9 ^ x3 ;
  assign n25 = n24 ^ x2 ;
  assign n26 = ~n24 & n25 ;
  assign n27 = n26 ^ n20 ;
  assign n28 = n27 ^ n24 ;
  assign n29 = ~n23 & ~n28 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n30 ^ n24 ;
  assign n32 = n18 & ~n31 ;
  assign n33 = n32 ^ n18 ;
  assign y0 = n33 ;
endmodule
