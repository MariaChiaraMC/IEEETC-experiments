module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 ;
  output y0 ;
  wire n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 ;
  assign n22 = x3 ^ x2 ;
  assign n23 = x3 & ~n22 ;
  assign n24 = x1 & n23 ;
  assign n25 = n24 ^ n22 ;
  assign n32 = x0 & ~n25 ;
  assign n27 = ~x1 & ~x6 ;
  assign n28 = ~x5 & n27 ;
  assign n33 = x4 & n28 ;
  assign n19 = ~x2 & ~x3 ;
  assign n20 = x1 & ~n19 ;
  assign n34 = x7 & n20 ;
  assign n35 = ~n33 & ~n34 ;
  assign n36 = ~n32 & n35 ;
  assign n21 = x10 & n20 ;
  assign n26 = x8 & ~n25 ;
  assign n29 = x9 & n28 ;
  assign n30 = ~n26 & ~n29 ;
  assign n31 = ~n21 & n30 ;
  assign n37 = n36 ^ n31 ;
  assign n38 = n31 ^ x11 ;
  assign n39 = n38 ^ n37 ;
  assign n45 = x16 & ~x17 ;
  assign n46 = ~x14 & ~n45 ;
  assign n47 = ~x15 & ~n46 ;
  assign n48 = ~x12 & ~n47 ;
  assign n49 = ~x13 & ~n48 ;
  assign n40 = ~x16 & x17 ;
  assign n41 = x14 & ~n40 ;
  assign n42 = x15 & ~n41 ;
  assign n43 = x12 & ~n42 ;
  assign n44 = x13 & ~n43 ;
  assign n50 = n49 ^ n44 ;
  assign n51 = ~x11 & n50 ;
  assign n52 = n51 ^ n44 ;
  assign n53 = n39 & n52 ;
  assign n54 = n53 ^ n51 ;
  assign n55 = n54 ^ n44 ;
  assign n56 = n55 ^ x11 ;
  assign n57 = n37 & ~n56 ;
  assign n58 = n57 ^ n36 ;
  assign y0 = ~n58 ;
endmodule
