module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n13 = ~x3 & x4 ;
  assign n14 = x6 & n13 ;
  assign n15 = x5 & ~x9 ;
  assign n16 = ~x1 & n15 ;
  assign n17 = ~x0 & ~x7 ;
  assign n18 = ~x2 & n17 ;
  assign n19 = n16 & n18 ;
  assign n20 = ~n14 & n19 ;
  assign n12 = x7 & ~x10 ;
  assign n21 = n20 ^ n12 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n20 ^ x9 ;
  assign n24 = n23 ^ n20 ;
  assign n25 = ~n22 & ~n24 ;
  assign n26 = n25 ^ n20 ;
  assign n27 = x8 & ~n26 ;
  assign n28 = n27 ^ n20 ;
  assign y0 = n28 ;
endmodule
