module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 ;
  assign n78 = x14 ^ x10 ;
  assign n86 = n78 ^ x14 ;
  assign n77 = x14 ^ x1 ;
  assign n79 = n78 ^ n77 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = n80 ^ x14 ;
  assign n82 = n79 ^ x0 ;
  assign n83 = n82 ^ n79 ;
  assign n84 = n83 ^ n81 ;
  assign n85 = ~n81 & ~n84 ;
  assign n87 = n86 ^ n85 ;
  assign n88 = n87 ^ n81 ;
  assign n89 = n79 ^ x3 ;
  assign n90 = n89 ^ n79 ;
  assign n91 = n90 ^ n86 ;
  assign n92 = n91 ^ n81 ;
  assign n93 = ~x2 & n92 ;
  assign n94 = n93 ^ n83 ;
  assign n95 = n90 ^ x14 ;
  assign n96 = n95 ^ n83 ;
  assign n97 = n86 & n96 ;
  assign n98 = n97 ^ n86 ;
  assign n99 = n94 & n98 ;
  assign n100 = n99 ^ n90 ;
  assign n101 = n100 ^ n83 ;
  assign n102 = ~n88 & ~n101 ;
  assign n103 = n102 ^ n97 ;
  assign n104 = n103 ^ n99 ;
  assign n105 = n104 ^ x10 ;
  assign n106 = n105 ^ n86 ;
  assign n107 = ~x13 & n106 ;
  assign n16 = x9 & x12 ;
  assign n17 = x10 & ~x13 ;
  assign n18 = n16 & n17 ;
  assign n108 = n107 ^ n18 ;
  assign n109 = n108 ^ n18 ;
  assign n19 = ~x1 & x5 ;
  assign n20 = x0 & n19 ;
  assign n21 = x5 & ~x6 ;
  assign n22 = x4 & ~x5 ;
  assign n23 = ~n21 & ~n22 ;
  assign n24 = ~n20 & ~n23 ;
  assign n25 = n24 ^ x13 ;
  assign n26 = x0 & x3 ;
  assign n27 = n26 ^ x1 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = n26 ^ x6 ;
  assign n30 = ~n28 & ~n29 ;
  assign n31 = n30 ^ n26 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = ~n25 & n32 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ n26 ;
  assign n36 = n35 ^ x13 ;
  assign n37 = n24 & ~n36 ;
  assign n38 = n37 ^ n24 ;
  assign n39 = x2 & ~n38 ;
  assign n43 = x2 ^ x1 ;
  assign n40 = x1 ^ x0 ;
  assign n41 = n40 ^ x2 ;
  assign n50 = n43 ^ n41 ;
  assign n42 = n41 ^ x2 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = n44 ^ n41 ;
  assign n46 = n42 ^ x5 ;
  assign n47 = n46 ^ n42 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = ~n45 & ~n48 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = n51 ^ n45 ;
  assign n53 = n41 ^ x6 ;
  assign n54 = n49 ^ n45 ;
  assign n55 = ~n53 & ~n54 ;
  assign n56 = n55 ^ n41 ;
  assign n57 = ~n52 & n56 ;
  assign n58 = n57 ^ n41 ;
  assign n59 = n58 ^ n40 ;
  assign n60 = n59 ^ n41 ;
  assign n61 = n60 ^ x13 ;
  assign n62 = n61 ^ n60 ;
  assign n63 = n62 ^ x9 ;
  assign n64 = x4 ^ x3 ;
  assign n65 = ~x3 & ~n64 ;
  assign n66 = n65 ^ n60 ;
  assign n67 = n66 ^ x3 ;
  assign n68 = ~n63 & n67 ;
  assign n69 = n68 ^ n65 ;
  assign n70 = n69 ^ x3 ;
  assign n71 = ~x9 & ~n70 ;
  assign n72 = n71 ^ x9 ;
  assign n73 = ~n39 & ~n72 ;
  assign n74 = ~x10 & ~n73 ;
  assign n75 = n74 ^ n18 ;
  assign n76 = n75 ^ n18 ;
  assign n110 = n109 ^ n76 ;
  assign n111 = n18 ^ x12 ;
  assign n112 = n111 ^ n18 ;
  assign n113 = n112 ^ n109 ;
  assign n114 = ~n109 & n113 ;
  assign n115 = n114 ^ n109 ;
  assign n116 = n110 & ~n115 ;
  assign n117 = n116 ^ n114 ;
  assign n118 = n117 ^ n18 ;
  assign n119 = n118 ^ n109 ;
  assign n120 = ~x11 & ~n119 ;
  assign n121 = n120 ^ n18 ;
  assign y0 = n121 ;
endmodule
