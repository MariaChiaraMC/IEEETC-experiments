module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 ;
  assign n18 = ~x15 & ~x16 ;
  assign n19 = ~x4 & x6 ;
  assign n20 = n18 & n19 ;
  assign n21 = ~x12 & ~x14 ;
  assign n22 = x1 & x3 ;
  assign n23 = n21 & n22 ;
  assign n24 = n20 & n23 ;
  assign n25 = x15 & x16 ;
  assign n26 = x14 & n25 ;
  assign n27 = x12 & n26 ;
  assign n28 = ~n24 & ~n27 ;
  assign n29 = ~x11 & ~x13 ;
  assign n30 = ~n28 & n29 ;
  assign n31 = x12 ^ x11 ;
  assign n32 = n31 ^ x13 ;
  assign n33 = x14 ^ x11 ;
  assign n34 = n25 ^ x11 ;
  assign n35 = n33 & n34 ;
  assign n36 = n35 ^ x11 ;
  assign n37 = n36 ^ n31 ;
  assign n38 = n32 & ~n37 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n39 ^ x11 ;
  assign n41 = n40 ^ x13 ;
  assign n42 = n31 & ~n41 ;
  assign n43 = n42 ^ n31 ;
  assign n44 = ~n30 & ~n43 ;
  assign y0 = ~n44 ;
endmodule
