module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n9 = x2 & x6 ;
  assign n10 = ~x5 & ~n9 ;
  assign n11 = x3 & ~n10 ;
  assign n12 = x6 ^ x1 ;
  assign n13 = x1 ^ x0 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = x6 ^ x2 ;
  assign n16 = n15 ^ x2 ;
  assign n17 = x5 ^ x2 ;
  assign n18 = n16 & n17 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = n19 ^ n12 ;
  assign n21 = ~n14 & n20 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = n22 ^ x2 ;
  assign n24 = n23 ^ n13 ;
  assign n25 = n12 & ~n24 ;
  assign n26 = n25 ^ n12 ;
  assign n27 = n26 ^ x1 ;
  assign n28 = ~n11 & ~n27 ;
  assign y0 = ~n28 ;
endmodule
