module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n11 = x1 & ~x9 ;
  assign n12 = n11 ^ x9 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = ~x1 & ~x4 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = n15 ^ n11 ;
  assign n17 = n13 & ~n16 ;
  assign n18 = n17 ^ n11 ;
  assign n19 = x7 & n18 ;
  assign n20 = n19 ^ n11 ;
  assign n21 = ~x8 & n20 ;
  assign n22 = x7 ^ x1 ;
  assign n23 = n22 ^ x1 ;
  assign n24 = n23 ^ x9 ;
  assign n27 = ~x4 & ~x5 ;
  assign n28 = n27 ^ x9 ;
  assign n29 = ~x9 & ~n28 ;
  assign n25 = x8 & ~n22 ;
  assign n32 = n29 ^ n25 ;
  assign n26 = n25 ^ n24 ;
  assign n30 = n29 ^ x9 ;
  assign n31 = n26 & ~n30 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = n24 & n33 ;
  assign n35 = n34 ^ n29 ;
  assign n36 = n35 ^ n31 ;
  assign n37 = ~n21 & ~n36 ;
  assign y0 = ~n37 ;
endmodule
