module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 ;
  assign n17 = ~x6 & ~x7 ;
  assign n18 = x3 & ~x5 ;
  assign n19 = n17 & n18 ;
  assign n20 = x10 ^ x8 ;
  assign n21 = n19 & n20 ;
  assign n22 = x15 ^ x14 ;
  assign n23 = n22 ^ x13 ;
  assign n24 = x15 ^ x13 ;
  assign n25 = ~x3 & ~x11 ;
  assign n26 = ~x8 & x10 ;
  assign n27 = ~x12 & n26 ;
  assign n28 = n25 & n27 ;
  assign n29 = n28 ^ x13 ;
  assign n30 = x13 & n29 ;
  assign n31 = n30 ^ x13 ;
  assign n32 = n24 & n31 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ x13 ;
  assign n35 = n34 ^ n28 ;
  assign n36 = n23 & n35 ;
  assign n37 = ~n21 & ~n36 ;
  assign n38 = x7 ^ x6 ;
  assign n39 = x7 ^ x4 ;
  assign n40 = x7 ^ x5 ;
  assign n41 = ~x7 & ~n40 ;
  assign n42 = n41 ^ x7 ;
  assign n43 = ~n39 & ~n42 ;
  assign n44 = n43 ^ n41 ;
  assign n45 = n44 ^ x7 ;
  assign n46 = n45 ^ x5 ;
  assign n47 = ~n38 & ~n46 ;
  assign n48 = n47 ^ x7 ;
  assign n49 = ~x9 & ~n48 ;
  assign n50 = ~n37 & n49 ;
  assign n51 = x4 & n18 ;
  assign n52 = ~n17 & n51 ;
  assign n53 = ~n50 & ~n52 ;
  assign n54 = ~x0 & ~x2 ;
  assign n55 = x1 & n54 ;
  assign n56 = ~n53 & n55 ;
  assign n57 = ~x1 & ~x3 ;
  assign n58 = x0 & n57 ;
  assign n59 = ~x7 & n58 ;
  assign n60 = ~n56 & ~n59 ;
  assign y0 = ~n60 ;
endmodule
