module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 ;
  assign n9 = ~x6 & x7 ;
  assign n10 = ~x1 & n9 ;
  assign n11 = x4 & ~x5 ;
  assign n12 = ~x4 & x5 ;
  assign n13 = ~x2 & n12 ;
  assign n14 = ~n11 & ~n13 ;
  assign n15 = n10 & ~n14 ;
  assign n16 = x1 & x2 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = x6 ^ x2 ;
  assign n19 = x6 & n18 ;
  assign n20 = x1 & n19 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n11 & n21 ;
  assign n23 = x2 & n12 ;
  assign n24 = ~x6 & ~x7 ;
  assign n25 = x5 & n24 ;
  assign n26 = ~x2 & n25 ;
  assign n27 = ~x5 & x6 ;
  assign n28 = x7 & n27 ;
  assign n29 = ~x4 & n28 ;
  assign n30 = ~n26 & ~n29 ;
  assign n31 = n30 ^ x1 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = n32 ^ n23 ;
  assign n34 = x5 & ~n24 ;
  assign n35 = n34 ^ x4 ;
  assign n36 = x4 & n35 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = n37 ^ x4 ;
  assign n39 = ~n33 & ~n38 ;
  assign n40 = n39 ^ n36 ;
  assign n41 = n40 ^ x4 ;
  assign n42 = ~n23 & n41 ;
  assign n43 = n42 ^ n23 ;
  assign n44 = ~n22 & ~n43 ;
  assign n45 = n44 ^ x3 ;
  assign n46 = n45 ^ n44 ;
  assign n47 = x4 & ~x7 ;
  assign n48 = ~x2 & ~n47 ;
  assign n49 = n27 & ~n48 ;
  assign n50 = n18 ^ x7 ;
  assign n51 = n50 ^ x5 ;
  assign n52 = x7 ^ x4 ;
  assign n53 = x6 ^ x4 ;
  assign n54 = n52 & n53 ;
  assign n55 = n54 ^ x4 ;
  assign n56 = n55 ^ n50 ;
  assign n57 = n51 & ~n56 ;
  assign n58 = n57 ^ n54 ;
  assign n59 = n58 ^ x4 ;
  assign n60 = n59 ^ x5 ;
  assign n61 = n50 & ~n60 ;
  assign n62 = n61 ^ n50 ;
  assign n65 = x6 ^ x5 ;
  assign n81 = ~x4 & ~n65 ;
  assign n82 = n81 ^ x5 ;
  assign n83 = ~n25 & n82 ;
  assign n63 = ~x2 & x6 ;
  assign n68 = n63 ^ x6 ;
  assign n64 = n63 ^ x4 ;
  assign n66 = n65 ^ n64 ;
  assign n67 = n66 ^ x6 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = n64 ^ n63 ;
  assign n71 = n70 ^ x6 ;
  assign n72 = n71 ^ x6 ;
  assign n73 = ~n66 & ~n72 ;
  assign n74 = n73 ^ n66 ;
  assign n75 = ~n71 & ~n74 ;
  assign n76 = n75 ^ x6 ;
  assign n77 = ~n69 & n76 ;
  assign n78 = n77 ^ n73 ;
  assign n79 = n78 ^ x6 ;
  assign n80 = n79 ^ n68 ;
  assign n84 = n83 ^ n80 ;
  assign n85 = ~x1 & ~n84 ;
  assign n86 = n85 ^ n83 ;
  assign n87 = ~n62 & n86 ;
  assign n88 = ~n49 & n87 ;
  assign n89 = n88 ^ n44 ;
  assign n90 = ~n46 & n89 ;
  assign n91 = n90 ^ n44 ;
  assign n92 = n91 ^ n15 ;
  assign n93 = n17 & ~n92 ;
  assign n94 = n93 ^ n90 ;
  assign n95 = n94 ^ n44 ;
  assign n96 = n95 ^ n16 ;
  assign n97 = ~n15 & ~n96 ;
  assign n98 = n97 ^ n15 ;
  assign y0 = n98 ;
endmodule
