module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;
  assign n11 = x2 & ~x4 ;
  assign n12 = ~x3 & x6 ;
  assign n13 = n12 ^ x7 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n12 ^ x1 ;
  assign n16 = ~n14 & n15 ;
  assign n17 = n16 ^ n12 ;
  assign n18 = ~n11 & n17 ;
  assign n19 = ~x5 & ~n18 ;
  assign n20 = ~x8 & ~x9 ;
  assign n21 = n20 ^ x6 ;
  assign n22 = x7 ^ x5 ;
  assign n23 = n20 ^ x5 ;
  assign n24 = ~n22 & n23 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = ~n21 & ~n25 ;
  assign n27 = n26 ^ x6 ;
  assign n28 = ~n19 & ~n27 ;
  assign n31 = x2 & x8 ;
  assign n29 = x5 & ~x7 ;
  assign n30 = ~x9 & n29 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = n30 ^ x0 ;
  assign n34 = n30 ^ x3 ;
  assign n35 = n30 & n34 ;
  assign n36 = n35 ^ n30 ;
  assign n37 = n33 & n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = n38 ^ n30 ;
  assign n40 = n39 ^ x3 ;
  assign n41 = n32 & n40 ;
  assign n42 = n41 ^ n30 ;
  assign n43 = n28 & ~n42 ;
  assign y0 = n43 ;
endmodule
