// Benchmark "bdd_orig/ctrl_untilsat.pla_dbb_orig_22" written by ABC on Mon Jul 12 07:22:59 2021

module \bdd_orig/ctrl_untilsat.pla_dbb_orig_22  ( 
    x0, x1, x2, x3, x4, x5, x6,
    z0  );
  input  x0, x1, x2, x3, x4, x5, x6;
  output z0;
  wire new_n9_, new_n10_, new_n11_, new_n12_, new_n13_, new_n14_, new_n15_,
    new_n16_;
  assign new_n9_ = x0 & x1;
  assign new_n10_ = x5 & x6;
  assign new_n11_ = x4 & ~new_n10_;
  assign new_n12_ = ~x2 & ~new_n11_;
  assign new_n13_ = new_n9_ & ~new_n12_;
  assign new_n14_ = x2 & x4;
  assign new_n15_ = ~new_n9_ & ~new_n14_;
  assign new_n16_ = x3 & ~new_n15_;
  assign z0 = ~new_n13_ & new_n16_;
endmodule


