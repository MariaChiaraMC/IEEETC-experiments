module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 ;
  assign n33 = ~x30 & ~x31 ;
  assign n34 = ~x28 & ~x29 ;
  assign n35 = n33 & n34 ;
  assign n36 = ~x24 & ~x27 ;
  assign n37 = ~x25 & ~x26 ;
  assign n38 = n36 & n37 ;
  assign n39 = ~n35 & n38 ;
  assign n40 = ~x22 & ~x23 ;
  assign n41 = ~x20 & n40 ;
  assign n42 = ~x21 & n41 ;
  assign n43 = ~n39 & n42 ;
  assign n44 = ~x17 & ~x18 ;
  assign n45 = ~x16 & n44 ;
  assign n46 = ~x19 & n45 ;
  assign n47 = ~n43 & n46 ;
  assign n48 = ~x12 & ~x15 ;
  assign n49 = ~x13 & n48 ;
  assign n50 = ~x14 & n49 ;
  assign n51 = ~n47 & n50 ;
  assign n52 = ~x8 & ~x11 ;
  assign n53 = ~x9 & n52 ;
  assign n54 = ~x10 & n53 ;
  assign n55 = ~n51 & n54 ;
  assign n56 = ~x4 & ~x7 ;
  assign n57 = ~x5 & n56 ;
  assign n58 = ~x6 & n57 ;
  assign n59 = ~n55 & n58 ;
  assign n60 = ~x1 & ~x2 ;
  assign n61 = ~x0 & n60 ;
  assign n62 = ~x3 & n61 ;
  assign n63 = ~n59 & n62 ;
  assign y0 = n63 ;
endmodule
