module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 ;
  assign n9 = ~x1 & ~x3 ;
  assign n10 = x4 & ~n9 ;
  assign n11 = x4 ^ x3 ;
  assign n17 = n11 ^ x4 ;
  assign n12 = n11 ^ x5 ;
  assign n13 = n12 ^ x4 ;
  assign n14 = x6 ^ x5 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = n13 & ~n15 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = x7 ^ x4 ;
  assign n21 = n16 ^ n13 ;
  assign n22 = n20 & n21 ;
  assign n23 = n22 ^ x4 ;
  assign n24 = ~n19 & ~n23 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = n25 ^ x3 ;
  assign n27 = n26 ^ x4 ;
  assign n28 = n27 ^ x1 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = ~x3 & ~x5 ;
  assign n31 = ~x6 & n30 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = n29 & ~n32 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = ~n10 & ~n34 ;
  assign n36 = x2 & ~n35 ;
  assign n37 = ~x4 & x5 ;
  assign n38 = ~x7 & n37 ;
  assign n39 = ~x3 & n38 ;
  assign n40 = x4 & ~x6 ;
  assign n41 = ~x6 & ~x7 ;
  assign n42 = n9 & n41 ;
  assign n43 = ~n40 & ~n42 ;
  assign n44 = ~n39 & n43 ;
  assign n45 = x3 & ~n41 ;
  assign n46 = ~x4 & x7 ;
  assign n47 = x6 & n46 ;
  assign n48 = ~n45 & ~n47 ;
  assign n49 = ~x5 & ~n48 ;
  assign n50 = x1 & ~n31 ;
  assign n51 = ~x2 & ~n50 ;
  assign n52 = ~n49 & n51 ;
  assign n53 = n44 & n52 ;
  assign n54 = ~x0 & ~n53 ;
  assign n55 = ~n36 & n54 ;
  assign y0 = n55 ;
endmodule
