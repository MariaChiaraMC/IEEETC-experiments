// Benchmark "./pla/newapla.pla_dbb_orig_3NonExact" written by ABC on Fri Nov 20 10:25:37 2020

module \./pla/newapla.pla_dbb_orig_3NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = ~x0;
endmodule


