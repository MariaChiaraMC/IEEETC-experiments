module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 ;
  assign n18 = ~x7 & x10 ;
  assign n19 = ~x16 & n18 ;
  assign n20 = ~x11 & ~x12 ;
  assign n21 = ~n19 & n20 ;
  assign n26 = ~x13 & ~x15 ;
  assign n22 = x15 & x16 ;
  assign n27 = n26 ^ n22 ;
  assign n23 = n22 ^ x14 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ x11 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = n29 ^ x12 ;
  assign n31 = n30 ^ n29 ;
  assign n34 = n26 ^ n24 ;
  assign n35 = n34 ^ n27 ;
  assign n36 = n35 ^ n29 ;
  assign n37 = ~n29 & n36 ;
  assign n32 = n24 & ~n27 ;
  assign n40 = n37 ^ n32 ;
  assign n33 = n32 ^ n31 ;
  assign n38 = n37 ^ n29 ;
  assign n39 = ~n33 & ~n38 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = ~n31 & n41 ;
  assign n43 = n42 ^ n37 ;
  assign n44 = n43 ^ n39 ;
  assign n45 = n44 ^ n23 ;
  assign n46 = ~n21 & n45 ;
  assign y0 = n46 ;
endmodule
