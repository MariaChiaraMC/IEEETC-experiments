module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 ;
  assign n18 = ~x3 & ~x4 ;
  assign n19 = x14 & ~x15 ;
  assign n20 = ~n18 & ~n19 ;
  assign n21 = x1 & ~n20 ;
  assign n22 = x3 & x4 ;
  assign n23 = ~x1 & x4 ;
  assign n24 = ~x11 & n23 ;
  assign n25 = ~n22 & ~n24 ;
  assign n26 = n25 ^ x3 ;
  assign n27 = ~x14 & x15 ;
  assign n28 = ~x6 & ~x7 ;
  assign n29 = ~x16 & ~n28 ;
  assign n30 = n27 & ~n29 ;
  assign n31 = x12 ^ x4 ;
  assign n32 = n19 & ~n31 ;
  assign n33 = n32 ^ x4 ;
  assign n34 = ~n30 & ~n33 ;
  assign n35 = x13 & ~n34 ;
  assign n36 = x14 & x16 ;
  assign n37 = ~x11 & ~n36 ;
  assign n38 = x12 & ~x15 ;
  assign n39 = ~x11 & x13 ;
  assign n40 = n38 & n39 ;
  assign n41 = ~n37 & ~n40 ;
  assign n42 = ~n35 & ~n41 ;
  assign n43 = x13 ^ x4 ;
  assign n44 = ~x11 & n43 ;
  assign n45 = n44 ^ x4 ;
  assign n46 = ~x12 & ~n45 ;
  assign n47 = ~n42 & ~n46 ;
  assign n48 = n47 ^ n25 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = n49 ^ n26 ;
  assign n51 = x6 ^ x5 ;
  assign n52 = x8 & x10 ;
  assign n53 = ~x16 & n52 ;
  assign n54 = x9 & n53 ;
  assign n55 = x12 ^ x11 ;
  assign n56 = n55 ^ n53 ;
  assign n57 = x14 ^ x13 ;
  assign n58 = x11 & n57 ;
  assign n59 = n58 ^ n54 ;
  assign n60 = ~n56 & n59 ;
  assign n61 = n60 ^ n58 ;
  assign n62 = n54 & n61 ;
  assign n63 = n62 ^ x6 ;
  assign n64 = n63 ^ n62 ;
  assign n65 = n64 ^ n51 ;
  assign n66 = x16 ^ x14 ;
  assign n67 = ~x16 & n66 ;
  assign n68 = n67 ^ n62 ;
  assign n69 = n68 ^ x16 ;
  assign n70 = ~n65 & n69 ;
  assign n71 = n70 ^ n67 ;
  assign n72 = n71 ^ x16 ;
  assign n73 = n51 & ~n72 ;
  assign n74 = n73 ^ x5 ;
  assign n75 = ~x7 & ~n74 ;
  assign n76 = n75 ^ x1 ;
  assign n77 = ~x1 & n76 ;
  assign n78 = n77 ^ n47 ;
  assign n79 = n78 ^ x1 ;
  assign n80 = ~n50 & n79 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n81 ^ x1 ;
  assign n83 = n26 & ~n82 ;
  assign n84 = n83 ^ n25 ;
  assign n85 = ~n21 & n84 ;
  assign n86 = x0 & ~n85 ;
  assign n87 = ~x2 & ~n86 ;
  assign n88 = x1 ^ x0 ;
  assign n89 = ~x12 & ~x13 ;
  assign n90 = x15 ^ x14 ;
  assign n91 = ~n89 & ~n90 ;
  assign n92 = x3 & ~n91 ;
  assign n93 = n92 ^ x1 ;
  assign n94 = n93 ^ n92 ;
  assign n95 = ~x5 & n28 ;
  assign n96 = n95 ^ x13 ;
  assign n97 = n96 ^ x13 ;
  assign n98 = ~x9 & ~x10 ;
  assign n99 = ~x8 & n98 ;
  assign n100 = n99 ^ x13 ;
  assign n101 = n100 ^ x13 ;
  assign n102 = ~n97 & ~n101 ;
  assign n103 = n102 ^ x13 ;
  assign n104 = x3 & n103 ;
  assign n105 = n104 ^ x13 ;
  assign n106 = n105 ^ n92 ;
  assign n107 = n94 & n106 ;
  assign n108 = n107 ^ n92 ;
  assign n109 = ~n88 & ~n108 ;
  assign n110 = n109 ^ x0 ;
  assign n111 = x4 ^ x3 ;
  assign n112 = ~n110 & n111 ;
  assign n113 = n87 & ~n112 ;
  assign n114 = ~x13 & n38 ;
  assign n115 = ~n19 & ~n57 ;
  assign n116 = ~x16 & ~n115 ;
  assign n117 = ~n114 & ~n116 ;
  assign n118 = n18 & ~n117 ;
  assign n119 = ~x12 & x15 ;
  assign n120 = x13 & n119 ;
  assign n121 = n120 ^ x3 ;
  assign n122 = n121 ^ x3 ;
  assign n123 = n22 ^ x3 ;
  assign n124 = n123 ^ x3 ;
  assign n125 = n122 & n124 ;
  assign n126 = n125 ^ x3 ;
  assign n127 = x0 & ~n126 ;
  assign n128 = n127 ^ x3 ;
  assign n129 = ~n118 & n128 ;
  assign n130 = ~x1 & ~n129 ;
  assign n131 = x14 & x15 ;
  assign n132 = ~x1 & x3 ;
  assign n133 = ~n18 & ~n132 ;
  assign n136 = n133 ^ n23 ;
  assign n137 = n136 ^ n133 ;
  assign n134 = n133 ^ x12 ;
  assign n135 = n134 ^ n133 ;
  assign n138 = n137 ^ n135 ;
  assign n139 = n133 ^ x3 ;
  assign n140 = n139 ^ n133 ;
  assign n141 = n140 ^ n137 ;
  assign n142 = n137 & n141 ;
  assign n143 = n142 ^ n137 ;
  assign n144 = n138 & n143 ;
  assign n145 = n144 ^ n142 ;
  assign n146 = n145 ^ n133 ;
  assign n147 = n146 ^ n137 ;
  assign n148 = x0 & n147 ;
  assign n149 = n148 ^ n133 ;
  assign n150 = ~n131 & n149 ;
  assign n151 = x2 & ~n150 ;
  assign n152 = ~n130 & n151 ;
  assign n153 = ~n113 & ~n152 ;
  assign y0 = n153 ;
endmodule
