module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 ;
  assign n33 = x2 ^ x0 ;
  assign n34 = n33 ^ x4 ;
  assign n31 = x3 ^ x1 ;
  assign n45 = n31 ^ x4 ;
  assign n35 = n34 ^ x2 ;
  assign n36 = n35 ^ x4 ;
  assign n46 = n45 ^ n36 ;
  assign n32 = n31 ^ x3 ;
  assign n37 = n36 ^ n32 ;
  assign n38 = n37 ^ n31 ;
  assign n47 = n46 ^ n38 ;
  assign n48 = n47 ^ n31 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n39 ^ n34 ;
  assign n49 = n48 ^ n40 ;
  assign n50 = n49 ^ n34 ;
  assign n51 = n34 & ~n50 ;
  assign n52 = n51 ^ n38 ;
  assign n53 = n52 ^ n40 ;
  assign n54 = n53 ^ n34 ;
  assign n55 = n54 ^ n31 ;
  assign n56 = n40 ^ n34 ;
  assign n57 = n56 ^ n31 ;
  assign n58 = ~n53 & ~n57 ;
  assign n59 = n58 ^ n38 ;
  assign n60 = n59 ^ n40 ;
  assign n61 = n60 ^ n34 ;
  assign n62 = n61 ^ n31 ;
  assign n63 = ~n55 & ~n62 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n41 ^ n34 ;
  assign n43 = n42 ^ n31 ;
  assign n44 = ~n42 & ~n43 ;
  assign n64 = n63 ^ n44 ;
  assign n65 = n64 ^ n51 ;
  assign n66 = n65 ^ n38 ;
  assign n67 = n66 ^ n40 ;
  assign n68 = n67 ^ n34 ;
  assign n69 = n68 ^ n31 ;
  assign n8 = x0 & x2 ;
  assign n9 = n8 ^ x3 ;
  assign n19 = n9 ^ x3 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = n19 & ~n20 ;
  assign n11 = ~x0 & ~x3 ;
  assign n12 = n11 ^ x1 ;
  assign n7 = x3 ^ x2 ;
  assign n10 = n9 ^ n7 ;
  assign n13 = n12 ^ n10 ;
  assign n14 = n13 ^ n10 ;
  assign n15 = n10 ^ n9 ;
  assign n16 = n15 ^ x3 ;
  assign n17 = ~n14 & ~n16 ;
  assign n24 = n21 ^ n17 ;
  assign n18 = n17 ^ x4 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = ~n18 & n22 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = ~x4 & n25 ;
  assign n27 = n26 ^ n17 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = n28 ^ n23 ;
  assign n30 = n29 ^ n8 ;
  assign n70 = n69 ^ n30 ;
  assign n71 = x5 & ~n70 ;
  assign n72 = n71 ^ n69 ;
  assign y0 = ~n72 ;
endmodule
