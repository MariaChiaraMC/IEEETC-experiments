// Benchmark "./pla/shift.pla_res_0NonExact" written by ABC on Fri Nov 20 10:29:14 2020

module \./pla/shift.pla_res_0NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = x0;
endmodule


