module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 ;
  assign n22 = x1 ^ x0 ;
  assign n23 = x2 ^ x1 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = x5 ^ x3 ;
  assign n27 = x5 ^ x1 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = ~n26 & ~n28 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = n30 ^ n26 ;
  assign n32 = n25 & ~n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ n26 ;
  assign n35 = n22 & ~n34 ;
  assign n36 = ~x4 & n35 ;
  assign n37 = ~x19 & ~x20 ;
  assign n38 = n37 ^ x18 ;
  assign n39 = n38 ^ x18 ;
  assign n40 = ~x1 & x3 ;
  assign n41 = x0 & ~n40 ;
  assign n42 = ~x2 & ~x11 ;
  assign n43 = ~x0 & ~x1 ;
  assign n44 = ~x9 & ~n43 ;
  assign n45 = n42 & ~n44 ;
  assign n46 = ~n41 & n45 ;
  assign n47 = ~x5 & ~n46 ;
  assign n48 = ~x9 & ~x10 ;
  assign n49 = ~x8 & n48 ;
  assign n50 = ~x8 & ~x11 ;
  assign n51 = ~n49 & ~n50 ;
  assign n52 = x12 & ~x13 ;
  assign n53 = ~x6 & ~x7 ;
  assign n54 = n53 ^ x11 ;
  assign n55 = x13 ^ x11 ;
  assign n56 = n55 ^ x11 ;
  assign n57 = n54 & ~n56 ;
  assign n58 = n57 ^ x11 ;
  assign n59 = ~x11 & n48 ;
  assign n60 = n59 ^ n52 ;
  assign n61 = ~n58 & ~n60 ;
  assign n62 = n61 ^ n59 ;
  assign n63 = ~n52 & n62 ;
  assign n64 = n63 ^ n52 ;
  assign n65 = ~n51 & ~n64 ;
  assign n66 = ~n47 & n65 ;
  assign n67 = ~x12 & ~x13 ;
  assign n68 = x9 & n67 ;
  assign n69 = x5 ^ x2 ;
  assign n85 = n69 ^ x8 ;
  assign n70 = x8 ^ x5 ;
  assign n86 = n85 ^ n70 ;
  assign n87 = n86 ^ n69 ;
  assign n88 = n87 ^ n70 ;
  assign n71 = ~x0 & ~x2 ;
  assign n72 = ~x10 & x11 ;
  assign n73 = n53 & n72 ;
  assign n74 = n71 & n73 ;
  assign n75 = ~n40 & ~n74 ;
  assign n76 = n75 ^ n70 ;
  assign n77 = n76 ^ n70 ;
  assign n89 = n77 ^ n69 ;
  assign n90 = n88 & n89 ;
  assign n78 = x10 & ~x11 ;
  assign n79 = n78 ^ n70 ;
  assign n80 = n79 ^ n76 ;
  assign n81 = n80 ^ n70 ;
  assign n82 = n81 ^ n77 ;
  assign n83 = n82 ^ n69 ;
  assign n84 = ~n69 & ~n83 ;
  assign n91 = n90 ^ n84 ;
  assign n92 = n91 ^ n87 ;
  assign n93 = n92 ^ n69 ;
  assign n94 = n93 ^ n88 ;
  assign n95 = n73 ^ n70 ;
  assign n96 = n95 ^ n69 ;
  assign n97 = n96 ^ n69 ;
  assign n98 = ~n77 & ~n97 ;
  assign n99 = n98 ^ n90 ;
  assign n100 = n99 ^ n87 ;
  assign n101 = n100 ^ n88 ;
  assign n102 = n88 & ~n101 ;
  assign n103 = n102 ^ n69 ;
  assign n104 = n103 ^ n88 ;
  assign n105 = n94 & ~n104 ;
  assign n106 = n105 ^ n84 ;
  assign n107 = n106 ^ x5 ;
  assign n108 = n68 & n107 ;
  assign n109 = ~n66 & ~n108 ;
  assign n110 = ~x4 & ~n109 ;
  assign n111 = ~n73 & ~n78 ;
  assign n112 = x8 & x9 ;
  assign n113 = ~n111 & n112 ;
  assign n114 = n50 & n53 ;
  assign n115 = ~n48 & n114 ;
  assign n116 = ~n113 & ~n115 ;
  assign n117 = ~x4 & n67 ;
  assign n118 = x2 & n117 ;
  assign n119 = ~x3 & n118 ;
  assign n120 = ~n116 & n119 ;
  assign n121 = x1 & x2 ;
  assign n122 = n121 ^ x4 ;
  assign n123 = n122 ^ x3 ;
  assign n124 = n123 ^ n122 ;
  assign n125 = n122 ^ n121 ;
  assign n126 = ~n124 & n125 ;
  assign n127 = n126 ^ n122 ;
  assign n128 = ~x0 & ~n122 ;
  assign n129 = n128 ^ x5 ;
  assign n130 = ~n127 & ~n129 ;
  assign n131 = n130 ^ n128 ;
  assign n132 = ~x5 & n131 ;
  assign n133 = n132 ^ n121 ;
  assign n134 = n133 ^ x5 ;
  assign n135 = ~n120 & n134 ;
  assign n136 = ~n43 & ~n135 ;
  assign n137 = x9 & n50 ;
  assign n138 = ~x10 & n137 ;
  assign n139 = x12 & ~n138 ;
  assign n140 = ~x2 & ~n139 ;
  assign n141 = ~x1 & ~n140 ;
  assign n142 = x13 & ~n141 ;
  assign n143 = x4 & ~n142 ;
  assign n147 = x11 ^ x8 ;
  assign n144 = x11 ^ x10 ;
  assign n148 = n147 ^ n144 ;
  assign n145 = x11 ^ x9 ;
  assign n146 = n145 ^ n144 ;
  assign n149 = n148 ^ n146 ;
  assign n152 = x11 ^ x7 ;
  assign n157 = n152 ^ n144 ;
  assign n153 = n152 ^ n148 ;
  assign n154 = n153 ^ n144 ;
  assign n155 = n154 ^ x11 ;
  assign n150 = n144 ^ x11 ;
  assign n151 = n150 ^ n149 ;
  assign n156 = n155 ^ n151 ;
  assign n158 = n157 ^ n156 ;
  assign n159 = ~n149 & ~n158 ;
  assign n160 = n159 ^ x11 ;
  assign n161 = n160 ^ n150 ;
  assign n162 = ~x16 & n151 ;
  assign n163 = n162 ^ x16 ;
  assign n164 = n163 ^ n150 ;
  assign n165 = n164 ^ n157 ;
  assign n166 = n150 ^ x11 ;
  assign n167 = n166 ^ n157 ;
  assign n168 = x11 & n167 ;
  assign n169 = n168 ^ n150 ;
  assign n170 = n169 ^ n149 ;
  assign n171 = ~n165 & n170 ;
  assign n172 = n171 ^ x11 ;
  assign n173 = n172 ^ n149 ;
  assign n174 = n173 ^ n157 ;
  assign n175 = ~n161 & n174 ;
  assign n176 = n175 ^ n171 ;
  assign n177 = n176 ^ x11 ;
  assign n178 = n177 ^ n149 ;
  assign n179 = n178 ^ x11 ;
  assign n180 = n179 ^ n157 ;
  assign n181 = ~x6 & ~x17 ;
  assign n182 = n181 ^ n180 ;
  assign n183 = x15 ^ x13 ;
  assign n184 = n183 ^ x15 ;
  assign n185 = x15 ^ x12 ;
  assign n186 = ~n184 & n185 ;
  assign n187 = n186 ^ x15 ;
  assign n188 = n187 ^ n180 ;
  assign n189 = ~n182 & n188 ;
  assign n190 = n189 ^ n186 ;
  assign n191 = n190 ^ x15 ;
  assign n192 = n191 ^ n181 ;
  assign n193 = ~n180 & ~n192 ;
  assign n194 = n193 ^ n180 ;
  assign n195 = x2 & n194 ;
  assign n196 = ~x0 & x1 ;
  assign n197 = n72 ^ x12 ;
  assign n198 = x11 ^ x2 ;
  assign n199 = n198 ^ x2 ;
  assign n200 = x9 ^ x2 ;
  assign n201 = n199 & n200 ;
  assign n202 = n201 ^ x2 ;
  assign n203 = n202 ^ n72 ;
  assign n204 = n197 & ~n203 ;
  assign n205 = n204 ^ n201 ;
  assign n206 = n205 ^ x2 ;
  assign n207 = n206 ^ x12 ;
  assign n208 = ~n72 & ~n207 ;
  assign n209 = n208 ^ n72 ;
  assign n210 = ~n196 & n209 ;
  assign n211 = ~n195 & n210 ;
  assign n212 = n143 & n211 ;
  assign n213 = x5 & ~n212 ;
  assign n214 = n71 ^ x1 ;
  assign n215 = n214 ^ x4 ;
  assign n229 = n215 ^ x0 ;
  assign n216 = n215 ^ n71 ;
  assign n217 = n216 ^ n215 ;
  assign n228 = n217 ^ x0 ;
  assign n230 = n229 ^ n228 ;
  assign n219 = ~x8 & x11 ;
  assign n220 = x5 & x9 ;
  assign n221 = n219 & n220 ;
  assign n222 = ~x12 & n221 ;
  assign n223 = n222 ^ n216 ;
  assign n218 = n217 ^ n214 ;
  assign n224 = n223 ^ n218 ;
  assign n225 = n218 ^ x0 ;
  assign n226 = n224 & n225 ;
  assign n227 = n226 ^ x0 ;
  assign n231 = n230 ^ n227 ;
  assign n232 = n231 ^ n223 ;
  assign n233 = n230 ^ n229 ;
  assign n234 = n233 ^ n218 ;
  assign n235 = n229 & n234 ;
  assign n236 = ~x8 & ~x9 ;
  assign n237 = n72 & n236 ;
  assign n238 = x2 & n237 ;
  assign n239 = n229 ^ n223 ;
  assign n240 = n238 & ~n239 ;
  assign n241 = n240 ^ n238 ;
  assign n242 = n241 ^ n223 ;
  assign n243 = n242 ^ n218 ;
  assign n244 = n235 & n243 ;
  assign n245 = n244 ^ x0 ;
  assign n246 = ~n232 & ~n245 ;
  assign n247 = n246 ^ n235 ;
  assign n248 = n247 ^ n244 ;
  assign n249 = n248 ^ x0 ;
  assign n250 = n249 ^ n229 ;
  assign n251 = n250 ^ n230 ;
  assign n252 = n251 ^ x1 ;
  assign n253 = n252 ^ n217 ;
  assign n254 = ~n213 & n253 ;
  assign n255 = n254 ^ x3 ;
  assign n256 = n255 ^ n254 ;
  assign n257 = n256 ^ n136 ;
  assign n258 = ~x2 & x5 ;
  assign n259 = n258 ^ x1 ;
  assign n260 = n258 & ~n259 ;
  assign n261 = n260 ^ n254 ;
  assign n262 = n261 ^ n258 ;
  assign n263 = ~n257 & ~n262 ;
  assign n264 = n263 ^ n260 ;
  assign n265 = n264 ^ n258 ;
  assign n266 = ~n136 & n265 ;
  assign n267 = n266 ^ n136 ;
  assign n268 = ~n110 & ~n267 ;
  assign n269 = n268 ^ x18 ;
  assign n270 = n39 & n269 ;
  assign n271 = n270 ^ x18 ;
  assign n272 = x14 & n271 ;
  assign n273 = ~n36 & n272 ;
  assign y0 = ~n273 ;
endmodule
