module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 ;
  assign n11 = x7 & x9 ;
  assign n12 = ~x1 & n11 ;
  assign n13 = ~x5 & x6 ;
  assign n14 = ~x0 & n13 ;
  assign n15 = n12 & n14 ;
  assign n17 = x3 & ~x8 ;
  assign n16 = ~x3 & x8 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = x2 & n18 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n15 & n20 ;
  assign n23 = x2 & x8 ;
  assign n24 = x6 & ~x9 ;
  assign n25 = ~x7 & n24 ;
  assign n26 = n23 & n25 ;
  assign n168 = x1 & n26 ;
  assign n169 = n168 ^ x3 ;
  assign n71 = x7 & n24 ;
  assign n171 = ~x2 & ~x5 ;
  assign n172 = n71 & n171 ;
  assign n173 = ~x7 & x9 ;
  assign n174 = x5 & ~x6 ;
  assign n175 = n173 & n174 ;
  assign n176 = ~n172 & ~n175 ;
  assign n67 = x2 & x9 ;
  assign n170 = ~x7 & n67 ;
  assign n177 = n176 ^ n170 ;
  assign n178 = n177 ^ n176 ;
  assign n179 = n176 ^ x5 ;
  assign n180 = n179 ^ n176 ;
  assign n181 = n178 & n180 ;
  assign n182 = n181 ^ n176 ;
  assign n183 = ~x1 & ~n182 ;
  assign n184 = n183 ^ n176 ;
  assign n185 = ~x8 & ~n184 ;
  assign n89 = ~x1 & x7 ;
  assign n186 = x5 ^ x2 ;
  assign n187 = x9 ^ x5 ;
  assign n188 = n187 ^ x9 ;
  assign n30 = x8 & x9 ;
  assign n189 = n30 ^ x9 ;
  assign n190 = ~n188 & ~n189 ;
  assign n191 = n190 ^ x9 ;
  assign n192 = ~n186 & ~n191 ;
  assign n193 = n89 & n192 ;
  assign n194 = ~x7 & x8 ;
  assign n195 = x5 & ~x9 ;
  assign n196 = ~n67 & ~n195 ;
  assign n197 = ~n171 & n196 ;
  assign n198 = n194 & n197 ;
  assign n199 = ~n193 & ~n198 ;
  assign n200 = n199 ^ x6 ;
  assign n201 = n200 ^ n199 ;
  assign n202 = n201 ^ n185 ;
  assign n203 = ~x1 & ~x5 ;
  assign n204 = n173 & n203 ;
  assign n114 = ~x1 & ~x9 ;
  assign n205 = x8 & n114 ;
  assign n206 = n205 ^ x5 ;
  assign n207 = n206 ^ n205 ;
  assign n68 = x7 & x8 ;
  assign n208 = ~x9 & n68 ;
  assign n209 = n208 ^ n205 ;
  assign n210 = ~n207 & n209 ;
  assign n211 = n210 ^ n205 ;
  assign n212 = ~n204 & ~n211 ;
  assign n213 = n212 ^ x2 ;
  assign n214 = ~n212 & n213 ;
  assign n215 = n214 ^ n199 ;
  assign n216 = n215 ^ n212 ;
  assign n217 = n202 & n216 ;
  assign n218 = n217 ^ n214 ;
  assign n219 = n218 ^ n212 ;
  assign n220 = ~n185 & ~n219 ;
  assign n221 = n220 ^ n185 ;
  assign n222 = n221 ^ x0 ;
  assign n223 = n222 ^ n221 ;
  assign n78 = ~x6 & n11 ;
  assign n79 = ~x8 & n78 ;
  assign n224 = x8 ^ x6 ;
  assign n225 = n224 ^ x8 ;
  assign n36 = ~x7 & ~x8 ;
  assign n226 = n36 ^ x8 ;
  assign n227 = n225 & n226 ;
  assign n228 = n227 ^ x8 ;
  assign n229 = n114 & n228 ;
  assign n230 = ~n79 & ~n229 ;
  assign n231 = n171 & ~n230 ;
  assign n62 = x6 & ~x7 ;
  assign n232 = ~x1 & x5 ;
  assign n233 = n62 & n232 ;
  assign n234 = n23 & n233 ;
  assign n34 = x2 & x7 ;
  assign n235 = ~n13 & n34 ;
  assign n236 = x9 ^ x8 ;
  assign n237 = ~x6 & n203 ;
  assign n238 = n237 ^ x9 ;
  assign n239 = n238 ^ n237 ;
  assign n240 = n239 ^ n236 ;
  assign n241 = n174 ^ x1 ;
  assign n242 = ~n174 & ~n241 ;
  assign n243 = n242 ^ n237 ;
  assign n244 = n243 ^ n174 ;
  assign n245 = ~n240 & ~n244 ;
  assign n246 = n245 ^ n242 ;
  assign n247 = n246 ^ n174 ;
  assign n248 = ~n236 & ~n247 ;
  assign n249 = n235 & n248 ;
  assign n250 = ~n234 & ~n249 ;
  assign n251 = ~n231 & n250 ;
  assign n252 = n251 ^ n221 ;
  assign n253 = ~n223 & ~n252 ;
  assign n254 = n253 ^ n221 ;
  assign n255 = n254 ^ n168 ;
  assign n256 = n169 & n255 ;
  assign n257 = n256 ^ n253 ;
  assign n258 = n257 ^ n221 ;
  assign n259 = n258 ^ x3 ;
  assign n260 = ~n168 & n259 ;
  assign n261 = n260 ^ n168 ;
  assign n112 = ~x0 & x2 ;
  assign n54 = ~x8 & x9 ;
  assign n262 = ~x7 & n54 ;
  assign n263 = ~n208 & ~n262 ;
  assign n264 = n112 & ~n263 ;
  assign n122 = ~x2 & ~x9 ;
  assign n265 = ~n68 & ~n122 ;
  assign n266 = ~n36 & ~n67 ;
  assign n267 = x0 & ~n266 ;
  assign n268 = ~n265 & n267 ;
  assign n269 = ~n264 & ~n268 ;
  assign n270 = x6 & ~n269 ;
  assign n29 = ~x2 & ~x6 ;
  assign n271 = ~x0 & n29 ;
  assign n272 = n194 & n271 ;
  assign n273 = ~x1 & ~n272 ;
  assign n274 = ~n270 & n273 ;
  assign n275 = n262 & n271 ;
  assign n276 = n79 ^ x2 ;
  assign n277 = n276 ^ n79 ;
  assign n278 = ~n24 & n194 ;
  assign n279 = n278 ^ n79 ;
  assign n280 = ~n277 & n279 ;
  assign n281 = n280 ^ n79 ;
  assign n282 = x0 & n281 ;
  assign n283 = x1 & ~n282 ;
  assign n284 = ~n275 & n283 ;
  assign n285 = ~n274 & ~n284 ;
  assign n286 = n285 ^ x5 ;
  assign n287 = n286 ^ n285 ;
  assign n288 = n287 ^ x3 ;
  assign n144 = x2 ^ x1 ;
  assign n291 = n144 ^ x9 ;
  assign n289 = x8 ^ x7 ;
  assign n292 = n291 ^ n289 ;
  assign n296 = n292 ^ n144 ;
  assign n290 = n289 ^ n144 ;
  assign n293 = n292 ^ n290 ;
  assign n294 = ~n290 & n293 ;
  assign n295 = n294 ^ n290 ;
  assign n297 = n296 ^ n295 ;
  assign n304 = x2 ^ x0 ;
  assign n305 = n304 ^ x7 ;
  assign n298 = n144 ^ x2 ;
  assign n299 = n298 ^ n296 ;
  assign n300 = n144 ^ x8 ;
  assign n301 = n300 ^ n298 ;
  assign n302 = ~n299 & ~n301 ;
  assign n303 = n302 ^ n300 ;
  assign n306 = n305 ^ n303 ;
  assign n307 = n305 ^ n299 ;
  assign n308 = ~n298 & ~n307 ;
  assign n309 = n308 ^ n298 ;
  assign n310 = n309 ^ n296 ;
  assign n311 = n306 & ~n310 ;
  assign n312 = n311 ^ n305 ;
  assign n313 = ~n297 & n312 ;
  assign n314 = n313 ^ x6 ;
  assign n315 = ~x6 & ~n314 ;
  assign n316 = n315 ^ n285 ;
  assign n317 = n316 ^ x6 ;
  assign n318 = n288 & ~n317 ;
  assign n319 = n318 ^ n315 ;
  assign n320 = n319 ^ x6 ;
  assign n321 = x3 & ~n320 ;
  assign n322 = n321 ^ x3 ;
  assign n323 = n261 & ~n322 ;
  assign n22 = ~x0 & x1 ;
  assign n27 = x3 & n26 ;
  assign n28 = n22 & n27 ;
  assign n31 = ~x1 & ~x7 ;
  assign n32 = n30 & n31 ;
  assign n33 = n29 & n32 ;
  assign n35 = x8 & n34 ;
  assign n37 = n29 & n36 ;
  assign n38 = ~n35 & ~n37 ;
  assign n39 = n38 ^ x1 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = n40 ^ x9 ;
  assign n42 = x2 & n36 ;
  assign n43 = n42 ^ x6 ;
  assign n44 = n42 & n43 ;
  assign n45 = n44 ^ n38 ;
  assign n46 = n45 ^ n42 ;
  assign n47 = ~n41 & ~n46 ;
  assign n48 = n47 ^ n44 ;
  assign n49 = n48 ^ n42 ;
  assign n50 = ~x9 & n49 ;
  assign n51 = ~n33 & ~n50 ;
  assign n52 = x0 & ~n51 ;
  assign n53 = ~x1 & ~x2 ;
  assign n55 = x6 & n54 ;
  assign n56 = n53 & n55 ;
  assign n57 = x7 & n56 ;
  assign n58 = ~n52 & ~n57 ;
  assign n59 = x3 & ~n58 ;
  assign n60 = ~x5 & ~n59 ;
  assign n61 = x2 & ~x3 ;
  assign n63 = ~x8 & ~x9 ;
  assign n64 = n62 & n63 ;
  assign n65 = n61 & n64 ;
  assign n66 = x3 & ~x6 ;
  assign n69 = n67 & n68 ;
  assign n70 = n66 & n69 ;
  assign n72 = ~n23 & n71 ;
  assign n73 = x8 ^ x3 ;
  assign n74 = n72 & n73 ;
  assign n75 = ~n70 & ~n74 ;
  assign n76 = ~n65 & n75 ;
  assign n77 = n22 & ~n76 ;
  assign n80 = n54 & n62 ;
  assign n81 = n80 ^ x3 ;
  assign n82 = n81 ^ n80 ;
  assign n83 = ~n25 & ~n78 ;
  assign n84 = n83 ^ n80 ;
  assign n85 = n82 & ~n84 ;
  assign n86 = n85 ^ n80 ;
  assign n87 = ~n79 & ~n86 ;
  assign n88 = n53 & ~n87 ;
  assign n90 = ~x3 & x6 ;
  assign n91 = n30 & n90 ;
  assign n92 = n89 & n91 ;
  assign n93 = ~n27 & ~n92 ;
  assign n94 = ~n88 & n93 ;
  assign n95 = n94 ^ x0 ;
  assign n96 = n95 ^ n94 ;
  assign n97 = n96 ^ n77 ;
  assign n98 = x2 & n31 ;
  assign n99 = ~n12 & ~n98 ;
  assign n100 = ~x3 & ~n23 ;
  assign n101 = ~n99 & n100 ;
  assign n102 = n101 ^ x6 ;
  assign n103 = ~x6 & ~n102 ;
  assign n104 = n103 ^ n94 ;
  assign n105 = n104 ^ x6 ;
  assign n106 = ~n97 & n105 ;
  assign n107 = n106 ^ n103 ;
  assign n108 = n107 ^ x6 ;
  assign n109 = ~n77 & ~n108 ;
  assign n110 = n109 ^ n77 ;
  assign n111 = n60 & ~n110 ;
  assign n113 = x6 ^ x3 ;
  assign n115 = n114 ^ x9 ;
  assign n116 = x9 ^ x6 ;
  assign n117 = n116 ^ x9 ;
  assign n118 = n115 & ~n117 ;
  assign n119 = n118 ^ x9 ;
  assign n120 = n113 & n119 ;
  assign n121 = n112 & n120 ;
  assign n123 = n66 & n122 ;
  assign n124 = x1 & n123 ;
  assign n125 = n24 & n53 ;
  assign n126 = x0 & n125 ;
  assign n127 = n22 & n67 ;
  assign n128 = n127 ^ x3 ;
  assign n129 = n126 & ~n128 ;
  assign n130 = n129 ^ n127 ;
  assign n131 = ~x3 & n130 ;
  assign n132 = ~n124 & ~n131 ;
  assign n133 = ~n121 & n132 ;
  assign n134 = n36 & ~n133 ;
  assign n135 = x5 & ~n134 ;
  assign n136 = ~x2 & n17 ;
  assign n137 = ~x1 & x2 ;
  assign n138 = n61 & ~n137 ;
  assign n139 = ~n136 & ~n138 ;
  assign n140 = x0 & ~x6 ;
  assign n141 = x9 & n140 ;
  assign n142 = ~n139 & n141 ;
  assign n143 = ~x0 & x6 ;
  assign n145 = x3 ^ x2 ;
  assign n146 = n144 & ~n145 ;
  assign n147 = n143 & n146 ;
  assign n148 = n63 & n147 ;
  assign n149 = ~n142 & ~n148 ;
  assign n150 = n149 ^ x7 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = n151 ^ n135 ;
  assign n153 = n114 ^ n22 ;
  assign n154 = x3 & n153 ;
  assign n155 = n154 ^ n114 ;
  assign n156 = n29 & n155 ;
  assign n157 = n156 ^ x8 ;
  assign n158 = n156 & n157 ;
  assign n159 = n158 ^ n149 ;
  assign n160 = n159 ^ n156 ;
  assign n161 = ~n152 & ~n160 ;
  assign n162 = n161 ^ n158 ;
  assign n163 = n162 ^ n156 ;
  assign n164 = n135 & n163 ;
  assign n165 = n164 ^ n135 ;
  assign n166 = ~n111 & ~n165 ;
  assign n167 = ~n28 & ~n166 ;
  assign n324 = n323 ^ n167 ;
  assign n325 = n324 ^ n167 ;
  assign n326 = n53 & n262 ;
  assign n327 = n143 ^ n140 ;
  assign n328 = x5 & n327 ;
  assign n329 = n328 ^ n140 ;
  assign n330 = n326 & n329 ;
  assign n331 = n330 ^ n167 ;
  assign n332 = n331 ^ n167 ;
  assign n333 = ~n325 & ~n332 ;
  assign n334 = n333 ^ n167 ;
  assign n335 = x4 & n334 ;
  assign n336 = n335 ^ n167 ;
  assign n337 = ~n21 & n336 ;
  assign y0 = ~n337 ;
endmodule
