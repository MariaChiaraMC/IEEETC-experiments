module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n11 = x6 ^ x2 ;
  assign n12 = n11 ^ x0 ;
  assign n13 = ~x3 & ~x7 ;
  assign n14 = ~x4 & n13 ;
  assign n15 = ~x1 & ~x5 ;
  assign n16 = n14 & n15 ;
  assign n17 = n16 ^ n12 ;
  assign n18 = x6 ^ x0 ;
  assign n19 = x9 ^ x6 ;
  assign n20 = n19 ^ x6 ;
  assign n21 = n18 & n20 ;
  assign n22 = n21 ^ x6 ;
  assign n23 = n22 ^ n12 ;
  assign n24 = n17 & ~n23 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ x6 ;
  assign n27 = n26 ^ n16 ;
  assign n28 = n12 & ~n27 ;
  assign n29 = n28 ^ n12 ;
  assign y0 = n29 ;
endmodule
