module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 ;
  assign n9 = x3 & x5 ;
  assign n10 = x6 & x7 ;
  assign n11 = x0 & x1 ;
  assign n12 = n10 & n11 ;
  assign n13 = n9 & n12 ;
  assign n14 = ~x2 & n13 ;
  assign n40 = ~x1 & x3 ;
  assign n89 = x6 ^ x5 ;
  assign n90 = x5 ^ x0 ;
  assign n91 = ~n89 & n90 ;
  assign n92 = n89 ^ x2 ;
  assign n93 = n91 ^ n10 ;
  assign n94 = ~n92 & n93 ;
  assign n95 = n94 ^ n10 ;
  assign n96 = n91 & n95 ;
  assign n97 = n40 & n96 ;
  assign n20 = ~x0 & ~x3 ;
  assign n98 = x1 & ~n9 ;
  assign n99 = ~n20 & n98 ;
  assign n15 = ~x3 & ~x5 ;
  assign n100 = ~x2 & ~x6 ;
  assign n101 = ~n15 & n100 ;
  assign n102 = ~x7 & n101 ;
  assign n103 = n99 & n102 ;
  assign n104 = ~n97 & ~n103 ;
  assign n16 = n12 & n15 ;
  assign n54 = ~x6 & x7 ;
  assign n55 = ~x1 & n15 ;
  assign n56 = n54 & n55 ;
  assign n57 = x0 & n56 ;
  assign n36 = x0 & x6 ;
  assign n37 = ~x0 & ~x1 ;
  assign n38 = ~n36 & ~n37 ;
  assign n39 = ~x0 & ~x7 ;
  assign n41 = ~x7 & n40 ;
  assign n42 = ~n9 & ~n41 ;
  assign n43 = ~n39 & ~n42 ;
  assign n44 = ~n38 & n43 ;
  assign n45 = x5 & x6 ;
  assign n46 = ~x1 & ~n45 ;
  assign n47 = n20 & ~n46 ;
  assign n48 = x5 & ~x6 ;
  assign n49 = n48 ^ x7 ;
  assign n50 = n47 & ~n49 ;
  assign n51 = ~n44 & ~n50 ;
  assign n58 = n57 ^ n51 ;
  assign n59 = n58 ^ n51 ;
  assign n17 = x7 ^ x6 ;
  assign n18 = x7 ^ x3 ;
  assign n19 = n18 ^ x3 ;
  assign n21 = n20 ^ x3 ;
  assign n22 = n19 & n21 ;
  assign n23 = n22 ^ x3 ;
  assign n24 = n17 & n23 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n26 ^ x1 ;
  assign n28 = n10 ^ x0 ;
  assign n29 = ~n10 & ~n28 ;
  assign n30 = n29 ^ n24 ;
  assign n31 = n30 ^ n10 ;
  assign n32 = n27 & ~n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ n10 ;
  assign n35 = x1 & ~n34 ;
  assign n52 = n51 ^ n35 ;
  assign n53 = n52 ^ n51 ;
  assign n60 = n59 ^ n53 ;
  assign n61 = ~x5 & n10 ;
  assign n62 = ~x7 & n48 ;
  assign n63 = ~n61 & ~n62 ;
  assign n64 = x3 & ~n63 ;
  assign n65 = x6 & ~x7 ;
  assign n66 = n15 & n65 ;
  assign n67 = ~n64 & ~n66 ;
  assign n68 = n37 & ~n67 ;
  assign n69 = n68 ^ n51 ;
  assign n70 = n69 ^ n51 ;
  assign n71 = n70 ^ n59 ;
  assign n72 = ~n59 & n71 ;
  assign n73 = n72 ^ n59 ;
  assign n74 = n60 & ~n73 ;
  assign n75 = n74 ^ n72 ;
  assign n76 = n75 ^ n51 ;
  assign n77 = n76 ^ n59 ;
  assign n78 = x2 & ~n77 ;
  assign n79 = n78 ^ n51 ;
  assign n80 = ~n16 & n79 ;
  assign n105 = n104 ^ n80 ;
  assign n106 = n105 ^ n80 ;
  assign n81 = ~x3 & x7 ;
  assign n82 = x0 & ~x2 ;
  assign n83 = ~x5 & ~x6 ;
  assign n84 = n82 & ~n83 ;
  assign n85 = n81 & n84 ;
  assign n86 = ~x1 & n85 ;
  assign n87 = n86 ^ n80 ;
  assign n88 = n87 ^ n80 ;
  assign n107 = n106 ^ n88 ;
  assign n108 = n98 ^ n48 ;
  assign n109 = n98 ^ x3 ;
  assign n110 = n109 ^ n98 ;
  assign n111 = n110 ^ n108 ;
  assign n112 = n36 ^ x1 ;
  assign n113 = ~n98 & ~n112 ;
  assign n114 = n113 ^ n36 ;
  assign n115 = n111 & n114 ;
  assign n116 = n115 ^ n113 ;
  assign n117 = n116 ^ n36 ;
  assign n118 = n117 ^ n98 ;
  assign n119 = n108 & ~n118 ;
  assign n120 = n119 ^ n48 ;
  assign n123 = n120 ^ x0 ;
  assign n124 = n123 ^ n120 ;
  assign n121 = n120 ^ n40 ;
  assign n122 = n121 ^ n120 ;
  assign n125 = n124 ^ n122 ;
  assign n126 = x3 ^ x1 ;
  assign n127 = ~x5 & ~n126 ;
  assign n128 = n127 ^ x1 ;
  assign n129 = n128 ^ n120 ;
  assign n130 = n129 ^ n120 ;
  assign n131 = n130 ^ n124 ;
  assign n132 = ~n124 & n131 ;
  assign n133 = n132 ^ n124 ;
  assign n134 = n125 & ~n133 ;
  assign n135 = n134 ^ n132 ;
  assign n136 = n135 ^ n120 ;
  assign n137 = n136 ^ n124 ;
  assign n138 = ~x7 & ~n137 ;
  assign n139 = n138 ^ n120 ;
  assign n140 = x2 & n139 ;
  assign n141 = n140 ^ n80 ;
  assign n142 = n141 ^ n80 ;
  assign n143 = n142 ^ n106 ;
  assign n144 = n106 & ~n143 ;
  assign n145 = n144 ^ n106 ;
  assign n146 = ~n107 & n145 ;
  assign n147 = n146 ^ n144 ;
  assign n148 = n147 ^ n80 ;
  assign n149 = n148 ^ n106 ;
  assign n150 = x4 & n149 ;
  assign n151 = n150 ^ n80 ;
  assign n152 = ~n14 & n151 ;
  assign y0 = ~n152 ;
endmodule
