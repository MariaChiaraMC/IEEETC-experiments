module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 ;
  assign n19 = ~x9 & ~x11 ;
  assign n20 = x10 & n19 ;
  assign n21 = x7 ^ x6 ;
  assign n22 = x7 ^ x4 ;
  assign n23 = x7 ^ x5 ;
  assign n24 = ~x7 & ~n23 ;
  assign n25 = n24 ^ x7 ;
  assign n26 = ~n22 & ~n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n27 ^ x7 ;
  assign n29 = n28 ^ x5 ;
  assign n30 = ~n21 & ~n29 ;
  assign n31 = n30 ^ x7 ;
  assign n32 = n20 & ~n31 ;
  assign n33 = ~x3 & ~x12 ;
  assign n34 = x13 & x15 ;
  assign n35 = ~x8 & ~n34 ;
  assign n36 = ~x13 & ~x15 ;
  assign n37 = n36 ^ x14 ;
  assign n38 = n35 & ~n37 ;
  assign n39 = n33 & n38 ;
  assign n40 = n32 & n39 ;
  assign n41 = ~x6 & ~x7 ;
  assign n42 = x3 & x4 ;
  assign n43 = ~x5 & n42 ;
  assign n44 = ~n41 & n43 ;
  assign n45 = ~n40 & ~n44 ;
  assign n17 = x0 & ~x7 ;
  assign n18 = ~x3 & n17 ;
  assign n46 = n45 ^ n18 ;
  assign n47 = n46 ^ n18 ;
  assign n48 = ~x0 & ~x2 ;
  assign n49 = n48 ^ n18 ;
  assign n50 = n49 ^ n18 ;
  assign n51 = ~n47 & n50 ;
  assign n52 = n51 ^ n18 ;
  assign n53 = x1 & n52 ;
  assign n54 = n53 ^ n18 ;
  assign y0 = n54 ;
endmodule
