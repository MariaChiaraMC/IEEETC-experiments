module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 ;
  assign n18 = x3 ^ x2 ;
  assign n16 = x3 ^ x1 ;
  assign n25 = n18 ^ n16 ;
  assign n17 = n16 ^ x3 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = n17 ^ x4 ;
  assign n22 = n21 ^ n17 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n20 & n23 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n26 ^ n20 ;
  assign n28 = n16 ^ x5 ;
  assign n29 = n24 ^ n20 ;
  assign n30 = ~n28 & n29 ;
  assign n31 = n30 ^ n16 ;
  assign n32 = n27 & n31 ;
  assign n33 = n32 ^ n16 ;
  assign n34 = n33 ^ x1 ;
  assign n35 = n34 ^ n16 ;
  assign n36 = ~x0 & n35 ;
  assign y0 = n36 ;
endmodule
