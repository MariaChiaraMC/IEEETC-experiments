module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 ;
  output y0 ;
  wire n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 ;
  assign n23 = ~x0 & ~x1 ;
  assign n24 = ~x4 & ~n23 ;
  assign n25 = x1 ^ x0 ;
  assign n26 = x2 & n25 ;
  assign n27 = n26 ^ x0 ;
  assign n28 = n27 ^ x5 ;
  assign n29 = n28 ^ n24 ;
  assign n30 = x5 ^ x3 ;
  assign n31 = x5 ^ x1 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = ~n30 & ~n32 ;
  assign n34 = n33 ^ x5 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = ~n29 & ~n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ n30 ;
  assign n39 = n24 & ~n38 ;
  assign n40 = ~x20 & ~x21 ;
  assign n41 = n40 ^ x19 ;
  assign n42 = n41 ^ x19 ;
  assign n43 = x2 & ~x3 ;
  assign n44 = ~x6 & x8 ;
  assign n45 = n43 & n44 ;
  assign n46 = ~x2 & ~x12 ;
  assign n47 = n46 ^ x13 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = n46 ^ x10 ;
  assign n50 = n48 & ~n49 ;
  assign n51 = n50 ^ x10 ;
  assign n61 = ~x8 & x9 ;
  assign n62 = ~x11 & n61 ;
  assign n54 = x11 & ~x12 ;
  assign n52 = n46 ^ x9 ;
  assign n53 = n52 ^ n47 ;
  assign n55 = n54 ^ n53 ;
  assign n56 = n55 ^ n53 ;
  assign n57 = n53 ^ n47 ;
  assign n58 = n57 ^ n46 ;
  assign n59 = n58 ^ n50 ;
  assign n60 = n56 & n59 ;
  assign n63 = n62 ^ n60 ;
  assign n64 = ~x10 & n63 ;
  assign n65 = n64 ^ n60 ;
  assign n66 = n65 ^ n48 ;
  assign n67 = ~n51 & n66 ;
  assign n68 = n67 ^ n60 ;
  assign n69 = n68 ^ n64 ;
  assign n70 = n69 ^ n48 ;
  assign n71 = n70 ^ x13 ;
  assign n72 = x4 & n71 ;
  assign n73 = x2 ^ x1 ;
  assign n74 = x0 & ~x13 ;
  assign n75 = n74 ^ x2 ;
  assign n76 = n75 ^ n74 ;
  assign n77 = n76 ^ n73 ;
  assign n78 = x15 ^ x12 ;
  assign n79 = x13 & n78 ;
  assign n80 = n79 ^ x12 ;
  assign n81 = ~x17 & ~n80 ;
  assign n82 = ~x13 & ~x18 ;
  assign n83 = x9 & ~n82 ;
  assign n84 = ~x10 & x11 ;
  assign n85 = x6 & ~x7 ;
  assign n86 = n84 & ~n85 ;
  assign n87 = ~n83 & n86 ;
  assign n88 = ~x7 & x16 ;
  assign n89 = ~x9 & ~n88 ;
  assign n90 = n87 & ~n89 ;
  assign n91 = n90 ^ n73 ;
  assign n92 = n81 & ~n91 ;
  assign n93 = n92 ^ n74 ;
  assign n94 = n77 & ~n93 ;
  assign n95 = n94 ^ n92 ;
  assign n96 = ~n73 & n95 ;
  assign n97 = n96 ^ n92 ;
  assign n98 = n97 ^ n94 ;
  assign n99 = n98 ^ x2 ;
  assign n100 = ~n72 & ~n99 ;
  assign n101 = ~x3 & ~n100 ;
  assign n102 = ~n45 & ~n101 ;
  assign n103 = ~x1 & x3 ;
  assign n104 = ~x2 & n103 ;
  assign n105 = ~x0 & ~x2 ;
  assign n106 = ~x3 & ~n105 ;
  assign n108 = ~x12 & ~x13 ;
  assign n109 = x9 & n108 ;
  assign n107 = x3 ^ x1 ;
  assign n110 = n109 ^ n107 ;
  assign n111 = n110 ^ x3 ;
  assign n112 = n111 ^ x3 ;
  assign n113 = n112 ^ n107 ;
  assign n139 = n113 ^ n107 ;
  assign n140 = n139 ^ x3 ;
  assign n114 = x10 ^ x9 ;
  assign n115 = ~x6 & ~x7 ;
  assign n116 = ~x11 & n115 ;
  assign n117 = n108 & n116 ;
  assign n118 = n117 ^ x11 ;
  assign n119 = n118 ^ n117 ;
  assign n120 = ~x12 & n115 ;
  assign n121 = ~x13 & ~n120 ;
  assign n122 = n121 ^ n117 ;
  assign n123 = n122 ^ n117 ;
  assign n124 = n119 & ~n123 ;
  assign n125 = n124 ^ n117 ;
  assign n126 = n125 ^ x10 ;
  assign n127 = n114 & ~n126 ;
  assign n128 = n127 ^ n124 ;
  assign n129 = n128 ^ n117 ;
  assign n130 = n129 ^ x9 ;
  assign n131 = ~x10 & ~n130 ;
  assign n132 = n131 ^ x10 ;
  assign n133 = n132 ^ n117 ;
  assign n134 = ~x8 & ~n133 ;
  assign n135 = n134 ^ n107 ;
  assign n136 = n135 ^ n113 ;
  assign n137 = n136 ^ n107 ;
  assign n138 = n137 ^ x3 ;
  assign n141 = n140 ^ n138 ;
  assign n142 = x3 & n141 ;
  assign n143 = n142 ^ n113 ;
  assign n144 = n143 ^ n140 ;
  assign n150 = n107 ^ x2 ;
  assign n145 = x8 & ~x11 ;
  assign n146 = x10 & n145 ;
  assign n147 = n146 ^ x2 ;
  assign n148 = n140 ^ n113 ;
  assign n149 = n147 & n148 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = n151 ^ n147 ;
  assign n153 = n152 ^ x3 ;
  assign n154 = ~n143 & n153 ;
  assign n155 = n154 ^ n113 ;
  assign n156 = n155 ^ x3 ;
  assign n157 = n156 ^ n140 ;
  assign n158 = n144 & n157 ;
  assign n159 = n158 ^ n113 ;
  assign n160 = n159 ^ x3 ;
  assign n161 = n160 ^ n140 ;
  assign n162 = n161 ^ x1 ;
  assign n163 = ~n106 & ~n162 ;
  assign n164 = n163 ^ x4 ;
  assign n165 = n164 ^ n163 ;
  assign n166 = ~x1 & ~x3 ;
  assign n167 = n54 & n61 ;
  assign n168 = n166 & n167 ;
  assign n169 = n168 ^ n163 ;
  assign n170 = n165 & ~n169 ;
  assign n171 = n170 ^ n163 ;
  assign n172 = ~n104 & n171 ;
  assign n173 = n102 & n172 ;
  assign n174 = x5 & ~n173 ;
  assign n175 = n103 & n109 ;
  assign n176 = n175 ^ x2 ;
  assign n177 = x8 & n115 ;
  assign n178 = n84 & n177 ;
  assign n179 = n178 ^ n176 ;
  assign n180 = n179 ^ n175 ;
  assign n181 = n180 ^ n179 ;
  assign n182 = ~x0 & ~x3 ;
  assign n183 = ~x8 & n116 ;
  assign n184 = ~n178 & ~n183 ;
  assign n185 = ~x0 & n109 ;
  assign n186 = ~n184 & n185 ;
  assign n187 = x10 & n183 ;
  assign n188 = n23 & n108 ;
  assign n189 = n187 & n188 ;
  assign n190 = ~n186 & ~n189 ;
  assign n191 = ~n182 & n190 ;
  assign n192 = ~x5 & ~n191 ;
  assign n193 = n192 ^ n179 ;
  assign n194 = n193 ^ n176 ;
  assign n195 = n181 & ~n194 ;
  assign n196 = n195 ^ n192 ;
  assign n197 = ~n146 & ~n183 ;
  assign n198 = ~n192 & n197 ;
  assign n199 = n198 ^ n176 ;
  assign n200 = ~n196 & n199 ;
  assign n201 = n200 ^ n198 ;
  assign n202 = n176 & n201 ;
  assign n203 = n202 ^ n195 ;
  assign n204 = n203 ^ x2 ;
  assign n205 = n204 ^ n192 ;
  assign n206 = ~x4 & n205 ;
  assign n207 = ~n146 & n184 ;
  assign n208 = x9 & ~n207 ;
  assign n209 = ~n187 & ~n208 ;
  assign n210 = n108 & ~n209 ;
  assign n211 = ~x4 & n210 ;
  assign n212 = n43 & n211 ;
  assign n213 = ~x9 & n84 ;
  assign n214 = x2 & ~x8 ;
  assign n215 = n213 & n214 ;
  assign n216 = ~x4 & ~n215 ;
  assign n217 = n166 & ~n216 ;
  assign n218 = ~n212 & ~n217 ;
  assign n219 = x0 & ~n218 ;
  assign n220 = ~n206 & ~n219 ;
  assign n221 = x3 & x4 ;
  assign n222 = ~x5 & n221 ;
  assign n223 = n222 ^ x1 ;
  assign n224 = n222 ^ x0 ;
  assign n225 = n224 ^ x0 ;
  assign n226 = x4 ^ x2 ;
  assign n227 = n226 ^ x2 ;
  assign n228 = n227 ^ x0 ;
  assign n229 = n210 ^ x3 ;
  assign n230 = ~x3 & ~n229 ;
  assign n231 = n230 ^ x2 ;
  assign n232 = n231 ^ x3 ;
  assign n233 = n228 & ~n232 ;
  assign n234 = n233 ^ n230 ;
  assign n235 = n234 ^ x3 ;
  assign n236 = ~x0 & ~n235 ;
  assign n237 = n236 ^ x0 ;
  assign n238 = ~n225 & ~n237 ;
  assign n239 = n238 ^ x0 ;
  assign n240 = n223 & n239 ;
  assign n241 = n240 ^ x1 ;
  assign n242 = n220 & ~n241 ;
  assign n243 = ~n174 & n242 ;
  assign n244 = n243 ^ x19 ;
  assign n245 = n42 & n244 ;
  assign n246 = n245 ^ x19 ;
  assign n247 = x14 & n246 ;
  assign n248 = ~n39 & n247 ;
  assign y0 = ~n248 ;
endmodule
