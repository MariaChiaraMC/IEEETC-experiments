module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 ;
  assign n9 = ~x0 & ~x1 ;
  assign n10 = ~x2 & n9 ;
  assign n14 = ~x6 & ~x7 ;
  assign n15 = x5 & ~n14 ;
  assign n11 = ~x5 & ~x7 ;
  assign n12 = ~x4 & n11 ;
  assign n13 = ~x3 & ~n12 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = ~x3 & x6 ;
  assign n19 = x4 & ~n18 ;
  assign n20 = n19 ^ n13 ;
  assign n21 = n17 & n20 ;
  assign n22 = n21 ^ n13 ;
  assign n23 = n10 & ~n22 ;
  assign y0 = n23 ;
endmodule
