module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 ;
  assign n7 = x1 & x2 ;
  assign n8 = ~x4 & x5 ;
  assign n9 = x0 & n8 ;
  assign n10 = n7 & n9 ;
  assign n11 = x2 ^ x1 ;
  assign n38 = n11 ^ x5 ;
  assign n39 = n11 & n38 ;
  assign n40 = x0 & n39 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = x4 & n41 ;
  assign n43 = x1 & ~x2 ;
  assign n44 = ~x0 & n43 ;
  assign n45 = n8 & n44 ;
  assign n46 = ~n42 & ~n45 ;
  assign n12 = n11 ^ x4 ;
  assign n13 = n12 ^ x5 ;
  assign n14 = n13 ^ x0 ;
  assign n15 = n14 ^ x2 ;
  assign n16 = n15 ^ x5 ;
  assign n17 = n16 ^ x2 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = n16 ^ x4 ;
  assign n20 = n19 ^ x5 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = n21 ^ n13 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n23 ^ n16 ;
  assign n25 = ~x2 & n24 ;
  assign n26 = n25 ^ n13 ;
  assign n27 = n26 ^ n18 ;
  assign n28 = n22 ^ x2 ;
  assign n29 = n28 ^ n18 ;
  assign n30 = n13 & n29 ;
  assign n31 = n30 ^ x2 ;
  assign n32 = n27 & ~n31 ;
  assign n33 = n18 & n32 ;
  assign n34 = n33 ^ n25 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ n13 ;
  assign n47 = n46 ^ n37 ;
  assign n48 = ~x3 & ~n47 ;
  assign n49 = n48 ^ n37 ;
  assign n50 = ~n10 & ~n49 ;
  assign y0 = ~n50 ;
endmodule
