module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n9 = ~x0 & x1 ;
  assign n10 = ~x7 & n9 ;
  assign n11 = ~x2 & ~x3 ;
  assign n12 = ~n10 & n11 ;
  assign n17 = ~x4 & ~x6 ;
  assign n13 = x6 & x7 ;
  assign n18 = n17 ^ n13 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = n15 ^ x2 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n20 ^ x3 ;
  assign n22 = n21 ^ n20 ;
  assign n25 = n17 ^ n15 ;
  assign n26 = n25 ^ n18 ;
  assign n27 = n26 ^ n20 ;
  assign n28 = ~n20 & n27 ;
  assign n23 = n15 & ~n18 ;
  assign n31 = n28 ^ n23 ;
  assign n24 = n23 ^ n22 ;
  assign n29 = n28 ^ n20 ;
  assign n30 = ~n24 & ~n29 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = ~n22 & n32 ;
  assign n34 = n33 ^ n28 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n35 ^ n14 ;
  assign n37 = ~n12 & n36 ;
  assign y0 = n37 ;
endmodule
