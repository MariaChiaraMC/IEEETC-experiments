module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 ;
  assign n17 = x2 & ~x14 ;
  assign n18 = ~x8 & n17 ;
  assign n19 = x3 & n18 ;
  assign n20 = x4 & x15 ;
  assign n21 = x1 & n20 ;
  assign n22 = n19 & n21 ;
  assign n23 = x5 & x7 ;
  assign n24 = x10 ^ x7 ;
  assign n25 = ~n23 & n24 ;
  assign n26 = x6 & n25 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = n22 & ~n27 ;
  assign n29 = x8 & x10 ;
  assign n30 = ~x2 & n29 ;
  assign n31 = ~x4 & n30 ;
  assign n32 = x3 & ~x6 ;
  assign n33 = ~x14 & n32 ;
  assign n34 = n23 & n33 ;
  assign n35 = n31 & n34 ;
  assign n36 = ~x3 & ~x7 ;
  assign n39 = ~x4 & ~x5 ;
  assign n40 = x6 & n39 ;
  assign n37 = x6 & x10 ;
  assign n38 = n18 & ~n37 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = x4 & x5 ;
  assign n43 = x10 & n42 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = n44 ^ n43 ;
  assign n46 = n45 ^ n41 ;
  assign n47 = x11 & x14 ;
  assign n48 = n47 ^ n30 ;
  assign n49 = n30 & n48 ;
  assign n50 = n49 ^ n43 ;
  assign n51 = n50 ^ n30 ;
  assign n52 = ~n46 & ~n51 ;
  assign n53 = n52 ^ n49 ;
  assign n54 = n53 ^ n30 ;
  assign n55 = n41 & n54 ;
  assign n56 = n55 ^ n38 ;
  assign n57 = n36 & n56 ;
  assign n58 = ~n35 & ~n57 ;
  assign n59 = ~x1 & ~x15 ;
  assign n60 = ~n58 & n59 ;
  assign n61 = ~n28 & ~n60 ;
  assign n62 = x9 & ~n61 ;
  assign n63 = ~x1 & x10 ;
  assign n64 = ~x6 & n63 ;
  assign n65 = x15 ^ x7 ;
  assign n66 = n39 ^ x15 ;
  assign n67 = n66 ^ n39 ;
  assign n68 = ~x9 & n42 ;
  assign n69 = n68 ^ n39 ;
  assign n70 = ~n67 & n69 ;
  assign n71 = n70 ^ n39 ;
  assign n72 = ~n65 & n71 ;
  assign n73 = n64 & n72 ;
  assign n74 = n19 & n73 ;
  assign n75 = ~n62 & ~n74 ;
  assign n76 = ~x12 & ~x13 ;
  assign n77 = ~x0 & n76 ;
  assign n78 = ~n75 & n77 ;
  assign y0 = n78 ;
endmodule
