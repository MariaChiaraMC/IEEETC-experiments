module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ;
  assign n13 = x8 ^ x4 ;
  assign n23 = n13 ^ x1 ;
  assign n14 = n13 ^ x2 ;
  assign n15 = n14 ^ n13 ;
  assign n24 = n15 ^ x6 ;
  assign n25 = n23 & n24 ;
  assign n16 = x8 ^ x7 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n16 ^ x8 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = n17 & ~n19 ;
  assign n31 = n25 ^ n20 ;
  assign n21 = n20 ^ n15 ;
  assign n22 = n21 ^ n17 ;
  assign n26 = n16 ^ n13 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = n27 ^ n23 ;
  assign n29 = n28 ^ x6 ;
  assign n30 = n22 & ~n29 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = n32 ^ n26 ;
  assign n34 = n33 ^ n23 ;
  assign n35 = n34 ^ x6 ;
  assign n36 = x6 & ~n35 ;
  assign n37 = n36 ^ x6 ;
  assign n38 = n37 ^ x8 ;
  assign n39 = n38 ^ x6 ;
  assign y0 = n39 ;
endmodule
