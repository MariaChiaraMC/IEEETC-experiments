module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n15 = ~x2 & ~x3 ;
  assign n16 = ~x0 & x4 ;
  assign n17 = ~x1 & x5 ;
  assign n18 = n16 & n17 ;
  assign n19 = n15 & n18 ;
  assign n20 = x7 ^ x6 ;
  assign n21 = n20 ^ x7 ;
  assign n22 = ~x11 & ~x13 ;
  assign n23 = ~x10 & n22 ;
  assign n24 = ~x7 & x12 ;
  assign n25 = x9 ^ x8 ;
  assign n26 = n24 & n25 ;
  assign n27 = n23 & n26 ;
  assign n28 = n27 ^ x7 ;
  assign n29 = ~n21 & n28 ;
  assign n30 = n29 ^ x7 ;
  assign n31 = n19 & n30 ;
  assign y0 = n31 ;
endmodule
