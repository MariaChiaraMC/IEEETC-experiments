module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 ;
  assign n9 = x4 & x5 ;
  assign n10 = x6 & x7 ;
  assign n11 = n9 & n10 ;
  assign n12 = x0 & ~x1 ;
  assign n13 = ~n11 & n12 ;
  assign n14 = ~x2 & n13 ;
  assign n32 = ~x6 & ~x7 ;
  assign n46 = x0 & x2 ;
  assign n47 = ~n32 & ~n46 ;
  assign n48 = ~x1 & ~n47 ;
  assign n49 = x4 & ~n48 ;
  assign n50 = x1 & x2 ;
  assign n51 = ~x5 & ~n10 ;
  assign n52 = n50 & ~n51 ;
  assign n53 = ~x0 & ~x2 ;
  assign n54 = ~n9 & n53 ;
  assign n55 = ~n46 & ~n54 ;
  assign n56 = ~n52 & ~n55 ;
  assign n57 = ~n49 & n56 ;
  assign n15 = x1 ^ x0 ;
  assign n16 = n15 ^ x4 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n18 ^ x1 ;
  assign n20 = ~n18 & n19 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = n15 ^ x2 ;
  assign n24 = n23 ^ x5 ;
  assign n30 = n24 ^ x5 ;
  assign n25 = n24 ^ n15 ;
  assign n26 = n25 ^ n17 ;
  assign n27 = n26 ^ n18 ;
  assign n28 = ~n17 & n27 ;
  assign n29 = n28 ^ n25 ;
  assign n31 = n30 ^ n29 ;
  assign n33 = n32 ^ n25 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = ~n32 & ~n34 ;
  assign n36 = n35 ^ n17 ;
  assign n37 = n31 & ~n36 ;
  assign n38 = n37 ^ n25 ;
  assign n39 = n38 ^ n18 ;
  assign n40 = n39 ^ x1 ;
  assign n41 = n22 & n40 ;
  assign n42 = n41 ^ n28 ;
  assign n43 = n42 ^ n37 ;
  assign n44 = n43 ^ n17 ;
  assign n45 = n44 ^ n15 ;
  assign n58 = n57 ^ n45 ;
  assign n59 = n58 ^ n57 ;
  assign n60 = ~x4 & ~x5 ;
  assign n61 = n32 ^ x1 ;
  assign n62 = ~x2 & n61 ;
  assign n63 = n62 ^ x1 ;
  assign n64 = n60 & n63 ;
  assign n65 = n64 ^ n57 ;
  assign n66 = n65 ^ n57 ;
  assign n67 = n59 & ~n66 ;
  assign n68 = n67 ^ n57 ;
  assign n69 = x3 & n68 ;
  assign n70 = n69 ^ n57 ;
  assign n71 = ~n14 & n70 ;
  assign y0 = ~n71 ;
endmodule
