module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 ;
  assign n7 = x1 ^ x0 ;
  assign n8 = n7 ^ x2 ;
  assign n10 = n8 ^ x2 ;
  assign n9 = n8 ^ x1 ;
  assign n11 = n10 ^ n9 ;
  assign n16 = n11 ^ n8 ;
  assign n17 = n16 ^ n10 ;
  assign n18 = n17 ^ n10 ;
  assign n19 = x4 & x5 ;
  assign n20 = n19 ^ n8 ;
  assign n21 = n20 ^ n8 ;
  assign n22 = n21 ^ n10 ;
  assign n23 = n18 & ~n22 ;
  assign n12 = n8 ^ x3 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n13 ^ n10 ;
  assign n15 = n11 & n14 ;
  assign n24 = n23 ^ n15 ;
  assign n25 = n24 ^ n11 ;
  assign n26 = n15 ^ n10 ;
  assign n27 = n26 ^ n17 ;
  assign n28 = n10 & n27 ;
  assign n29 = n28 ^ n15 ;
  assign n30 = n25 & n29 ;
  assign n31 = n30 ^ n23 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = n32 ^ n11 ;
  assign n34 = n33 ^ n10 ;
  assign n35 = n34 ^ n17 ;
  assign n36 = n35 ^ x2 ;
  assign y0 = n36 ;
endmodule
