module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 ;
  assign n15 = x7 & ~x8 ;
  assign n16 = x6 & n15 ;
  assign n17 = ~x10 & ~n16 ;
  assign n18 = ~x4 & ~x10 ;
  assign n19 = x13 & ~n18 ;
  assign n20 = n19 ^ x12 ;
  assign n21 = n20 ^ x11 ;
  assign n30 = n21 ^ n20 ;
  assign n22 = ~x3 & ~x9 ;
  assign n23 = x2 & ~n22 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n24 ^ n20 ;
  assign n26 = n21 ^ n19 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n25 & ~n28 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n31 ^ n25 ;
  assign n33 = n20 ^ x0 ;
  assign n34 = n29 ^ n25 ;
  assign n35 = n33 & n34 ;
  assign n36 = n35 ^ n20 ;
  assign n37 = n32 & n36 ;
  assign n38 = n37 ^ n20 ;
  assign n39 = n38 ^ x12 ;
  assign n40 = n39 ^ n20 ;
  assign n41 = ~n17 & n40 ;
  assign n42 = x7 ^ x6 ;
  assign n43 = n42 ^ n15 ;
  assign n44 = ~x5 & ~n43 ;
  assign n45 = n44 ^ n15 ;
  assign n46 = ~x4 & n45 ;
  assign n47 = n16 ^ x10 ;
  assign n48 = x11 ^ x10 ;
  assign n49 = n48 ^ x10 ;
  assign n50 = n47 & n49 ;
  assign n51 = n50 ^ x10 ;
  assign n52 = ~x1 & n51 ;
  assign n53 = ~n46 & ~n52 ;
  assign n54 = x12 & ~n53 ;
  assign n55 = ~n41 & ~n54 ;
  assign y0 = ~n55 ;
endmodule
