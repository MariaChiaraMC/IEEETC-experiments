module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 ;
  assign n11 = x3 & x5 ;
  assign n24 = ~x7 & x8 ;
  assign n12 = ~x0 & ~x8 ;
  assign n13 = ~x1 & n12 ;
  assign n15 = x4 & ~x7 ;
  assign n14 = ~x4 & x7 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = x2 & n16 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n13 & n18 ;
  assign n25 = n24 ^ n19 ;
  assign n26 = n25 ^ n19 ;
  assign n20 = x0 & ~x2 ;
  assign n21 = x1 & n20 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ n19 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = n19 ^ x4 ;
  assign n29 = n28 ^ n19 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n26 & ~n30 ;
  assign n32 = n31 ^ n26 ;
  assign n33 = n27 & n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n34 ^ n19 ;
  assign n36 = n35 ^ n26 ;
  assign n37 = ~x6 & n36 ;
  assign n38 = n37 ^ n19 ;
  assign n39 = n11 & n38 ;
  assign n40 = x0 & x1 ;
  assign n41 = x7 & ~x8 ;
  assign n42 = n40 & n41 ;
  assign n43 = ~x4 & x5 ;
  assign n44 = ~x2 & ~x3 ;
  assign n45 = n43 & n44 ;
  assign n46 = n42 & n45 ;
  assign n47 = x2 & ~x3 ;
  assign n48 = ~x0 & n47 ;
  assign n49 = x5 & ~x7 ;
  assign n50 = n48 & n49 ;
  assign n51 = x3 & ~x5 ;
  assign n52 = ~x2 & ~x7 ;
  assign n53 = n51 & n52 ;
  assign n54 = ~n20 & ~n53 ;
  assign n55 = x5 ^ x3 ;
  assign n56 = x7 ^ x5 ;
  assign n57 = ~n55 & n56 ;
  assign n58 = x0 & n57 ;
  assign n59 = n58 ^ x0 ;
  assign n60 = ~n54 & ~n59 ;
  assign n61 = ~n50 & ~n60 ;
  assign n64 = n61 ^ x3 ;
  assign n65 = n64 ^ n61 ;
  assign n62 = n61 ^ n20 ;
  assign n63 = n62 ^ n61 ;
  assign n66 = n65 ^ n63 ;
  assign n67 = x5 & x7 ;
  assign n68 = n67 ^ n61 ;
  assign n69 = n68 ^ n61 ;
  assign n70 = n69 ^ n65 ;
  assign n71 = n65 & n70 ;
  assign n72 = n71 ^ n65 ;
  assign n73 = n66 & n72 ;
  assign n74 = n73 ^ n71 ;
  assign n75 = n74 ^ n61 ;
  assign n76 = n75 ^ n65 ;
  assign n77 = x1 & ~n76 ;
  assign n78 = n77 ^ n61 ;
  assign n79 = x8 & ~n78 ;
  assign n80 = n40 & n53 ;
  assign n81 = ~n79 & ~n80 ;
  assign n82 = x4 & ~n81 ;
  assign n85 = ~x1 & x3 ;
  assign n83 = ~x1 & ~n43 ;
  assign n84 = x7 & ~n83 ;
  assign n86 = n85 ^ n84 ;
  assign n87 = x5 ^ x4 ;
  assign n88 = x2 & x3 ;
  assign n89 = n88 ^ x5 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = n88 ^ n44 ;
  assign n92 = n90 & n91 ;
  assign n93 = n92 ^ n88 ;
  assign n94 = ~n87 & n93 ;
  assign n95 = n94 ^ n84 ;
  assign n96 = n95 ^ n94 ;
  assign n97 = n96 ^ n86 ;
  assign n98 = ~x5 & ~n15 ;
  assign n99 = x4 & x5 ;
  assign n100 = x2 & ~n99 ;
  assign n101 = n100 ^ n98 ;
  assign n102 = ~n98 & ~n101 ;
  assign n103 = n102 ^ n94 ;
  assign n104 = n103 ^ n98 ;
  assign n105 = ~n97 & n104 ;
  assign n106 = n105 ^ n102 ;
  assign n107 = n106 ^ n98 ;
  assign n108 = n86 & ~n107 ;
  assign n109 = n108 ^ n84 ;
  assign n110 = n12 & n109 ;
  assign n123 = ~x1 & ~x5 ;
  assign n124 = x0 & ~x4 ;
  assign n125 = n123 & n124 ;
  assign n111 = n47 & n49 ;
  assign n112 = x1 & n111 ;
  assign n113 = n21 & n51 ;
  assign n114 = ~x3 & x5 ;
  assign n115 = x0 & n114 ;
  assign n116 = x7 ^ x2 ;
  assign n117 = n115 & n116 ;
  assign n118 = ~n113 & ~n117 ;
  assign n119 = ~n112 & n118 ;
  assign n120 = ~x4 & ~n119 ;
  assign n126 = n125 ^ n120 ;
  assign n127 = n126 ^ n120 ;
  assign n121 = n120 ^ n44 ;
  assign n122 = n121 ^ n120 ;
  assign n128 = n127 ^ n122 ;
  assign n129 = n120 ^ x7 ;
  assign n130 = n129 ^ n120 ;
  assign n131 = n130 ^ n127 ;
  assign n132 = n127 & ~n131 ;
  assign n133 = n132 ^ n127 ;
  assign n134 = n128 & n133 ;
  assign n135 = n134 ^ n132 ;
  assign n136 = n135 ^ n120 ;
  assign n137 = n136 ^ n127 ;
  assign n138 = x8 & n137 ;
  assign n139 = n138 ^ n120 ;
  assign n140 = ~n110 & ~n139 ;
  assign n141 = ~n82 & n140 ;
  assign n142 = n141 ^ x6 ;
  assign n143 = n142 ^ n141 ;
  assign n158 = n24 & n123 ;
  assign n159 = n11 & n41 ;
  assign n160 = ~n158 & ~n159 ;
  assign n161 = x0 & ~n160 ;
  assign n162 = ~x0 & x5 ;
  assign n163 = n24 ^ x3 ;
  assign n164 = n163 ^ x1 ;
  assign n165 = n164 ^ n24 ;
  assign n166 = n165 ^ n162 ;
  assign n167 = x8 ^ x1 ;
  assign n168 = ~x8 & ~n167 ;
  assign n169 = n168 ^ n24 ;
  assign n170 = n169 ^ x8 ;
  assign n171 = ~n166 & ~n170 ;
  assign n172 = n171 ^ n168 ;
  assign n173 = n172 ^ x8 ;
  assign n174 = n162 & ~n173 ;
  assign n175 = ~n161 & ~n174 ;
  assign n144 = x8 ^ x7 ;
  assign n145 = n144 ^ n56 ;
  assign n146 = x1 ^ x0 ;
  assign n147 = n146 ^ x0 ;
  assign n148 = x8 ^ x0 ;
  assign n149 = ~n147 & ~n148 ;
  assign n150 = n149 ^ x0 ;
  assign n151 = n150 ^ n144 ;
  assign n152 = n145 & n151 ;
  assign n153 = n152 ^ n149 ;
  assign n154 = n153 ^ x0 ;
  assign n155 = n154 ^ n56 ;
  assign n156 = ~n144 & n155 ;
  assign n157 = n156 ^ n144 ;
  assign n176 = n175 ^ n157 ;
  assign n177 = n176 ^ n175 ;
  assign n178 = n175 ^ x3 ;
  assign n179 = n178 ^ n175 ;
  assign n180 = ~n177 & ~n179 ;
  assign n181 = n180 ^ n175 ;
  assign n182 = ~x4 & ~n181 ;
  assign n183 = n182 ^ n175 ;
  assign n184 = ~x2 & ~n183 ;
  assign n188 = x7 & x8 ;
  assign n189 = x5 & n188 ;
  assign n190 = x3 & n189 ;
  assign n185 = ~x3 & x7 ;
  assign n186 = ~x8 & n11 ;
  assign n187 = ~n185 & ~n186 ;
  assign n191 = n190 ^ n187 ;
  assign n192 = n191 ^ n190 ;
  assign n193 = n190 ^ n41 ;
  assign n194 = n193 ^ n190 ;
  assign n195 = ~n192 & ~n194 ;
  assign n196 = n195 ^ n190 ;
  assign n197 = x1 & n196 ;
  assign n198 = n197 ^ n190 ;
  assign n199 = x0 & n198 ;
  assign n200 = ~x7 & ~x8 ;
  assign n201 = n114 & n200 ;
  assign n202 = ~x1 & n201 ;
  assign n203 = ~n199 & ~n202 ;
  assign n204 = x4 & ~n20 ;
  assign n205 = ~n203 & n204 ;
  assign n206 = ~n184 & ~n205 ;
  assign n207 = n206 ^ n141 ;
  assign n208 = ~n143 & n207 ;
  assign n209 = n208 ^ n141 ;
  assign n210 = ~n46 & n209 ;
  assign n211 = n210 ^ x9 ;
  assign n212 = n211 ^ n210 ;
  assign n213 = n44 & n188 ;
  assign n214 = x5 & ~x6 ;
  assign n215 = n124 & n214 ;
  assign n216 = n213 & n215 ;
  assign n217 = ~x3 & ~x5 ;
  assign n218 = n41 & n217 ;
  assign n219 = ~x4 & ~x6 ;
  assign n220 = n218 & n219 ;
  assign n221 = ~x2 & n220 ;
  assign n222 = ~n99 & n185 ;
  assign n223 = ~x5 & ~x7 ;
  assign n224 = x3 & x4 ;
  assign n225 = n223 & n224 ;
  assign n226 = ~x6 & n225 ;
  assign n227 = ~n222 & ~n226 ;
  assign n228 = ~x8 & ~n227 ;
  assign n229 = ~x6 & n99 ;
  assign n230 = n24 & n229 ;
  assign n231 = ~n228 & ~n230 ;
  assign n232 = n20 & ~n231 ;
  assign n233 = x2 & n124 ;
  assign n234 = ~n114 & n233 ;
  assign n235 = n214 ^ n24 ;
  assign n236 = n235 ^ n234 ;
  assign n237 = n41 ^ x3 ;
  assign n238 = n24 & n237 ;
  assign n239 = n238 ^ n41 ;
  assign n240 = n236 & n239 ;
  assign n241 = n240 ^ n238 ;
  assign n242 = n241 ^ n41 ;
  assign n243 = n242 ^ n24 ;
  assign n244 = n234 & n243 ;
  assign n245 = ~n232 & ~n244 ;
  assign n246 = x3 & ~x4 ;
  assign n247 = n41 & n246 ;
  assign n248 = n247 ^ x4 ;
  assign n249 = n248 ^ n247 ;
  assign n250 = ~x3 & n24 ;
  assign n251 = n250 ^ n247 ;
  assign n252 = n251 ^ n247 ;
  assign n253 = n249 & n252 ;
  assign n254 = n253 ^ n247 ;
  assign n255 = x5 & n254 ;
  assign n256 = n255 ^ n247 ;
  assign n257 = x2 & n256 ;
  assign n258 = n67 & ~n88 ;
  assign n259 = n224 ^ x4 ;
  assign n260 = x8 & ~n259 ;
  assign n261 = n260 ^ x4 ;
  assign n262 = n258 & ~n261 ;
  assign n263 = ~n257 & ~n262 ;
  assign n264 = n263 ^ x0 ;
  assign n265 = n264 ^ n263 ;
  assign n266 = n265 ^ x6 ;
  assign n267 = ~x7 & n11 ;
  assign n268 = n267 ^ x2 ;
  assign n269 = n268 ^ n267 ;
  assign n270 = n269 ^ x4 ;
  assign n271 = n218 ^ n190 ;
  assign n272 = ~n190 & n271 ;
  assign n273 = n272 ^ n267 ;
  assign n274 = n273 ^ n190 ;
  assign n275 = n270 & n274 ;
  assign n276 = n275 ^ n272 ;
  assign n277 = n276 ^ n190 ;
  assign n278 = x4 & ~n277 ;
  assign n279 = n278 ^ x4 ;
  assign n280 = ~x3 & ~x4 ;
  assign n281 = ~x5 & x8 ;
  assign n282 = n280 & n281 ;
  assign n283 = ~n186 & ~n282 ;
  assign n284 = n52 & ~n283 ;
  assign n285 = n284 ^ n279 ;
  assign n286 = ~n279 & n285 ;
  assign n287 = n286 ^ n263 ;
  assign n288 = n287 ^ n279 ;
  assign n289 = ~n266 & ~n288 ;
  assign n290 = n289 ^ n286 ;
  assign n291 = n290 ^ n279 ;
  assign n292 = x6 & ~n291 ;
  assign n293 = n292 ^ x6 ;
  assign n294 = n245 & ~n293 ;
  assign n295 = ~n221 & n294 ;
  assign n296 = n295 ^ x1 ;
  assign n297 = n296 ^ n295 ;
  assign n298 = n24 & n48 ;
  assign n299 = n43 & n298 ;
  assign n300 = n246 & n281 ;
  assign n301 = x4 & ~x8 ;
  assign n302 = n114 & n301 ;
  assign n303 = ~n300 & ~n302 ;
  assign n304 = ~x7 & n20 ;
  assign n305 = ~n303 & n304 ;
  assign n306 = n189 & n280 ;
  assign n307 = x3 & n301 ;
  assign n308 = ~n223 & n307 ;
  assign n309 = ~n306 & ~n308 ;
  assign n310 = n309 ^ x0 ;
  assign n311 = n310 ^ n309 ;
  assign n312 = n15 ^ x3 ;
  assign n313 = n312 ^ n15 ;
  assign n314 = n16 & n313 ;
  assign n315 = n314 ^ n15 ;
  assign n316 = ~x5 & n315 ;
  assign n317 = x8 & n316 ;
  assign n318 = n317 ^ n309 ;
  assign n319 = ~n311 & ~n318 ;
  assign n320 = n319 ^ n309 ;
  assign n321 = x2 & ~n320 ;
  assign n322 = ~n305 & ~n321 ;
  assign n323 = n322 ^ x6 ;
  assign n324 = n323 ^ n322 ;
  assign n325 = n124 ^ x7 ;
  assign n326 = x2 & n325 ;
  assign n327 = n326 ^ x7 ;
  assign n328 = ~n14 & n327 ;
  assign n329 = n281 & n328 ;
  assign n330 = ~x0 & ~x5 ;
  assign n331 = ~x4 & n88 ;
  assign n332 = n200 & n331 ;
  assign n333 = ~n213 & ~n332 ;
  assign n334 = n330 & ~n333 ;
  assign n335 = ~n15 & ~n185 ;
  assign n336 = n162 & ~n246 ;
  assign n337 = ~n301 & n336 ;
  assign n338 = n335 & n337 ;
  assign n339 = x2 & n338 ;
  assign n340 = ~n334 & ~n339 ;
  assign n341 = ~n329 & n340 ;
  assign n342 = n341 ^ n322 ;
  assign n343 = ~n324 & n342 ;
  assign n344 = n343 ^ n322 ;
  assign n345 = ~n299 & n344 ;
  assign n346 = n345 ^ n295 ;
  assign n347 = n297 & n346 ;
  assign n348 = n347 ^ n295 ;
  assign n349 = ~n216 & n348 ;
  assign n350 = n349 ^ n210 ;
  assign n351 = ~n212 & n350 ;
  assign n352 = n351 ^ n210 ;
  assign n353 = ~n39 & n352 ;
  assign y0 = ~n353 ;
endmodule
