module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 ;
  assign n9 = x1 & ~x2 ;
  assign n10 = x6 & n9 ;
  assign n11 = x2 & x5 ;
  assign n12 = n11 ^ x0 ;
  assign n13 = x7 ^ x0 ;
  assign n14 = n13 ^ x0 ;
  assign n15 = n12 & n14 ;
  assign n16 = n15 ^ x0 ;
  assign n17 = ~n10 & ~n16 ;
  assign n18 = n17 ^ x0 ;
  assign n19 = x1 & x6 ;
  assign n20 = n19 ^ n11 ;
  assign n21 = ~x7 & n20 ;
  assign n22 = n18 & ~n21 ;
  assign n23 = ~x3 & ~n22 ;
  assign n24 = x6 ^ x5 ;
  assign n25 = ~x1 & x2 ;
  assign n26 = n25 ^ x6 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = n25 ^ n9 ;
  assign n29 = n27 & n28 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = n24 & n30 ;
  assign n32 = ~x0 & n31 ;
  assign n33 = x3 & ~x7 ;
  assign n34 = n19 & n33 ;
  assign n35 = ~n32 & ~n34 ;
  assign n45 = ~x1 & ~x2 ;
  assign n46 = ~x5 & ~x6 ;
  assign n47 = ~n45 & ~n46 ;
  assign n48 = x1 & x2 ;
  assign n49 = x5 & x6 ;
  assign n50 = ~n48 & ~n49 ;
  assign n51 = x3 & ~n50 ;
  assign n52 = n47 & ~n51 ;
  assign n36 = x2 ^ x1 ;
  assign n37 = ~x5 & x6 ;
  assign n38 = n37 ^ x2 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = x5 & ~x6 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = ~n39 & n41 ;
  assign n43 = n42 ^ n37 ;
  assign n44 = n36 & n43 ;
  assign n53 = n52 ^ n44 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = n52 ^ x3 ;
  assign n56 = n55 ^ n52 ;
  assign n57 = n54 & n56 ;
  assign n58 = n57 ^ n52 ;
  assign n59 = ~x0 & ~n58 ;
  assign n60 = n59 ^ n52 ;
  assign n61 = n60 ^ x7 ;
  assign n62 = n61 ^ n60 ;
  assign n63 = x2 & n40 ;
  assign n64 = n63 ^ n60 ;
  assign n65 = ~n62 & ~n64 ;
  assign n66 = n65 ^ n60 ;
  assign n67 = n35 & n66 ;
  assign n68 = n67 ^ x4 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = ~x0 & x3 ;
  assign n71 = ~n47 & n70 ;
  assign n72 = n33 & ~n63 ;
  assign n73 = ~n19 & n72 ;
  assign n74 = ~x0 & ~n51 ;
  assign n75 = x3 & n31 ;
  assign n76 = ~n44 & ~n70 ;
  assign n77 = ~n75 & n76 ;
  assign n78 = x7 & ~n77 ;
  assign n79 = ~n74 & n78 ;
  assign n80 = ~n73 & ~n79 ;
  assign n81 = ~n71 & n80 ;
  assign n82 = n81 ^ n67 ;
  assign n83 = n69 & n82 ;
  assign n84 = n83 ^ n67 ;
  assign n85 = ~n23 & n84 ;
  assign y0 = ~n85 ;
endmodule
