module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 ;
  output y0 ;
  wire n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 ;
  assign n19 = ~x15 & ~x16 ;
  assign n20 = ~x0 & n19 ;
  assign n21 = ~x6 & ~x7 ;
  assign n22 = ~x8 & n21 ;
  assign n23 = ~x14 & x17 ;
  assign n24 = ~n22 & n23 ;
  assign n25 = n24 ^ x13 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n26 ^ n20 ;
  assign n28 = x8 & x9 ;
  assign n29 = n21 & ~n28 ;
  assign n30 = ~x10 & n29 ;
  assign n31 = ~x2 & x14 ;
  assign n32 = n30 & n31 ;
  assign n33 = x17 & ~n32 ;
  assign n34 = x4 & n29 ;
  assign n35 = ~x14 & ~n34 ;
  assign n36 = ~x3 & n35 ;
  assign n37 = n33 & ~n36 ;
  assign n38 = x3 & ~x5 ;
  assign n39 = ~x10 & n38 ;
  assign n40 = x1 & ~x14 ;
  assign n41 = ~x12 & ~x17 ;
  assign n42 = ~x11 & n41 ;
  assign n43 = n40 & n42 ;
  assign n44 = ~n39 & n43 ;
  assign n45 = n44 ^ n37 ;
  assign n46 = ~n37 & n45 ;
  assign n47 = n46 ^ n24 ;
  assign n48 = n47 ^ n37 ;
  assign n49 = ~n27 & n48 ;
  assign n50 = n49 ^ n46 ;
  assign n51 = n50 ^ n37 ;
  assign n52 = n20 & ~n51 ;
  assign n53 = n52 ^ n20 ;
  assign y0 = n53 ;
endmodule
