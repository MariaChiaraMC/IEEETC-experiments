module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 ;
  assign n9 = ~x4 & ~x7 ;
  assign n10 = x3 ^ x1 ;
  assign n11 = n10 ^ x5 ;
  assign n12 = x3 ^ x2 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = x6 ^ x3 ;
  assign n15 = n14 ^ x6 ;
  assign n16 = x6 ^ x5 ;
  assign n17 = n16 ^ x6 ;
  assign n18 = n15 & n17 ;
  assign n19 = n18 ^ x6 ;
  assign n20 = n19 ^ n11 ;
  assign n21 = n13 & ~n20 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = n22 ^ x6 ;
  assign n24 = n23 ^ n12 ;
  assign n25 = ~n11 & ~n24 ;
  assign n26 = n25 ^ n11 ;
  assign n27 = n9 & ~n26 ;
  assign n28 = x5 & x7 ;
  assign n29 = ~x1 & x3 ;
  assign n30 = ~x3 & x4 ;
  assign n31 = ~x6 & n30 ;
  assign n32 = ~n29 & ~n31 ;
  assign n33 = n28 & ~n32 ;
  assign n36 = x7 ^ x1 ;
  assign n34 = x6 ^ x1 ;
  assign n37 = n36 ^ n34 ;
  assign n35 = n34 ^ n10 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = n38 ^ x4 ;
  assign n40 = n39 ^ x1 ;
  assign n41 = n40 ^ x1 ;
  assign n42 = n41 ^ n37 ;
  assign n43 = x5 ^ x1 ;
  assign n44 = n43 ^ x7 ;
  assign n45 = ~n34 & ~n44 ;
  assign n46 = n45 ^ n40 ;
  assign n47 = ~n42 & ~n46 ;
  assign n48 = n47 ^ n37 ;
  assign n49 = n48 ^ n42 ;
  assign n50 = x4 ^ x1 ;
  assign n51 = n50 ^ n37 ;
  assign n52 = n46 ^ n37 ;
  assign n53 = n52 ^ n42 ;
  assign n54 = ~n51 & ~n53 ;
  assign n55 = n54 ^ n40 ;
  assign n56 = n55 ^ n37 ;
  assign n57 = n56 ^ n42 ;
  assign n58 = n49 & ~n57 ;
  assign n59 = n58 ^ n54 ;
  assign n60 = n59 ^ n40 ;
  assign n61 = n60 ^ n37 ;
  assign n62 = n61 ^ n42 ;
  assign n63 = ~n33 & n62 ;
  assign n64 = ~x2 & ~n63 ;
  assign n68 = ~x5 & ~x7 ;
  assign n69 = ~n28 & ~n68 ;
  assign n70 = ~x6 & n69 ;
  assign n71 = x2 & ~x3 ;
  assign n72 = ~x2 & ~x5 ;
  assign n73 = x3 & n72 ;
  assign n74 = ~n71 & ~n73 ;
  assign n75 = n70 & ~n74 ;
  assign n76 = x6 & ~x7 ;
  assign n77 = x3 & x5 ;
  assign n78 = ~x2 & n77 ;
  assign n79 = n76 & n78 ;
  assign n80 = ~n75 & ~n79 ;
  assign n81 = x4 & ~n80 ;
  assign n82 = ~x4 & ~x5 ;
  assign n83 = x7 ^ x3 ;
  assign n84 = n83 ^ x7 ;
  assign n85 = x7 ^ x6 ;
  assign n86 = n85 ^ x7 ;
  assign n87 = ~n84 & ~n86 ;
  assign n88 = n87 ^ x7 ;
  assign n89 = n82 & n88 ;
  assign n90 = x2 & n89 ;
  assign n91 = ~n81 & ~n90 ;
  assign n65 = x6 & x7 ;
  assign n66 = x5 & n65 ;
  assign n67 = n30 & n66 ;
  assign n92 = n91 ^ n67 ;
  assign n93 = ~x1 & ~n92 ;
  assign n94 = n93 ^ n91 ;
  assign n95 = ~n64 & n94 ;
  assign n96 = n95 ^ x0 ;
  assign n97 = n96 ^ n95 ;
  assign n98 = x5 & ~x6 ;
  assign n99 = x4 & n98 ;
  assign n100 = ~n82 & ~n99 ;
  assign n101 = ~x1 & ~x3 ;
  assign n102 = x7 & n101 ;
  assign n103 = ~n100 & n102 ;
  assign n104 = x3 & ~x7 ;
  assign n105 = n99 & n104 ;
  assign n106 = ~x6 & ~x7 ;
  assign n107 = ~n77 & ~n106 ;
  assign n108 = x3 & ~x6 ;
  assign n109 = ~x1 & x4 ;
  assign n110 = ~n108 & n109 ;
  assign n111 = ~n107 & n110 ;
  assign n112 = ~x3 & ~x5 ;
  assign n113 = ~x4 & n65 ;
  assign n114 = n112 & n113 ;
  assign n115 = ~n111 & ~n114 ;
  assign n116 = ~n105 & n115 ;
  assign n117 = n116 ^ x2 ;
  assign n118 = n117 ^ n116 ;
  assign n119 = n118 ^ n103 ;
  assign n128 = x4 & ~x5 ;
  assign n129 = ~n68 & ~n128 ;
  assign n130 = ~n76 & ~n129 ;
  assign n120 = n98 ^ x5 ;
  assign n121 = n120 ^ n98 ;
  assign n122 = n98 ^ n76 ;
  assign n123 = n122 ^ n98 ;
  assign n124 = ~n121 & n123 ;
  assign n125 = n124 ^ n98 ;
  assign n126 = x4 & n125 ;
  assign n127 = n126 ^ n98 ;
  assign n131 = n130 ^ n127 ;
  assign n132 = n131 ^ n127 ;
  assign n133 = n127 ^ n113 ;
  assign n134 = n133 ^ n127 ;
  assign n135 = ~n132 & ~n134 ;
  assign n136 = n135 ^ n127 ;
  assign n137 = x3 & ~n136 ;
  assign n138 = n137 ^ n127 ;
  assign n139 = ~x1 & ~n138 ;
  assign n140 = ~x3 & ~x4 ;
  assign n141 = n66 & n140 ;
  assign n142 = ~x3 & ~n68 ;
  assign n143 = n104 ^ x5 ;
  assign n144 = x4 & ~n143 ;
  assign n145 = n144 ^ x5 ;
  assign n146 = ~n142 & n145 ;
  assign n147 = ~x6 & n146 ;
  assign n148 = ~n141 & ~n147 ;
  assign n149 = x1 & n148 ;
  assign n150 = n149 ^ n139 ;
  assign n151 = ~n139 & n150 ;
  assign n152 = n151 ^ n116 ;
  assign n153 = n152 ^ n139 ;
  assign n154 = ~n119 & n153 ;
  assign n155 = n154 ^ n151 ;
  assign n156 = n155 ^ n139 ;
  assign n157 = ~n103 & ~n156 ;
  assign n158 = n157 ^ n103 ;
  assign n159 = n158 ^ n95 ;
  assign n160 = n97 & ~n159 ;
  assign n161 = n160 ^ n95 ;
  assign n162 = ~n27 & n161 ;
  assign y0 = ~n162 ;
endmodule
