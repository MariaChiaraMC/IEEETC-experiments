module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 ;
  assign n17 = x2 ^ x0 ;
  assign n32 = x1 & ~x3 ;
  assign n18 = x5 & ~x6 ;
  assign n19 = ~x4 & n18 ;
  assign n20 = x10 & ~x11 ;
  assign n21 = ~x7 & n20 ;
  assign n22 = ~x8 & ~x12 ;
  assign n23 = x9 & n22 ;
  assign n24 = n21 & n23 ;
  assign n25 = x14 & x15 ;
  assign n26 = x14 ^ x13 ;
  assign n27 = n26 ^ x15 ;
  assign n28 = n25 & n27 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n24 & n29 ;
  assign n31 = ~n19 & n30 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = x4 & x5 ;
  assign n36 = x1 & ~x6 ;
  assign n37 = n36 ^ x7 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = n36 ^ x3 ;
  assign n40 = n38 & ~n39 ;
  assign n41 = n40 ^ n36 ;
  assign n42 = n35 & n41 ;
  assign n43 = n42 ^ n31 ;
  assign n44 = ~n34 & n43 ;
  assign n45 = n44 ^ n31 ;
  assign n46 = n45 ^ x2 ;
  assign n47 = n17 & ~n46 ;
  assign n48 = n47 ^ n44 ;
  assign n49 = n48 ^ n31 ;
  assign n50 = n49 ^ x0 ;
  assign n51 = ~x2 & ~n50 ;
  assign n52 = n51 ^ x2 ;
  assign y0 = ~n52 ;
endmodule
