module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 ;
  assign n23 = x5 ^ x1 ;
  assign n24 = ~x0 & n23 ;
  assign n27 = ~x6 & x7 ;
  assign n25 = x2 & ~x3 ;
  assign n26 = ~x4 & n25 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = n27 ^ x5 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n30 ^ n24 ;
  assign n32 = n28 & ~n31 ;
  assign n33 = n32 ^ n26 ;
  assign n34 = n24 & n33 ;
  assign n35 = n34 ^ x0 ;
  assign n17 = ~x2 & ~x3 ;
  assign n18 = ~x4 & x13 ;
  assign n19 = n17 & n18 ;
  assign n36 = n35 ^ n19 ;
  assign n37 = n36 ^ n19 ;
  assign n20 = ~x9 & ~x10 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = n21 ^ n19 ;
  assign n38 = n37 ^ n22 ;
  assign n39 = x3 ^ x2 ;
  assign n40 = n39 ^ x3 ;
  assign n41 = n40 ^ x4 ;
  assign n42 = n41 ^ x4 ;
  assign n43 = ~x4 & ~x5 ;
  assign n44 = x7 & n43 ;
  assign n45 = n42 ^ n39 ;
  assign n46 = n45 ^ n42 ;
  assign n47 = n44 & ~n46 ;
  assign n48 = n47 ^ x4 ;
  assign n49 = ~x5 & n27 ;
  assign n50 = n49 ^ x4 ;
  assign n51 = ~n45 & ~n50 ;
  assign n52 = n51 ^ n42 ;
  assign n53 = n52 ^ n45 ;
  assign n54 = n48 & ~n53 ;
  assign n55 = n42 & n54 ;
  assign n56 = n55 ^ n47 ;
  assign n57 = ~x1 & n56 ;
  assign n58 = ~x3 & ~x7 ;
  assign n59 = ~x4 & ~n58 ;
  assign n60 = x5 & ~n59 ;
  assign n61 = ~x5 & x7 ;
  assign n62 = x6 & ~n61 ;
  assign n63 = ~n26 & n62 ;
  assign n64 = x4 ^ x1 ;
  assign n65 = n64 ^ x4 ;
  assign n66 = x2 & x5 ;
  assign n67 = n66 ^ x4 ;
  assign n68 = n65 & ~n67 ;
  assign n69 = n68 ^ x4 ;
  assign n70 = x3 & n69 ;
  assign n71 = n70 ^ x1 ;
  assign n72 = n63 & n71 ;
  assign n73 = ~n60 & n72 ;
  assign n74 = x0 & ~n73 ;
  assign n75 = ~n57 & n74 ;
  assign n76 = n75 ^ n19 ;
  assign n77 = n76 ^ n19 ;
  assign n78 = n77 ^ n37 ;
  assign n79 = n37 & ~n78 ;
  assign n80 = n79 ^ n37 ;
  assign n81 = n38 & n80 ;
  assign n82 = n81 ^ n79 ;
  assign n83 = n82 ^ n19 ;
  assign n84 = n83 ^ n37 ;
  assign n85 = ~x12 & n84 ;
  assign n86 = n85 ^ n19 ;
  assign n87 = ~x8 & n86 ;
  assign n15 = x12 ^ x11 ;
  assign n88 = n87 ^ n15 ;
  assign n16 = n15 ^ x12 ;
  assign n89 = n88 ^ n16 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = n90 ^ n15 ;
  assign n92 = n15 ^ x9 ;
  assign n93 = n15 ^ x10 ;
  assign n94 = n92 & n93 ;
  assign n95 = n88 ^ n15 ;
  assign n96 = ~n90 & n95 ;
  assign n97 = n96 ^ n91 ;
  assign n98 = n94 & n97 ;
  assign n99 = n98 ^ n96 ;
  assign n100 = n91 & n99 ;
  assign n101 = n100 ^ n96 ;
  assign n102 = n101 ^ x12 ;
  assign y0 = n102 ;
endmodule
