module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 ;
  assign n16 = ~x3 & ~x4 ;
  assign n17 = x1 ^ x0 ;
  assign n18 = ~x8 & ~x9 ;
  assign n19 = ~x7 & n18 ;
  assign n20 = ~x6 & ~n19 ;
  assign n21 = ~x10 & ~x11 ;
  assign n22 = ~x13 & ~x14 ;
  assign n23 = ~x7 & n22 ;
  assign n24 = n23 ^ x12 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = x14 ^ x13 ;
  assign n27 = x8 & x9 ;
  assign n28 = n27 ^ x14 ;
  assign n29 = x13 ^ x7 ;
  assign n30 = n29 ^ x14 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = ~n27 & ~n31 ;
  assign n33 = n32 ^ n27 ;
  assign n34 = n28 & ~n33 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = n35 ^ n27 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = ~n26 & ~n37 ;
  assign n39 = n38 ^ n30 ;
  assign n40 = n39 ^ n23 ;
  assign n41 = ~n25 & n40 ;
  assign n42 = n41 ^ n23 ;
  assign n43 = n21 & n42 ;
  assign n44 = n20 & ~n43 ;
  assign n45 = ~x2 & ~x5 ;
  assign n46 = ~n44 & n45 ;
  assign n47 = x1 & ~n46 ;
  assign n48 = n17 & n47 ;
  assign n49 = n48 ^ n17 ;
  assign n50 = n16 & n49 ;
  assign y0 = n50 ;
endmodule
