module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 ;
  assign n16 = x9 & ~x14 ;
  assign n17 = x8 & ~n16 ;
  assign n18 = x6 & ~x11 ;
  assign n19 = ~n17 & n18 ;
  assign n20 = x4 & x7 ;
  assign n21 = ~x13 & n20 ;
  assign n22 = n19 & n21 ;
  assign n23 = ~x8 & x9 ;
  assign n24 = x0 & x2 ;
  assign n25 = ~n23 & n24 ;
  assign n26 = ~x14 & ~n25 ;
  assign n27 = ~x12 & ~n26 ;
  assign n28 = n22 & n27 ;
  assign n29 = x3 & ~x5 ;
  assign n30 = ~x1 & x10 ;
  assign n31 = n30 ^ x14 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = x1 & ~x10 ;
  assign n34 = x9 & ~n33 ;
  assign n35 = ~x0 & ~x2 ;
  assign n36 = ~n34 & n35 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = n32 & n37 ;
  assign n39 = n38 ^ n30 ;
  assign n40 = ~x9 & ~n30 ;
  assign n41 = n40 ^ n29 ;
  assign n42 = ~n39 & n41 ;
  assign n43 = n42 ^ n40 ;
  assign n44 = n29 & n43 ;
  assign n45 = n44 ^ n29 ;
  assign n46 = n28 & n45 ;
  assign y0 = n46 ;
endmodule
