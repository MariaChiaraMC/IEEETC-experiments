module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 ;
  assign n30 = x9 & ~x10 ;
  assign n15 = ~x6 & x13 ;
  assign n16 = ~x11 & n15 ;
  assign n31 = n30 ^ n16 ;
  assign n39 = n31 ^ n16 ;
  assign n17 = x3 & x8 ;
  assign n18 = n17 ^ x6 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = n17 ^ x0 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n19 & n21 ;
  assign n23 = n22 ^ n17 ;
  assign n24 = x10 & n23 ;
  assign n25 = n24 ^ n17 ;
  assign n26 = ~x9 & n25 ;
  assign n27 = ~x11 & ~n26 ;
  assign n28 = ~x13 & ~n27 ;
  assign n29 = n28 ^ n16 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = n33 ^ n16 ;
  assign n35 = n32 ^ x12 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = n34 & ~n37 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = n40 ^ n34 ;
  assign n42 = ~x6 & x10 ;
  assign n43 = x8 & n42 ;
  assign n44 = x11 & ~n43 ;
  assign n45 = ~x9 & ~n44 ;
  assign n46 = n45 ^ n16 ;
  assign n47 = n38 ^ n34 ;
  assign n48 = ~n46 & n47 ;
  assign n49 = n48 ^ n16 ;
  assign n50 = n41 & ~n49 ;
  assign n51 = n50 ^ n16 ;
  assign n52 = n51 ^ n30 ;
  assign n53 = n52 ^ n16 ;
  assign y0 = n53 ;
endmodule
