module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 ;
  assign n9 = ~x5 & ~x6 ;
  assign n10 = x1 & n9 ;
  assign n11 = x0 & ~x1 ;
  assign n12 = x6 & x7 ;
  assign n13 = n11 & n12 ;
  assign n14 = ~x5 & n13 ;
  assign n15 = ~n10 & ~n14 ;
  assign n16 = ~x3 & ~x4 ;
  assign n17 = ~n15 & n16 ;
  assign n18 = ~x2 & n17 ;
  assign n21 = ~x1 & ~x2 ;
  assign n22 = x6 & ~x7 ;
  assign n23 = ~x4 & n22 ;
  assign n24 = x4 & ~x6 ;
  assign n25 = ~n23 & ~n24 ;
  assign n26 = n21 & ~n25 ;
  assign n27 = ~x6 & x7 ;
  assign n19 = ~x2 & x4 ;
  assign n28 = n19 & n22 ;
  assign n29 = ~n27 & ~n28 ;
  assign n30 = x1 & ~n29 ;
  assign n31 = ~n26 & ~n30 ;
  assign n20 = n12 & n19 ;
  assign n32 = n31 ^ n20 ;
  assign n33 = x5 & ~n32 ;
  assign n34 = n33 ^ n31 ;
  assign n47 = ~n23 & ~n27 ;
  assign n48 = ~x2 & ~x4 ;
  assign n49 = n47 & ~n48 ;
  assign n35 = x7 ^ x1 ;
  assign n36 = n35 ^ x2 ;
  assign n37 = n36 ^ n9 ;
  assign n38 = x2 ^ x1 ;
  assign n39 = n38 ^ x5 ;
  assign n40 = ~x5 & n39 ;
  assign n41 = n40 ^ x2 ;
  assign n42 = n41 ^ x5 ;
  assign n43 = n37 & n42 ;
  assign n44 = n43 ^ n40 ;
  assign n45 = n44 ^ x5 ;
  assign n46 = ~n9 & ~n45 ;
  assign n50 = n49 ^ n46 ;
  assign n51 = n50 ^ x1 ;
  assign n58 = n51 ^ n50 ;
  assign n52 = n51 ^ x4 ;
  assign n53 = n52 ^ n50 ;
  assign n54 = n51 ^ n49 ;
  assign n55 = n54 ^ x4 ;
  assign n56 = n55 ^ n53 ;
  assign n57 = ~n53 & n56 ;
  assign n59 = n58 ^ n57 ;
  assign n60 = n59 ^ n53 ;
  assign n61 = n50 ^ n9 ;
  assign n62 = n57 ^ n53 ;
  assign n63 = ~n61 & ~n62 ;
  assign n64 = n63 ^ n50 ;
  assign n65 = ~n60 & n64 ;
  assign n66 = n65 ^ n50 ;
  assign n67 = n66 ^ n46 ;
  assign n68 = n67 ^ n50 ;
  assign n69 = n68 ^ x3 ;
  assign n70 = n69 ^ n68 ;
  assign n76 = x5 ^ x4 ;
  assign n77 = n76 ^ x7 ;
  assign n71 = n38 ^ x4 ;
  assign n87 = n77 ^ n71 ;
  assign n88 = n87 ^ x2 ;
  assign n78 = n77 ^ x5 ;
  assign n79 = n78 ^ n71 ;
  assign n101 = n88 ^ n79 ;
  assign n90 = n71 ^ x7 ;
  assign n91 = n90 ^ n77 ;
  assign n92 = n91 ^ x5 ;
  assign n93 = n92 ^ n77 ;
  assign n94 = n93 ^ n71 ;
  assign n102 = n101 ^ n94 ;
  assign n103 = n94 ^ n79 ;
  assign n72 = x6 ^ x5 ;
  assign n73 = n72 ^ n71 ;
  assign n74 = n73 ^ x2 ;
  assign n81 = n74 ^ n71 ;
  assign n82 = n81 ^ n79 ;
  assign n83 = n82 ^ x2 ;
  assign n104 = n103 ^ n83 ;
  assign n75 = n74 ^ x2 ;
  assign n80 = n79 ^ n75 ;
  assign n84 = n83 ^ n80 ;
  assign n85 = n84 ^ n74 ;
  assign n86 = n85 ^ n79 ;
  assign n89 = n88 ^ n86 ;
  assign n95 = n94 ^ n89 ;
  assign n96 = n95 ^ n83 ;
  assign n105 = n104 ^ n96 ;
  assign n106 = ~n102 & ~n105 ;
  assign n97 = n96 ^ n83 ;
  assign n98 = n94 ^ n83 ;
  assign n99 = n98 ^ n96 ;
  assign n100 = ~n97 & ~n99 ;
  assign n107 = n106 ^ n100 ;
  assign n108 = n107 ^ n74 ;
  assign n109 = n108 ^ n83 ;
  assign n110 = n109 ^ n96 ;
  assign n111 = n100 ^ n88 ;
  assign n112 = n111 ^ n96 ;
  assign n113 = n103 ^ n96 ;
  assign n114 = n88 ^ n74 ;
  assign n115 = n114 ^ n83 ;
  assign n116 = n113 & ~n115 ;
  assign n117 = n116 ^ n79 ;
  assign n118 = n117 ^ n94 ;
  assign n119 = ~n112 & n118 ;
  assign n120 = n119 ^ n79 ;
  assign n121 = n120 ^ n88 ;
  assign n122 = n121 ^ n96 ;
  assign n123 = n110 & ~n122 ;
  assign n124 = n123 ^ n116 ;
  assign n125 = n124 ^ n119 ;
  assign n126 = n125 ^ n74 ;
  assign n127 = n126 ^ n94 ;
  assign n128 = n127 ^ n83 ;
  assign n129 = n128 ^ x4 ;
  assign n130 = n129 ^ n84 ;
  assign n131 = n130 ^ n68 ;
  assign n132 = n70 & ~n131 ;
  assign n133 = n132 ^ n68 ;
  assign n134 = n34 & n133 ;
  assign n135 = ~x0 & ~n134 ;
  assign n136 = x5 & ~x7 ;
  assign n137 = x3 & n136 ;
  assign n138 = n24 & n137 ;
  assign n139 = n21 & n138 ;
  assign n140 = ~n135 & ~n139 ;
  assign n141 = ~n18 & n140 ;
  assign y0 = ~n141 ;
endmodule
