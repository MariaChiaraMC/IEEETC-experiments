module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 ;
  assign n8 = x2 ^ x1 ;
  assign n9 = x4 ^ x3 ;
  assign n10 = n9 ^ x3 ;
  assign n11 = ~x5 & ~x6 ;
  assign n12 = n11 ^ x3 ;
  assign n13 = ~n10 & ~n12 ;
  assign n14 = n13 ^ x3 ;
  assign n15 = n14 ^ x2 ;
  assign n16 = ~n8 & ~n15 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n17 ^ x3 ;
  assign n19 = n18 ^ x1 ;
  assign n20 = x2 & n19 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = ~x0 & n21 ;
  assign y0 = ~n22 ;
endmodule
