module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 ;
  assign n11 = ~x5 & x7 ;
  assign n12 = ~x2 & n11 ;
  assign n13 = ~x0 & x3 ;
  assign n14 = n12 & n13 ;
  assign n15 = x6 & n14 ;
  assign n16 = ~x0 & x4 ;
  assign n17 = x2 & ~x7 ;
  assign n18 = ~x5 & ~x6 ;
  assign n19 = n17 & n18 ;
  assign n20 = x3 & ~n19 ;
  assign n21 = n16 & ~n20 ;
  assign n22 = ~x2 & x7 ;
  assign n23 = x6 & n22 ;
  assign n24 = n23 ^ x2 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = x6 & ~x7 ;
  assign n27 = ~x3 & ~n26 ;
  assign n28 = n27 ^ n23 ;
  assign n29 = n28 ^ n23 ;
  assign n30 = n25 & ~n29 ;
  assign n31 = n30 ^ n23 ;
  assign n32 = ~x5 & n31 ;
  assign n33 = n32 ^ n23 ;
  assign n34 = n21 & n33 ;
  assign n35 = ~x3 & ~x4 ;
  assign n36 = x5 & ~x7 ;
  assign n37 = n36 ^ n18 ;
  assign n38 = n37 ^ n18 ;
  assign n39 = n18 ^ x6 ;
  assign n40 = n39 ^ n18 ;
  assign n41 = n38 & n40 ;
  assign n42 = n41 ^ n18 ;
  assign n43 = x0 & n42 ;
  assign n44 = n43 ^ n18 ;
  assign n45 = n35 & n44 ;
  assign n46 = x2 & n45 ;
  assign n47 = ~n34 & ~n46 ;
  assign n48 = x3 & ~x4 ;
  assign n52 = x6 ^ x5 ;
  assign n49 = x6 ^ x0 ;
  assign n50 = n49 ^ x7 ;
  assign n59 = n52 ^ n50 ;
  assign n51 = n50 ^ x6 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n52 ^ x2 ;
  assign n55 = n54 ^ x7 ;
  assign n56 = n55 ^ x6 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n53 & ~n57 ;
  assign n60 = n59 ^ n58 ;
  assign n61 = n60 ^ n53 ;
  assign n62 = n52 ^ x7 ;
  assign n63 = n58 ^ n53 ;
  assign n64 = n62 & n63 ;
  assign n65 = n64 ^ n52 ;
  assign n66 = n61 & n65 ;
  assign n67 = n66 ^ n52 ;
  assign n68 = n67 ^ n52 ;
  assign n69 = n48 & n68 ;
  assign n70 = n47 & ~n69 ;
  assign n71 = ~n15 & n70 ;
  assign n72 = x9 & ~n71 ;
  assign n73 = ~x0 & ~n36 ;
  assign n74 = x3 & ~n11 ;
  assign n75 = ~n73 & n74 ;
  assign n76 = ~x2 & ~x6 ;
  assign n77 = ~x4 & ~x5 ;
  assign n78 = n77 ^ x9 ;
  assign n79 = n76 & ~n78 ;
  assign n80 = n79 ^ x9 ;
  assign n81 = n75 & ~n80 ;
  assign n82 = x6 ^ x4 ;
  assign n83 = n82 ^ x2 ;
  assign n84 = x6 ^ x2 ;
  assign n85 = n26 ^ x2 ;
  assign n86 = ~x2 & n85 ;
  assign n87 = n86 ^ x2 ;
  assign n88 = n84 & ~n87 ;
  assign n89 = n88 ^ n86 ;
  assign n90 = n89 ^ x2 ;
  assign n91 = n90 ^ n26 ;
  assign n92 = n83 & n91 ;
  assign n93 = n92 ^ n26 ;
  assign n94 = n81 & ~n93 ;
  assign n95 = ~x7 & ~x9 ;
  assign n96 = ~x0 & x2 ;
  assign n97 = n95 & n96 ;
  assign n98 = ~x3 & n97 ;
  assign n99 = n77 & n98 ;
  assign n100 = ~n94 & ~n99 ;
  assign n101 = ~n72 & n100 ;
  assign n102 = x1 & ~n101 ;
  assign n127 = x4 & x6 ;
  assign n128 = x9 & ~n127 ;
  assign n129 = x7 & ~n128 ;
  assign n130 = x2 ^ x0 ;
  assign n131 = x9 ^ x3 ;
  assign n132 = n131 ^ x9 ;
  assign n133 = n132 ^ n130 ;
  assign n134 = x4 ^ x2 ;
  assign n135 = x4 & ~n134 ;
  assign n136 = n135 ^ x9 ;
  assign n137 = n136 ^ x4 ;
  assign n138 = ~n133 & ~n137 ;
  assign n139 = n138 ^ n135 ;
  assign n140 = n139 ^ x4 ;
  assign n141 = n130 & n140 ;
  assign n142 = n141 ^ n130 ;
  assign n143 = n142 ^ x6 ;
  assign n144 = n143 ^ n142 ;
  assign n103 = ~x2 & ~x4 ;
  assign n145 = x3 ^ x0 ;
  assign n146 = n103 & ~n145 ;
  assign n147 = n146 ^ n142 ;
  assign n148 = ~n144 & n147 ;
  assign n149 = n148 ^ n142 ;
  assign n150 = n129 & n149 ;
  assign n151 = n48 ^ n17 ;
  assign n152 = x9 ^ x0 ;
  assign n153 = n152 ^ x0 ;
  assign n154 = ~x0 & x6 ;
  assign n155 = n154 ^ x0 ;
  assign n156 = ~n153 & n155 ;
  assign n157 = n156 ^ x0 ;
  assign n158 = n157 ^ n48 ;
  assign n159 = n151 & n158 ;
  assign n160 = n159 ^ n156 ;
  assign n161 = n160 ^ x0 ;
  assign n162 = n161 ^ n17 ;
  assign n163 = n48 & n162 ;
  assign n164 = n163 ^ n48 ;
  assign n165 = ~n150 & ~n164 ;
  assign n166 = ~x1 & ~n165 ;
  assign n123 = ~x7 & x9 ;
  assign n167 = n13 & n127 ;
  assign n168 = n123 & n167 ;
  assign n169 = ~x2 & n168 ;
  assign n170 = ~n166 & ~n169 ;
  assign n104 = n95 & n103 ;
  assign n105 = x2 & x9 ;
  assign n106 = x4 & x7 ;
  assign n107 = n106 ^ x3 ;
  assign n108 = n107 ^ n106 ;
  assign n109 = ~x4 & ~x7 ;
  assign n110 = n109 ^ n106 ;
  assign n111 = ~n108 & n110 ;
  assign n112 = n111 ^ n106 ;
  assign n113 = n105 & n112 ;
  assign n114 = ~n104 & ~n113 ;
  assign n115 = ~x6 & ~n114 ;
  assign n116 = x2 & x6 ;
  assign n117 = ~x3 & ~x9 ;
  assign n118 = ~n116 & n117 ;
  assign n119 = n106 & n118 ;
  assign n120 = ~n115 & ~n119 ;
  assign n121 = ~x1 & ~n120 ;
  assign n122 = ~x3 & x4 ;
  assign n124 = n122 & n123 ;
  assign n125 = n76 & n124 ;
  assign n126 = ~n121 & ~n125 ;
  assign n171 = n170 ^ n126 ;
  assign n172 = n171 ^ n170 ;
  assign n173 = n170 ^ x0 ;
  assign n174 = n173 ^ n170 ;
  assign n175 = ~n172 & n174 ;
  assign n176 = n175 ^ n170 ;
  assign n177 = x5 & ~n176 ;
  assign n178 = n177 ^ n170 ;
  assign n179 = ~n102 & n178 ;
  assign n180 = ~x8 & ~n179 ;
  assign n181 = ~x2 & x5 ;
  assign n182 = n26 & n181 ;
  assign n183 = x2 & ~x5 ;
  assign n184 = ~x6 & x7 ;
  assign n185 = n183 & n184 ;
  assign n186 = ~n182 & ~n185 ;
  assign n187 = x1 & ~x4 ;
  assign n188 = ~x9 & n187 ;
  assign n189 = ~n186 & n188 ;
  assign n190 = ~x1 & x2 ;
  assign n191 = x7 & x9 ;
  assign n192 = n127 & n191 ;
  assign n193 = n190 & n192 ;
  assign n194 = ~x5 & n193 ;
  assign n195 = ~n189 & ~n194 ;
  assign n196 = n13 & ~n195 ;
  assign n197 = x0 & ~x2 ;
  assign n198 = n191 & n197 ;
  assign n199 = ~n97 & ~n198 ;
  assign n200 = ~x5 & ~n199 ;
  assign n201 = ~x0 & x9 ;
  assign n202 = x2 & x5 ;
  assign n203 = ~x7 & n202 ;
  assign n204 = n201 & n203 ;
  assign n205 = ~n200 & ~n204 ;
  assign n206 = x1 & ~n205 ;
  assign n207 = ~n17 & ~n22 ;
  assign n208 = x0 & ~x1 ;
  assign n209 = ~x5 & ~n191 ;
  assign n210 = n208 & n209 ;
  assign n211 = ~n207 & n210 ;
  assign n212 = ~n206 & ~n211 ;
  assign n213 = n127 & ~n212 ;
  assign n214 = n77 & n184 ;
  assign n215 = ~n182 & ~n214 ;
  assign n216 = x1 & ~n215 ;
  assign n217 = n216 ^ x2 ;
  assign n218 = n217 ^ n216 ;
  assign n219 = x1 & ~x6 ;
  assign n220 = x5 & x7 ;
  assign n221 = ~x4 & n220 ;
  assign n222 = n219 & n221 ;
  assign n223 = ~x1 & ~x7 ;
  assign n224 = n52 ^ x6 ;
  assign n225 = ~x4 & ~x6 ;
  assign n226 = n225 ^ x6 ;
  assign n227 = n224 & n226 ;
  assign n228 = n227 ^ x6 ;
  assign n229 = n223 & n228 ;
  assign n230 = ~n222 & ~n229 ;
  assign n231 = n230 ^ n216 ;
  assign n232 = n231 ^ n216 ;
  assign n233 = n218 & ~n232 ;
  assign n234 = n233 ^ n216 ;
  assign n235 = x9 & n234 ;
  assign n236 = n235 ^ n216 ;
  assign n237 = ~x0 & n236 ;
  assign n239 = ~x1 & ~n184 ;
  assign n240 = x4 & n202 ;
  assign n241 = ~n239 & n240 ;
  assign n238 = n197 & n222 ;
  assign n242 = n241 ^ n238 ;
  assign n243 = n242 ^ n238 ;
  assign n244 = x7 ^ x1 ;
  assign n245 = x0 & n244 ;
  assign n246 = n245 ^ x1 ;
  assign n247 = n246 ^ n238 ;
  assign n248 = n247 ^ n238 ;
  assign n249 = n243 & ~n248 ;
  assign n250 = n249 ^ n238 ;
  assign n251 = ~x9 & n250 ;
  assign n252 = n251 ^ n238 ;
  assign n253 = ~n237 & ~n252 ;
  assign n254 = ~n213 & n253 ;
  assign n255 = n254 ^ x3 ;
  assign n256 = n255 ^ n254 ;
  assign n258 = ~x5 & ~x7 ;
  assign n257 = x1 ^ x0 ;
  assign n259 = n258 ^ n257 ;
  assign n260 = n259 ^ x4 ;
  assign n261 = n260 ^ n259 ;
  assign n262 = n261 ^ n257 ;
  assign n263 = n257 ^ n220 ;
  assign n264 = x1 & ~n263 ;
  assign n265 = n259 ^ n257 ;
  assign n266 = n261 & n265 ;
  assign n267 = n266 ^ n262 ;
  assign n268 = n264 & n267 ;
  assign n269 = n268 ^ n266 ;
  assign n270 = n262 & n269 ;
  assign n271 = n270 ^ n266 ;
  assign n272 = n76 & n271 ;
  assign n273 = x0 & x7 ;
  assign n274 = ~x6 & n190 ;
  assign n275 = n77 & n274 ;
  assign n276 = n273 & n275 ;
  assign n277 = x0 & x6 ;
  assign n278 = n187 & n277 ;
  assign n279 = n203 & n278 ;
  assign n280 = ~x9 & ~n279 ;
  assign n281 = ~n276 & n280 ;
  assign n282 = ~n12 & ~n203 ;
  assign n283 = x4 & ~n282 ;
  assign n284 = n283 ^ x2 ;
  assign n285 = n284 ^ n283 ;
  assign n286 = n283 ^ n220 ;
  assign n287 = n286 ^ n283 ;
  assign n288 = n285 & n287 ;
  assign n289 = n288 ^ n283 ;
  assign n290 = ~x1 & n289 ;
  assign n291 = n290 ^ n283 ;
  assign n292 = n154 & n291 ;
  assign n293 = n281 & ~n292 ;
  assign n294 = ~n272 & n293 ;
  assign n295 = n183 ^ n181 ;
  assign n296 = x7 ^ x4 ;
  assign n297 = n181 ^ x7 ;
  assign n298 = n296 & n297 ;
  assign n299 = n298 ^ x7 ;
  assign n300 = n295 & ~n299 ;
  assign n301 = n300 ^ n183 ;
  assign n302 = n219 & n301 ;
  assign n303 = n77 & n239 ;
  assign n304 = ~n207 & n303 ;
  assign n305 = ~n302 & ~n304 ;
  assign n306 = ~x0 & ~n305 ;
  assign n307 = x4 & n208 ;
  assign n308 = ~n181 & ~n183 ;
  assign n309 = ~n76 & n308 ;
  assign n310 = n309 ^ n184 ;
  assign n311 = n310 ^ n184 ;
  assign n312 = n184 ^ x7 ;
  assign n313 = n311 & ~n312 ;
  assign n314 = n313 ^ n184 ;
  assign n315 = n307 & n314 ;
  assign n316 = x9 & ~n315 ;
  assign n317 = ~n306 & n316 ;
  assign n318 = ~n294 & ~n317 ;
  assign n319 = n318 ^ n254 ;
  assign n320 = ~n256 & ~n319 ;
  assign n321 = n320 ^ n254 ;
  assign n322 = x8 & ~n321 ;
  assign n323 = ~n196 & ~n322 ;
  assign n324 = ~n180 & n323 ;
  assign y0 = ~n324 ;
endmodule
