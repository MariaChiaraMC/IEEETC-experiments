module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n17 = ~x0 & ~x2 ;
  assign n18 = ~x3 & n17 ;
  assign n19 = x6 & n18 ;
  assign n20 = ~x1 & n19 ;
  assign n21 = ~x4 & ~x7 ;
  assign n22 = x11 ^ x10 ;
  assign n23 = n21 & n22 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = x4 & x7 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = n25 & n27 ;
  assign n29 = n28 ^ n23 ;
  assign n30 = n20 & n29 ;
  assign y0 = n30 ;
endmodule
