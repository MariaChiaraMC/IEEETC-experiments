module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n15 = ~x9 & ~x12 ;
  assign n16 = ~x4 & n15 ;
  assign n17 = ~x5 & ~x13 ;
  assign n18 = ~x8 & n17 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = ~x6 & x10 ;
  assign n21 = n20 ^ x11 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = x3 & ~x10 ;
  assign n24 = n23 ^ n20 ;
  assign n25 = ~n22 & n24 ;
  assign n26 = n25 ^ n20 ;
  assign n27 = n26 ^ n16 ;
  assign n28 = n19 & n27 ;
  assign n29 = n28 ^ n25 ;
  assign n30 = n29 ^ n20 ;
  assign n31 = n30 ^ n18 ;
  assign n32 = n16 & n31 ;
  assign n33 = n32 ^ n16 ;
  assign y0 = n33 ;
endmodule
