module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 ;
  assign n10 = ~x0 & ~x7 ;
  assign n11 = x6 & ~x8 ;
  assign n12 = x5 & n11 ;
  assign n13 = n12 ^ x3 ;
  assign n21 = n13 ^ n12 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = ~x6 & x8 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = ~n15 & ~n19 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n22 ^ n15 ;
  assign n24 = n12 ^ x1 ;
  assign n25 = n20 ^ n15 ;
  assign n26 = ~n24 & ~n25 ;
  assign n27 = n26 ^ n12 ;
  assign n28 = n23 & ~n27 ;
  assign n29 = n28 ^ n12 ;
  assign n30 = n29 ^ x3 ;
  assign n31 = n30 ^ n12 ;
  assign n32 = n10 & ~n31 ;
  assign n45 = x0 & ~x1 ;
  assign n38 = x3 & ~x6 ;
  assign n46 = ~x7 & n38 ;
  assign n47 = n46 ^ x3 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = x6 & x7 ;
  assign n50 = ~x6 & ~x7 ;
  assign n51 = ~n49 & ~n50 ;
  assign n52 = n51 ^ n46 ;
  assign n53 = n52 ^ n46 ;
  assign n54 = ~n48 & ~n53 ;
  assign n55 = n54 ^ n46 ;
  assign n56 = ~x8 & n55 ;
  assign n57 = n56 ^ n46 ;
  assign n58 = n45 & n57 ;
  assign n33 = ~x0 & x7 ;
  assign n34 = x8 & n33 ;
  assign n35 = x3 & x6 ;
  assign n36 = n35 ^ x1 ;
  assign n37 = n36 ^ n35 ;
  assign n39 = ~x3 & x6 ;
  assign n40 = ~n38 & ~n39 ;
  assign n41 = n40 ^ n35 ;
  assign n42 = n37 & ~n41 ;
  assign n43 = n42 ^ n35 ;
  assign n44 = n34 & n43 ;
  assign n59 = n58 ^ n44 ;
  assign n60 = n59 ^ x5 ;
  assign n67 = n60 ^ n59 ;
  assign n61 = n60 ^ n45 ;
  assign n62 = n61 ^ n59 ;
  assign n63 = n60 ^ n58 ;
  assign n64 = n63 ^ n45 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = n62 & n65 ;
  assign n68 = n67 ^ n66 ;
  assign n69 = n68 ^ n62 ;
  assign n70 = x7 & ~x8 ;
  assign n71 = ~x6 & n70 ;
  assign n72 = n71 ^ n59 ;
  assign n73 = n66 ^ n62 ;
  assign n74 = n72 & n73 ;
  assign n75 = n74 ^ n59 ;
  assign n76 = n69 & n75 ;
  assign n77 = n76 ^ n59 ;
  assign n78 = n77 ^ n44 ;
  assign n79 = n78 ^ n59 ;
  assign n80 = ~n32 & ~n79 ;
  assign n81 = n80 ^ x4 ;
  assign n82 = n81 ^ n80 ;
  assign n98 = ~x3 & n11 ;
  assign n105 = ~x5 & ~x7 ;
  assign n106 = x5 & x7 ;
  assign n107 = ~n105 & ~n106 ;
  assign n108 = n98 & n107 ;
  assign n109 = ~n10 & n108 ;
  assign n110 = x6 ^ x0 ;
  assign n111 = n110 ^ n105 ;
  assign n120 = n111 ^ n105 ;
  assign n121 = n106 ^ x6 ;
  assign n122 = n121 ^ n105 ;
  assign n123 = n122 ^ n120 ;
  assign n124 = n120 & n123 ;
  assign n112 = n111 ^ x6 ;
  assign n113 = n112 ^ n105 ;
  assign n114 = n105 ^ x3 ;
  assign n115 = n114 ^ n113 ;
  assign n116 = n113 & ~n115 ;
  assign n129 = n124 ^ n116 ;
  assign n117 = n116 ^ n111 ;
  assign n118 = n117 ^ n113 ;
  assign n119 = n118 ^ x8 ;
  assign n125 = n124 ^ n113 ;
  assign n126 = n125 ^ n120 ;
  assign n127 = n126 ^ x8 ;
  assign n128 = n119 & ~n127 ;
  assign n130 = n129 ^ n128 ;
  assign n131 = ~x8 & n130 ;
  assign n132 = n131 ^ n124 ;
  assign n133 = n132 ^ n116 ;
  assign n134 = n133 ^ n128 ;
  assign n135 = ~n39 & n134 ;
  assign n136 = ~n109 & ~n135 ;
  assign n83 = x3 & x5 ;
  assign n84 = ~x3 & ~x5 ;
  assign n85 = x8 & n84 ;
  assign n86 = ~n83 & ~n85 ;
  assign n87 = x8 ^ x6 ;
  assign n88 = n10 & ~n87 ;
  assign n89 = ~n86 & n88 ;
  assign n90 = x7 & ~n84 ;
  assign n91 = x5 ^ x3 ;
  assign n92 = ~x8 & n91 ;
  assign n93 = n92 ^ x3 ;
  assign n94 = ~x6 & ~n93 ;
  assign n95 = n94 ^ x0 ;
  assign n96 = n95 ^ n94 ;
  assign n97 = ~x5 & n16 ;
  assign n99 = ~n97 & ~n98 ;
  assign n100 = n99 ^ n94 ;
  assign n101 = n96 & ~n100 ;
  assign n102 = n101 ^ n94 ;
  assign n103 = n90 & n102 ;
  assign n104 = ~n89 & ~n103 ;
  assign n137 = n136 ^ n104 ;
  assign n138 = x1 & n137 ;
  assign n139 = n138 ^ n136 ;
  assign n140 = n139 ^ n80 ;
  assign n141 = ~n82 & n140 ;
  assign n142 = n141 ^ n80 ;
  assign n143 = x2 & ~n142 ;
  assign n144 = ~x4 & x5 ;
  assign n145 = n38 & n144 ;
  assign n146 = ~x2 & x8 ;
  assign n147 = n33 & n146 ;
  assign n148 = n145 & n147 ;
  assign n149 = n148 ^ n143 ;
  assign n150 = n49 & n84 ;
  assign n151 = n150 ^ x0 ;
  assign n152 = n151 ^ n150 ;
  assign n153 = n150 ^ x7 ;
  assign n154 = n152 & ~n153 ;
  assign n155 = n154 ^ x7 ;
  assign n158 = ~x4 & x6 ;
  assign n156 = n150 ^ x3 ;
  assign n157 = n156 ^ n151 ;
  assign n159 = n158 ^ n157 ;
  assign n160 = n159 ^ n157 ;
  assign n161 = n157 ^ n151 ;
  assign n162 = n161 ^ n150 ;
  assign n163 = n162 ^ n154 ;
  assign n164 = n160 & ~n163 ;
  assign n165 = n164 ^ n145 ;
  assign n166 = ~x7 & n165 ;
  assign n167 = n166 ^ n164 ;
  assign n168 = n167 ^ n152 ;
  assign n169 = ~n155 & n168 ;
  assign n170 = n169 ^ n164 ;
  assign n171 = n170 ^ n166 ;
  assign n172 = n171 ^ n152 ;
  assign n173 = n172 ^ x0 ;
  assign n174 = n146 & n173 ;
  assign n176 = x4 & n49 ;
  assign n177 = n176 ^ n83 ;
  assign n175 = n83 ^ x2 ;
  assign n178 = n177 ^ n175 ;
  assign n179 = n178 ^ n177 ;
  assign n180 = n179 ^ n83 ;
  assign n181 = x6 ^ x4 ;
  assign n182 = n105 ^ x6 ;
  assign n183 = n182 ^ n105 ;
  assign n184 = n107 ^ n105 ;
  assign n185 = ~n183 & n184 ;
  assign n186 = n185 ^ n105 ;
  assign n187 = n181 & n186 ;
  assign n188 = n187 ^ n178 ;
  assign n189 = x3 & n188 ;
  assign n190 = n177 ^ n83 ;
  assign n191 = n179 & n190 ;
  assign n192 = n191 ^ n180 ;
  assign n193 = n189 & ~n192 ;
  assign n194 = n193 ^ n191 ;
  assign n195 = ~n180 & n194 ;
  assign n196 = n195 ^ n191 ;
  assign n197 = n196 ^ n176 ;
  assign n198 = ~x8 & n197 ;
  assign n199 = ~x0 & n198 ;
  assign n200 = ~x8 & n105 ;
  assign n201 = ~n158 & n200 ;
  assign n202 = ~x0 & x2 ;
  assign n203 = n201 & ~n202 ;
  assign n204 = x0 & ~x2 ;
  assign n205 = n204 ^ x4 ;
  assign n206 = n205 ^ n203 ;
  assign n207 = x4 ^ x3 ;
  assign n208 = n207 ^ n181 ;
  assign n209 = ~n181 & n208 ;
  assign n210 = n209 ^ x4 ;
  assign n211 = n210 ^ n181 ;
  assign n212 = ~n206 & n211 ;
  assign n213 = n212 ^ n209 ;
  assign n214 = n213 ^ n181 ;
  assign n215 = n203 & ~n214 ;
  assign n216 = ~n199 & ~n215 ;
  assign n217 = ~n174 & n216 ;
  assign n218 = n217 ^ x1 ;
  assign n219 = n218 ^ n217 ;
  assign n220 = ~x2 & ~x3 ;
  assign n221 = x4 & x5 ;
  assign n222 = n71 & n221 ;
  assign n223 = n220 & n222 ;
  assign n224 = n146 & n221 ;
  assign n225 = n46 & n224 ;
  assign n226 = n70 & n158 ;
  assign n227 = n84 & n226 ;
  assign n228 = ~n225 & ~n227 ;
  assign n229 = n228 ^ x0 ;
  assign n230 = n229 ^ n228 ;
  assign n231 = n230 ^ n223 ;
  assign n232 = x8 & n105 ;
  assign n233 = n232 ^ n144 ;
  assign n234 = n233 ^ n232 ;
  assign n235 = n232 ^ n70 ;
  assign n236 = n235 ^ n232 ;
  assign n237 = n234 & n236 ;
  assign n238 = n237 ^ n232 ;
  assign n239 = ~x6 & n238 ;
  assign n240 = n239 ^ n232 ;
  assign n241 = x3 & n240 ;
  assign n242 = x8 & n106 ;
  assign n243 = ~n200 & ~n242 ;
  assign n244 = x4 & n38 ;
  assign n245 = ~n39 & ~n244 ;
  assign n246 = ~n243 & ~n245 ;
  assign n247 = ~x3 & x8 ;
  assign n248 = n50 & n144 ;
  assign n249 = n247 & n248 ;
  assign n250 = ~n246 & ~n249 ;
  assign n251 = ~n241 & n250 ;
  assign n252 = n251 ^ x2 ;
  assign n253 = ~x2 & n252 ;
  assign n254 = n253 ^ n228 ;
  assign n255 = n254 ^ x2 ;
  assign n256 = ~n231 & n255 ;
  assign n257 = n256 ^ n253 ;
  assign n258 = n257 ^ x2 ;
  assign n259 = ~n223 & ~n258 ;
  assign n260 = n259 ^ n223 ;
  assign n261 = n260 ^ n217 ;
  assign n262 = ~n219 & ~n261 ;
  assign n263 = n262 ^ n217 ;
  assign n264 = n263 ^ n143 ;
  assign n265 = n149 & ~n264 ;
  assign n266 = n265 ^ n262 ;
  assign n267 = n266 ^ n217 ;
  assign n268 = n267 ^ n148 ;
  assign n269 = ~n143 & ~n268 ;
  assign n270 = n269 ^ n143 ;
  assign y0 = n270 ;
endmodule
