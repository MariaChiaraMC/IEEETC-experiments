module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 ;
  assign n9 = x5 & x6 ;
  assign n10 = ~x3 & ~n9 ;
  assign n11 = x2 & ~n10 ;
  assign n12 = ~x4 & n11 ;
  assign n13 = ~x3 & ~x4 ;
  assign n14 = ~n9 & ~n13 ;
  assign n15 = ~x4 & x5 ;
  assign n16 = ~x2 & ~n15 ;
  assign n17 = ~n14 & n16 ;
  assign n18 = x5 & x7 ;
  assign n19 = n18 ^ x5 ;
  assign n20 = n19 ^ x4 ;
  assign n28 = n20 ^ n19 ;
  assign n21 = x2 & ~x7 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n20 ^ n18 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n23 & n26 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = n19 ^ x3 ;
  assign n32 = n27 ^ n23 ;
  assign n33 = ~n31 & n32 ;
  assign n34 = n33 ^ n19 ;
  assign n35 = ~n30 & ~n34 ;
  assign n36 = n35 ^ n19 ;
  assign n37 = n36 ^ x5 ;
  assign n38 = n37 ^ n19 ;
  assign n39 = ~x6 & ~n38 ;
  assign n40 = ~n17 & ~n39 ;
  assign n41 = ~n12 & n40 ;
  assign n42 = ~x1 & ~n41 ;
  assign n43 = n18 ^ x4 ;
  assign n44 = x4 ^ x3 ;
  assign n45 = n44 ^ x4 ;
  assign n46 = ~n43 & n45 ;
  assign n47 = n46 ^ x4 ;
  assign n48 = x1 & n47 ;
  assign n52 = x7 ^ x4 ;
  assign n49 = n44 ^ x5 ;
  assign n50 = n49 ^ n44 ;
  assign n51 = n50 ^ x4 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n44 ^ x7 ;
  assign n55 = n54 ^ x4 ;
  assign n56 = n55 ^ x4 ;
  assign n57 = ~n50 & ~n56 ;
  assign n58 = n57 ^ n50 ;
  assign n59 = n55 & ~n58 ;
  assign n60 = n59 ^ x4 ;
  assign n61 = n53 & ~n60 ;
  assign n62 = n61 ^ n57 ;
  assign n63 = n62 ^ x4 ;
  assign n64 = n63 ^ x3 ;
  assign n65 = n64 ^ n52 ;
  assign n66 = n65 ^ x6 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = n67 ^ n48 ;
  assign n69 = ~x3 & ~x7 ;
  assign n70 = x1 & ~x4 ;
  assign n71 = ~n69 & ~n70 ;
  assign n72 = n71 ^ x5 ;
  assign n73 = x5 & ~n72 ;
  assign n74 = n73 ^ n65 ;
  assign n75 = n74 ^ x5 ;
  assign n76 = ~n68 & ~n75 ;
  assign n77 = n76 ^ n73 ;
  assign n78 = n77 ^ x5 ;
  assign n79 = ~n48 & n78 ;
  assign n80 = n79 ^ n48 ;
  assign n81 = ~x2 & n80 ;
  assign n82 = ~n42 & ~n81 ;
  assign y0 = ~n82 ;
endmodule
