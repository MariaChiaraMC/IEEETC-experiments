module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 ;
  assign n15 = ~x1 & ~x2 ;
  assign n16 = ~x5 & ~n15 ;
  assign n17 = x1 & x6 ;
  assign n18 = n17 ^ x3 ;
  assign n19 = x4 & ~n18 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = ~n16 & ~n20 ;
  assign n22 = x5 & n15 ;
  assign n23 = x1 & ~x4 ;
  assign n24 = ~x8 & ~x11 ;
  assign n25 = ~x10 & ~x12 ;
  assign n26 = ~x7 & ~x9 ;
  assign n27 = n25 & ~n26 ;
  assign n28 = x3 & ~x13 ;
  assign n29 = n27 & n28 ;
  assign n30 = n24 & n29 ;
  assign n31 = ~n23 & ~n30 ;
  assign n32 = n31 ^ x2 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = n33 ^ n22 ;
  assign n35 = x6 ^ x3 ;
  assign n36 = ~x3 & ~n35 ;
  assign n37 = n36 ^ n31 ;
  assign n38 = n37 ^ x3 ;
  assign n39 = n34 & n38 ;
  assign n40 = n39 ^ n36 ;
  assign n41 = n40 ^ x3 ;
  assign n42 = ~n22 & ~n41 ;
  assign n43 = n42 ^ n22 ;
  assign n44 = n21 & ~n43 ;
  assign n45 = ~x0 & ~n44 ;
  assign y0 = n45 ;
endmodule
