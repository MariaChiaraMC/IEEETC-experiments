module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 ;
  assign n15 = ~x4 & x11 ;
  assign n16 = x5 & x6 ;
  assign n17 = n15 & n16 ;
  assign n18 = x3 ^ x2 ;
  assign n19 = ~x7 & n18 ;
  assign n20 = n19 ^ x2 ;
  assign n21 = n17 & n20 ;
  assign n22 = ~x2 & ~x8 ;
  assign n23 = x1 & n22 ;
  assign n24 = ~x11 & n23 ;
  assign n25 = ~n21 & ~n24 ;
  assign n26 = ~x12 & ~x13 ;
  assign n27 = ~n25 & n26 ;
  assign n28 = ~x5 & x12 ;
  assign n29 = ~x6 & n28 ;
  assign n30 = n20 & ~n29 ;
  assign n31 = ~x13 & ~n28 ;
  assign n32 = x6 & x13 ;
  assign n33 = ~n31 & ~n32 ;
  assign n34 = x5 & ~x12 ;
  assign n35 = x11 ^ x4 ;
  assign n36 = ~n34 & ~n35 ;
  assign n37 = n33 & n36 ;
  assign n38 = n30 & n37 ;
  assign n39 = ~n27 & ~n38 ;
  assign n40 = x2 & ~x7 ;
  assign n41 = x13 ^ x6 ;
  assign n44 = ~n28 & n36 ;
  assign n42 = ~x4 & ~x5 ;
  assign n43 = ~x11 & n42 ;
  assign n45 = n44 ^ n43 ;
  assign n46 = n45 ^ n44 ;
  assign n47 = n46 ^ n41 ;
  assign n48 = x13 ^ x12 ;
  assign n49 = ~x12 & ~n48 ;
  assign n50 = n49 ^ n44 ;
  assign n51 = n50 ^ x12 ;
  assign n52 = ~n47 & ~n51 ;
  assign n53 = n52 ^ n49 ;
  assign n54 = n53 ^ x12 ;
  assign n55 = ~n41 & ~n54 ;
  assign n56 = n40 & n55 ;
  assign n57 = n39 & ~n56 ;
  assign n58 = ~x9 & ~x10 ;
  assign n59 = ~x0 & n58 ;
  assign n60 = ~n57 & n59 ;
  assign y0 = n60 ;
endmodule
