module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ;
  assign n18 = x15 ^ x12 ;
  assign n19 = x15 ^ x13 ;
  assign n20 = n19 ^ x13 ;
  assign n21 = x16 ^ x13 ;
  assign n22 = n20 & ~n21 ;
  assign n23 = n22 ^ x13 ;
  assign n24 = ~n18 & ~n23 ;
  assign n25 = n24 ^ x12 ;
  assign n26 = x14 & ~n25 ;
  assign n27 = x15 & x16 ;
  assign n28 = ~x14 & ~n27 ;
  assign n29 = ~x0 & ~n28 ;
  assign n30 = x12 ^ x11 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = ~x7 & x10 ;
  assign n33 = ~x16 & n32 ;
  assign n34 = ~x11 & n33 ;
  assign n35 = n34 ^ n29 ;
  assign n36 = n31 & n35 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = n29 & n37 ;
  assign n39 = ~n26 & n38 ;
  assign y0 = n39 ;
endmodule
