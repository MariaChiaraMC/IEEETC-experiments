module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;
  assign n8 = ~x5 & ~x6 ;
  assign n9 = x5 & x6 ;
  assign n10 = ~x0 & ~x1 ;
  assign n11 = x2 & ~n10 ;
  assign n12 = n9 & ~n11 ;
  assign n13 = n12 ^ x3 ;
  assign n14 = n13 ^ x3 ;
  assign n15 = n14 ^ n8 ;
  assign n31 = x2 & x6 ;
  assign n32 = x5 & n10 ;
  assign n33 = ~x2 & n32 ;
  assign n34 = x4 & ~n33 ;
  assign n35 = ~n31 & n34 ;
  assign n17 = x6 ^ x4 ;
  assign n16 = x5 ^ x4 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = n19 ^ x4 ;
  assign n21 = x4 ^ x2 ;
  assign n22 = x4 ^ x1 ;
  assign n23 = n21 & n22 ;
  assign n24 = n17 ^ x4 ;
  assign n25 = ~n19 & ~n24 ;
  assign n26 = n25 ^ n20 ;
  assign n27 = n23 & ~n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = ~n20 & n28 ;
  assign n30 = n29 ^ n25 ;
  assign n36 = n35 ^ n30 ;
  assign n37 = ~x3 & n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = n15 & ~n38 ;
  assign n40 = n39 ^ n37 ;
  assign n41 = n40 ^ n35 ;
  assign n42 = n41 ^ x3 ;
  assign n43 = ~n8 & n42 ;
  assign y0 = ~n43 ;
endmodule
