module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 ;
  assign n25 = x4 & ~x5 ;
  assign n26 = x10 & n25 ;
  assign n27 = ~x1 & n26 ;
  assign n28 = x1 & x5 ;
  assign n29 = ~x18 & n28 ;
  assign n30 = x4 & ~x17 ;
  assign n31 = ~x23 & ~n30 ;
  assign n32 = n29 & ~n31 ;
  assign n33 = ~n27 & ~n32 ;
  assign n34 = ~x14 & ~x15 ;
  assign n35 = x16 & ~n34 ;
  assign n36 = x2 & ~n35 ;
  assign n37 = ~n33 & n36 ;
  assign n38 = x14 & x15 ;
  assign n39 = x16 & n38 ;
  assign n40 = x11 & ~n39 ;
  assign n41 = x1 & ~x2 ;
  assign n42 = n26 & n41 ;
  assign n43 = n40 & n42 ;
  assign n44 = ~x18 & n43 ;
  assign n45 = ~n37 & ~n44 ;
  assign n46 = ~x0 & ~n45 ;
  assign n47 = x2 & n29 ;
  assign n48 = ~x0 & n47 ;
  assign n49 = ~n31 & ~n38 ;
  assign n50 = x7 & ~x17 ;
  assign n51 = ~n49 & ~n50 ;
  assign n52 = n48 & ~n51 ;
  assign n53 = ~x18 & n25 ;
  assign n54 = ~n39 & n53 ;
  assign n55 = ~x7 & ~n54 ;
  assign n56 = ~x1 & ~x2 ;
  assign n57 = ~x9 & n56 ;
  assign n58 = ~n55 & n57 ;
  assign n59 = ~n52 & ~n58 ;
  assign n60 = n59 ^ x3 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = ~x2 & x8 ;
  assign n63 = n25 & ~n35 ;
  assign n64 = ~x6 & ~n63 ;
  assign n65 = n56 & ~n64 ;
  assign n66 = ~n62 & ~n65 ;
  assign n69 = n66 ^ n47 ;
  assign n70 = n69 ^ n66 ;
  assign n67 = n66 ^ x17 ;
  assign n68 = n67 ^ n66 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = n66 ^ x6 ;
  assign n73 = n72 ^ n66 ;
  assign n74 = n73 ^ n70 ;
  assign n75 = n70 & n74 ;
  assign n76 = n75 ^ n70 ;
  assign n77 = ~n71 & n76 ;
  assign n78 = n77 ^ n75 ;
  assign n79 = n78 ^ n66 ;
  assign n80 = n79 ^ n70 ;
  assign n81 = ~x0 & ~n80 ;
  assign n82 = n81 ^ n66 ;
  assign n83 = n82 ^ n59 ;
  assign n84 = ~n61 & n83 ;
  assign n85 = n84 ^ n59 ;
  assign n86 = ~n46 & n85 ;
  assign n87 = x13 & ~n86 ;
  assign y0 = n87 ;
endmodule
