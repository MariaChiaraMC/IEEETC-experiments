module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 ;
  assign n22 = ~x0 & ~x2 ;
  assign n23 = ~x4 & n22 ;
  assign n24 = x3 & ~x5 ;
  assign n25 = x1 & ~n24 ;
  assign n26 = n23 & n25 ;
  assign n27 = x0 & ~x1 ;
  assign n28 = ~x2 & ~x3 ;
  assign n29 = ~x4 & x5 ;
  assign n30 = ~n28 & n29 ;
  assign n31 = n27 & n30 ;
  assign n32 = ~x2 & ~x11 ;
  assign n33 = x9 ^ x0 ;
  assign n34 = x9 ^ x1 ;
  assign n35 = n34 ^ x1 ;
  assign n36 = ~x1 & x3 ;
  assign n37 = n36 ^ x1 ;
  assign n38 = n35 & n37 ;
  assign n39 = n38 ^ x1 ;
  assign n40 = ~n33 & n39 ;
  assign n41 = n40 ^ x0 ;
  assign n42 = n32 & ~n41 ;
  assign n43 = ~x5 & ~n42 ;
  assign n44 = ~x9 & ~x10 ;
  assign n45 = n44 ^ x11 ;
  assign n46 = x12 & ~x13 ;
  assign n47 = ~x8 & ~n46 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = ~x6 & ~x7 ;
  assign n50 = n49 ^ x11 ;
  assign n51 = x13 ^ x11 ;
  assign n52 = n51 ^ x11 ;
  assign n53 = n50 & ~n52 ;
  assign n54 = n53 ^ x11 ;
  assign n55 = n54 ^ n45 ;
  assign n56 = ~n48 & ~n55 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n57 ^ x11 ;
  assign n59 = n58 ^ n47 ;
  assign n60 = ~n45 & n59 ;
  assign n61 = n60 ^ n45 ;
  assign n62 = ~n43 & ~n61 ;
  assign n63 = ~x12 & ~x13 ;
  assign n64 = ~x2 & x5 ;
  assign n65 = x10 & ~x11 ;
  assign n66 = x5 & n65 ;
  assign n67 = x11 & n49 ;
  assign n68 = ~x10 & n67 ;
  assign n69 = n68 ^ n36 ;
  assign n70 = n68 ^ n22 ;
  assign n71 = n70 ^ n22 ;
  assign n72 = x10 & n32 ;
  assign n73 = n72 ^ n22 ;
  assign n74 = ~n71 & ~n73 ;
  assign n75 = n74 ^ n22 ;
  assign n76 = n69 & n75 ;
  assign n77 = n76 ^ n36 ;
  assign n78 = ~n66 & ~n77 ;
  assign n79 = x8 & ~n78 ;
  assign n80 = ~n64 & ~n79 ;
  assign n81 = n63 & ~n80 ;
  assign n82 = x9 & n81 ;
  assign n83 = ~n62 & ~n82 ;
  assign n84 = ~x4 & ~n83 ;
  assign n85 = ~x0 & ~x1 ;
  assign n86 = x2 & ~n85 ;
  assign n87 = ~n65 & ~n68 ;
  assign n88 = x9 & ~n87 ;
  assign n89 = x8 & ~n88 ;
  assign n90 = n89 ^ n86 ;
  assign n92 = ~x8 & x11 ;
  assign n91 = ~x1 & n44 ;
  assign n93 = n92 ^ n91 ;
  assign n94 = n93 ^ n91 ;
  assign n95 = ~n44 & n49 ;
  assign n96 = ~x8 & ~n95 ;
  assign n97 = ~x4 & n63 ;
  assign n98 = ~n96 & n97 ;
  assign n99 = n98 ^ n91 ;
  assign n100 = ~n94 & n99 ;
  assign n101 = n100 ^ n91 ;
  assign n102 = n101 ^ n86 ;
  assign n103 = ~n90 & n102 ;
  assign n104 = n103 ^ n100 ;
  assign n105 = n104 ^ n91 ;
  assign n106 = n105 ^ n89 ;
  assign n107 = n86 & ~n106 ;
  assign n108 = n107 ^ n86 ;
  assign n109 = ~x5 & ~n108 ;
  assign n110 = x9 & x10 ;
  assign n111 = ~n44 & ~n110 ;
  assign n112 = ~x8 & ~x12 ;
  assign n113 = ~n92 & ~n112 ;
  assign n114 = ~n111 & ~n113 ;
  assign n115 = ~x15 & ~n114 ;
  assign n116 = ~x6 & ~n115 ;
  assign n117 = n116 ^ x2 ;
  assign n118 = n117 ^ n116 ;
  assign n119 = ~x10 & ~x11 ;
  assign n120 = ~x8 & x9 ;
  assign n121 = n119 & n120 ;
  assign n122 = x12 & ~n121 ;
  assign n123 = n122 ^ n116 ;
  assign n124 = ~n118 & n123 ;
  assign n125 = n124 ^ n116 ;
  assign n126 = ~x1 & n125 ;
  assign n127 = x13 & ~n126 ;
  assign n128 = x10 & n49 ;
  assign n129 = n128 ^ x7 ;
  assign n130 = n128 ^ x16 ;
  assign n131 = n128 ^ x8 ;
  assign n132 = n128 & n131 ;
  assign n133 = n132 ^ n128 ;
  assign n134 = n130 & n133 ;
  assign n135 = n134 ^ n132 ;
  assign n136 = n135 ^ n128 ;
  assign n137 = n136 ^ x8 ;
  assign n138 = n129 & n137 ;
  assign n139 = n138 ^ n128 ;
  assign n140 = n111 & n139 ;
  assign n141 = x11 & n140 ;
  assign n142 = x12 ^ x6 ;
  assign n143 = x10 & ~x15 ;
  assign n144 = ~n121 & ~n143 ;
  assign n145 = n144 ^ x12 ;
  assign n146 = n144 ^ x7 ;
  assign n147 = n144 & ~n146 ;
  assign n148 = n147 ^ n144 ;
  assign n149 = ~n145 & n148 ;
  assign n150 = n149 ^ n147 ;
  assign n151 = n150 ^ n144 ;
  assign n152 = n151 ^ x7 ;
  assign n153 = ~n142 & ~n152 ;
  assign n154 = n153 ^ x12 ;
  assign n155 = ~n141 & ~n154 ;
  assign n156 = ~x13 & ~n155 ;
  assign n157 = x6 & x9 ;
  assign n158 = x7 & n157 ;
  assign n159 = ~x13 & ~n49 ;
  assign n160 = ~x16 & ~n159 ;
  assign n161 = ~x13 & ~n112 ;
  assign n162 = x9 & ~n161 ;
  assign n163 = ~n160 & ~n162 ;
  assign n164 = ~x15 & ~n163 ;
  assign n165 = ~n158 & ~n164 ;
  assign n166 = x11 & ~n165 ;
  assign n167 = ~x13 & n65 ;
  assign n168 = ~x9 & n167 ;
  assign n169 = x15 & ~n168 ;
  assign n170 = n49 & ~n169 ;
  assign n171 = x10 & n158 ;
  assign n172 = x9 & ~x12 ;
  assign n173 = n143 & n172 ;
  assign n174 = ~n171 & ~n173 ;
  assign n175 = ~n170 & n174 ;
  assign n176 = x8 & ~n175 ;
  assign n177 = ~x17 & ~n176 ;
  assign n178 = ~n166 & n177 ;
  assign n179 = ~n156 & n178 ;
  assign n180 = x2 & ~n179 ;
  assign n181 = ~x2 & n110 ;
  assign n182 = x11 & n181 ;
  assign n183 = x13 & x16 ;
  assign n184 = x7 & n44 ;
  assign n185 = n183 & n184 ;
  assign n186 = n92 & n185 ;
  assign n187 = ~n182 & ~n186 ;
  assign n188 = ~x12 & ~n187 ;
  assign n189 = x4 & ~n27 ;
  assign n190 = ~n188 & n189 ;
  assign n191 = ~n180 & n190 ;
  assign n192 = ~n127 & n191 ;
  assign n193 = ~n109 & ~n192 ;
  assign n194 = x1 & x5 ;
  assign n195 = ~x0 & n194 ;
  assign n196 = ~n23 & ~n195 ;
  assign n197 = ~n193 & n196 ;
  assign n198 = ~x3 & ~n197 ;
  assign n199 = x4 & ~x5 ;
  assign n200 = n27 & n199 ;
  assign n201 = x4 ^ x2 ;
  assign n202 = n201 ^ x4 ;
  assign n203 = n202 ^ n201 ;
  assign n204 = n203 ^ x5 ;
  assign n205 = n203 & ~n204 ;
  assign n206 = n205 ^ n202 ;
  assign n207 = n206 ^ n203 ;
  assign n208 = n201 ^ x3 ;
  assign n214 = n208 ^ x0 ;
  assign n209 = n208 ^ n201 ;
  assign n210 = n209 ^ n202 ;
  assign n211 = n210 ^ n203 ;
  assign n212 = n202 & n211 ;
  assign n213 = n212 ^ n209 ;
  assign n215 = n214 ^ n213 ;
  assign n216 = n209 ^ x20 ;
  assign n217 = n216 ^ n214 ;
  assign n218 = ~x20 & n217 ;
  assign n219 = n218 ^ n202 ;
  assign n220 = ~n215 & n219 ;
  assign n221 = n220 ^ n209 ;
  assign n222 = n221 ^ n203 ;
  assign n223 = n222 ^ x5 ;
  assign n224 = n207 & ~n223 ;
  assign n225 = n224 ^ n212 ;
  assign n226 = n225 ^ n220 ;
  assign n227 = n226 ^ n202 ;
  assign n228 = n227 ^ x2 ;
  assign n229 = n228 ^ x1 ;
  assign n230 = n229 ^ n228 ;
  assign n231 = n230 ^ n200 ;
  assign n232 = n92 & n172 ;
  assign n233 = ~x3 & ~n232 ;
  assign n234 = n233 ^ n64 ;
  assign n235 = ~n233 & ~n234 ;
  assign n236 = n235 ^ n228 ;
  assign n237 = n236 ^ n233 ;
  assign n238 = n231 & ~n237 ;
  assign n239 = n238 ^ n235 ;
  assign n240 = n239 ^ n233 ;
  assign n241 = ~n200 & ~n240 ;
  assign n242 = n241 ^ n200 ;
  assign n243 = ~n198 & ~n242 ;
  assign n244 = ~n84 & n243 ;
  assign n245 = ~x19 & ~n244 ;
  assign n246 = ~x18 & n245 ;
  assign n247 = ~n31 & ~n246 ;
  assign n248 = ~n26 & n247 ;
  assign n249 = x14 & ~n248 ;
  assign y0 = n249 ;
endmodule
