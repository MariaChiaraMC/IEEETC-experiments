module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 ;
  output y0 ;
  wire n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 ;
  assign n23 = ~x0 & x2 ;
  assign n24 = x1 & x5 ;
  assign n25 = n23 & n24 ;
  assign n26 = x13 & x14 ;
  assign n27 = ~x12 & n26 ;
  assign n28 = ~x3 & n27 ;
  assign n29 = x12 & x14 ;
  assign n30 = n29 ^ x15 ;
  assign n31 = n30 ^ x15 ;
  assign n32 = x15 ^ x3 ;
  assign n33 = n31 & ~n32 ;
  assign n34 = n33 ^ x15 ;
  assign n35 = ~x13 & x15 ;
  assign n36 = n35 ^ x16 ;
  assign n37 = n34 & ~n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = ~x16 & n38 ;
  assign n40 = n39 ^ x16 ;
  assign n41 = ~n28 & n40 ;
  assign n42 = n25 & ~n41 ;
  assign n45 = ~x15 & n26 ;
  assign n43 = x9 & n23 ;
  assign n44 = ~x1 & n43 ;
  assign n46 = n45 ^ n44 ;
  assign n47 = n44 ^ x16 ;
  assign n48 = n47 ^ x16 ;
  assign n49 = ~x1 & ~x2 ;
  assign n50 = x0 & n49 ;
  assign n51 = ~x3 & n50 ;
  assign n52 = n51 ^ x16 ;
  assign n53 = ~n48 & n52 ;
  assign n54 = n53 ^ x16 ;
  assign n55 = ~n46 & ~n54 ;
  assign n56 = n55 ^ n45 ;
  assign n57 = ~n29 & ~n56 ;
  assign n58 = x3 & ~x8 ;
  assign n59 = n58 ^ x10 ;
  assign n60 = n59 ^ n58 ;
  assign n61 = ~x0 & x9 ;
  assign n62 = n61 ^ n58 ;
  assign n63 = n62 ^ n58 ;
  assign n64 = n60 & n63 ;
  assign n65 = n64 ^ n58 ;
  assign n66 = x1 & n65 ;
  assign n67 = n66 ^ n58 ;
  assign n68 = ~x2 & n67 ;
  assign n69 = n68 ^ x16 ;
  assign n70 = x13 & x15 ;
  assign n71 = n29 & n70 ;
  assign n72 = n71 ^ n68 ;
  assign n73 = n72 ^ n71 ;
  assign n74 = ~x8 & ~x12 ;
  assign n75 = n50 & n74 ;
  assign n76 = n75 ^ n71 ;
  assign n77 = ~n73 & ~n76 ;
  assign n78 = n77 ^ n71 ;
  assign n79 = ~n69 & n78 ;
  assign n80 = n79 ^ x16 ;
  assign n81 = ~n57 & n80 ;
  assign n82 = ~x5 & ~n81 ;
  assign n83 = ~n42 & ~n82 ;
  assign n84 = x4 & ~n83 ;
  assign n85 = x16 ^ x13 ;
  assign n86 = ~x15 & ~n85 ;
  assign n87 = n86 ^ x13 ;
  assign n88 = n25 & n87 ;
  assign n89 = ~x8 & n49 ;
  assign n90 = ~n88 & ~n89 ;
  assign n91 = x3 & x7 ;
  assign n92 = ~n90 & n91 ;
  assign n93 = n50 ^ x6 ;
  assign n94 = n93 ^ x3 ;
  assign n95 = n88 ^ x8 ;
  assign n96 = x6 & ~n95 ;
  assign n97 = n96 ^ x8 ;
  assign n98 = ~n94 & n97 ;
  assign n99 = n98 ^ n96 ;
  assign n100 = n99 ^ x8 ;
  assign n101 = n100 ^ x6 ;
  assign n102 = ~x3 & n101 ;
  assign n103 = ~n92 & ~n102 ;
  assign n104 = ~n84 & n103 ;
  assign n21 = ~x17 & ~x18 ;
  assign n22 = x19 & n21 ;
  assign n105 = n104 ^ n22 ;
  assign n106 = ~x11 & ~n105 ;
  assign n107 = n106 ^ n104 ;
  assign y0 = ~n107 ;
endmodule
