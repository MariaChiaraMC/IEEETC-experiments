module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 ;
  assign n16 = ~x7 & x10 ;
  assign n17 = x3 & x14 ;
  assign n18 = x6 & ~n17 ;
  assign n19 = ~x8 & ~n18 ;
  assign n20 = n16 & ~n19 ;
  assign n21 = x12 ^ x11 ;
  assign n22 = x9 & ~x13 ;
  assign n23 = ~x0 & n22 ;
  assign n24 = n23 ^ x12 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = ~x3 & ~x6 ;
  assign n28 = x13 & x14 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n27 & n29 ;
  assign n31 = n30 ^ n23 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = n26 & n32 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ n27 ;
  assign n36 = n21 & n35 ;
  assign n37 = n20 & n36 ;
  assign n38 = x0 & x14 ;
  assign n39 = x3 & x8 ;
  assign n40 = n22 & n39 ;
  assign n41 = ~x10 & ~x11 ;
  assign n42 = x6 & n41 ;
  assign n43 = n40 & n42 ;
  assign n44 = ~n38 & n43 ;
  assign n45 = ~n37 & ~n44 ;
  assign n46 = ~x4 & ~n45 ;
  assign n47 = ~x5 & n46 ;
  assign n48 = x14 ^ x10 ;
  assign n49 = x14 ^ x13 ;
  assign n50 = n49 ^ n48 ;
  assign n51 = x11 ^ x4 ;
  assign n52 = x13 & n51 ;
  assign n53 = n52 ^ x4 ;
  assign n54 = n50 & n53 ;
  assign n55 = n54 ^ n52 ;
  assign n56 = n55 ^ x4 ;
  assign n57 = n56 ^ x13 ;
  assign n58 = n48 & n57 ;
  assign n59 = n58 ^ x10 ;
  assign n60 = ~x3 & ~n59 ;
  assign n61 = x11 & x14 ;
  assign n62 = n61 ^ x10 ;
  assign n63 = n62 ^ n61 ;
  assign n64 = ~x0 & x4 ;
  assign n65 = ~x13 & x14 ;
  assign n70 = ~x11 & ~n65 ;
  assign n66 = x3 & ~x8 ;
  assign n67 = ~x1 & ~x6 ;
  assign n68 = ~n66 & ~n67 ;
  assign n69 = n65 & n68 ;
  assign n71 = n70 ^ n69 ;
  assign n72 = n69 ^ x7 ;
  assign n73 = n69 ^ x5 ;
  assign n74 = ~n69 & ~n73 ;
  assign n75 = n74 ^ n69 ;
  assign n76 = ~n72 & ~n75 ;
  assign n77 = n76 ^ n74 ;
  assign n78 = n77 ^ n69 ;
  assign n79 = n78 ^ x5 ;
  assign n80 = n71 & ~n79 ;
  assign n81 = n80 ^ n70 ;
  assign n82 = n64 & n81 ;
  assign n83 = x5 & x6 ;
  assign n84 = n70 & n83 ;
  assign n85 = x7 & n84 ;
  assign n86 = x4 & n85 ;
  assign n87 = ~x11 & x13 ;
  assign n88 = n87 ^ x4 ;
  assign n89 = n88 ^ x14 ;
  assign n92 = ~x5 & ~x6 ;
  assign n93 = x7 & ~x13 ;
  assign n94 = x8 & x11 ;
  assign n95 = n93 & n94 ;
  assign n96 = n92 & n95 ;
  assign n90 = x1 & x7 ;
  assign n91 = ~x5 & n90 ;
  assign n97 = n96 ^ n91 ;
  assign n98 = ~x4 & n97 ;
  assign n99 = n98 ^ n91 ;
  assign n100 = n89 & ~n99 ;
  assign n101 = n100 ^ n98 ;
  assign n102 = n101 ^ n91 ;
  assign n103 = n102 ^ x4 ;
  assign n104 = ~x14 & n103 ;
  assign n105 = ~n86 & ~n104 ;
  assign n106 = ~n82 & n105 ;
  assign n107 = n106 ^ n61 ;
  assign n108 = n63 & ~n107 ;
  assign n109 = n108 ^ n61 ;
  assign n110 = ~n39 & n64 ;
  assign n111 = x5 & ~x13 ;
  assign n112 = x3 & ~n67 ;
  assign n113 = n111 & ~n112 ;
  assign n114 = n110 & n113 ;
  assign n115 = n61 & n114 ;
  assign n116 = n115 ^ n60 ;
  assign n117 = n109 & ~n116 ;
  assign n118 = n117 ^ n115 ;
  assign n119 = ~n60 & n118 ;
  assign n120 = n119 ^ n60 ;
  assign n121 = ~x12 & n120 ;
  assign n122 = ~x4 & x14 ;
  assign n123 = n122 ^ x11 ;
  assign n124 = ~x8 & n93 ;
  assign n125 = ~x7 & x8 ;
  assign n126 = n87 & n125 ;
  assign n127 = ~n124 & ~n126 ;
  assign n128 = n92 & ~n127 ;
  assign n129 = n128 ^ n123 ;
  assign n130 = n129 ^ n122 ;
  assign n131 = n130 ^ n129 ;
  assign n132 = x13 & ~x14 ;
  assign n133 = n91 & n132 ;
  assign n134 = ~x2 & n111 ;
  assign n135 = ~n67 & n134 ;
  assign n136 = ~n133 & ~n135 ;
  assign n137 = n64 & ~n66 ;
  assign n138 = ~n136 & n137 ;
  assign n139 = n138 ^ n129 ;
  assign n140 = n139 ^ n123 ;
  assign n141 = n131 & ~n140 ;
  assign n142 = n141 ^ n138 ;
  assign n143 = x13 & ~n138 ;
  assign n144 = n143 ^ n123 ;
  assign n145 = ~n142 & ~n144 ;
  assign n146 = n145 ^ n143 ;
  assign n147 = ~n123 & n146 ;
  assign n148 = n147 ^ n141 ;
  assign n149 = n148 ^ x11 ;
  assign n150 = n149 ^ n138 ;
  assign n151 = x10 & ~n150 ;
  assign n153 = n151 ^ x12 ;
  assign n162 = n153 ^ n151 ;
  assign n152 = n151 ^ n41 ;
  assign n154 = n153 ^ n152 ;
  assign n155 = n154 ^ n153 ;
  assign n156 = n155 ^ n151 ;
  assign n157 = n154 ^ x14 ;
  assign n158 = n157 ^ x3 ;
  assign n159 = n158 ^ n154 ;
  assign n160 = n159 ^ n156 ;
  assign n161 = n156 & ~n160 ;
  assign n163 = n162 ^ n161 ;
  assign n164 = n163 ^ n156 ;
  assign n165 = n151 ^ x3 ;
  assign n166 = n161 ^ n156 ;
  assign n167 = n165 & n166 ;
  assign n168 = n167 ^ n151 ;
  assign n169 = n164 & ~n168 ;
  assign n170 = n169 ^ n151 ;
  assign n171 = n170 ^ x12 ;
  assign n172 = n171 ^ n151 ;
  assign n173 = ~n121 & ~n172 ;
  assign n174 = ~x9 & ~n173 ;
  assign n175 = x11 & ~x12 ;
  assign n176 = ~x1 & n38 ;
  assign n177 = ~x13 & ~n176 ;
  assign n178 = n175 & ~n177 ;
  assign n179 = ~x3 & n61 ;
  assign n180 = ~x13 & ~n179 ;
  assign n181 = x14 ^ x7 ;
  assign n187 = n181 ^ x14 ;
  assign n182 = n181 ^ x8 ;
  assign n183 = n182 ^ x14 ;
  assign n184 = x13 ^ x8 ;
  assign n185 = n184 ^ n183 ;
  assign n186 = n183 & ~n185 ;
  assign n188 = n187 ^ n186 ;
  assign n189 = n188 ^ n183 ;
  assign n190 = x14 ^ x6 ;
  assign n191 = n186 ^ n183 ;
  assign n192 = n190 & n191 ;
  assign n193 = n192 ^ x14 ;
  assign n194 = n189 & n193 ;
  assign n195 = n194 ^ x14 ;
  assign n196 = n195 ^ x7 ;
  assign n197 = n196 ^ x14 ;
  assign n198 = ~n180 & ~n197 ;
  assign n199 = x12 & ~n198 ;
  assign n200 = n199 ^ x9 ;
  assign n201 = n200 ^ n199 ;
  assign n202 = ~x11 & x12 ;
  assign n203 = n202 ^ n199 ;
  assign n204 = n203 ^ n200 ;
  assign n205 = n204 ^ x13 ;
  assign n211 = n205 ^ n200 ;
  assign n212 = n211 ^ n199 ;
  assign n206 = n205 ^ x14 ;
  assign n207 = n206 ^ x13 ;
  assign n208 = n207 ^ n206 ;
  assign n209 = n208 ^ n199 ;
  assign n210 = n209 ^ n201 ;
  assign n213 = n212 ^ n210 ;
  assign n214 = n201 & n213 ;
  assign n215 = n214 ^ n208 ;
  assign n216 = n215 ^ n212 ;
  assign n222 = n206 ^ n205 ;
  assign n217 = x0 & ~x11 ;
  assign n218 = n217 ^ n206 ;
  assign n219 = n212 ^ n208 ;
  assign n220 = n218 & n219 ;
  assign n221 = n220 ^ n214 ;
  assign n223 = n222 ^ n221 ;
  assign n224 = n223 ^ n218 ;
  assign n225 = n224 ^ n208 ;
  assign n226 = n212 & ~n225 ;
  assign n227 = n226 ^ n201 ;
  assign n228 = n216 & n227 ;
  assign n229 = n228 ^ n201 ;
  assign n230 = n229 ^ x9 ;
  assign n231 = n230 ^ n201 ;
  assign n232 = ~n178 & ~n231 ;
  assign n233 = ~x10 & ~n232 ;
  assign n234 = ~x10 & x12 ;
  assign n235 = n22 & n125 ;
  assign n236 = n234 & n235 ;
  assign n237 = n92 & n236 ;
  assign n238 = ~n233 & ~n237 ;
  assign n239 = ~n174 & n238 ;
  assign n240 = ~n47 & n239 ;
  assign y0 = ~n240 ;
endmodule
