module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 ;
  assign n33 = ~x24 & ~x30 ;
  assign n34 = ~x27 & n33 ;
  assign n35 = ~x25 & ~x31 ;
  assign n36 = ~x26 & n35 ;
  assign n37 = ~x5 & ~x6 ;
  assign n38 = ~x0 & ~x15 ;
  assign n39 = n37 & n38 ;
  assign n40 = n36 & n39 ;
  assign n41 = n34 & n40 ;
  assign n42 = ~x4 & ~x7 ;
  assign n43 = ~x2 & ~x13 ;
  assign n44 = n42 & n43 ;
  assign n45 = ~x11 & ~x21 ;
  assign n46 = n44 & n45 ;
  assign n47 = ~x20 & ~x23 ;
  assign n48 = ~x1 & ~x14 ;
  assign n49 = n47 & n48 ;
  assign n50 = ~x9 & ~x10 ;
  assign n51 = ~x8 & ~x22 ;
  assign n52 = n50 & n51 ;
  assign n53 = n49 & n52 ;
  assign n54 = n46 & n53 ;
  assign n55 = ~x17 & ~x29 ;
  assign n56 = ~x18 & n55 ;
  assign n57 = ~x19 & ~x28 ;
  assign n58 = ~x16 & n57 ;
  assign n59 = n56 & n58 ;
  assign n60 = ~x3 & ~x12 ;
  assign n61 = n59 & n60 ;
  assign n62 = n54 & n61 ;
  assign n63 = n41 & n62 ;
  assign y0 = n63 ;
endmodule
