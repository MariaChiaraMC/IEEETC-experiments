module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 ;
  assign n60 = x5 ^ x4 ;
  assign n61 = n60 ^ x2 ;
  assign n58 = x6 ^ x5 ;
  assign n46 = x6 ^ x3 ;
  assign n57 = n46 ^ x2 ;
  assign n59 = n58 ^ n57 ;
  assign n62 = n61 ^ n59 ;
  assign n63 = n62 ^ n61 ;
  assign n64 = n63 ^ n57 ;
  assign n65 = x6 ^ x2 ;
  assign n66 = n65 ^ n57 ;
  assign n67 = n66 ^ n61 ;
  assign n68 = n67 ^ n64 ;
  assign n69 = n68 ^ x6 ;
  assign n70 = n69 ^ n61 ;
  assign n71 = n70 ^ n57 ;
  assign n72 = n71 ^ x6 ;
  assign n78 = n72 ^ x6 ;
  assign n79 = n78 ^ n64 ;
  assign n80 = n79 ^ n69 ;
  assign n81 = n64 & n80 ;
  assign n73 = n72 ^ n64 ;
  assign n74 = n64 ^ n57 ;
  assign n75 = n74 ^ n64 ;
  assign n76 = n75 ^ n72 ;
  assign n77 = ~n73 & ~n76 ;
  assign n82 = n81 ^ n77 ;
  assign n83 = n82 ^ n64 ;
  assign n84 = n83 ^ n72 ;
  assign n85 = n78 ^ n72 ;
  assign n86 = n77 ^ n74 ;
  assign n87 = n86 ^ n72 ;
  assign n88 = n85 & ~n87 ;
  assign n89 = n88 ^ n77 ;
  assign n90 = n89 ^ n64 ;
  assign n91 = n90 ^ n78 ;
  assign n92 = n91 ^ n69 ;
  assign n93 = ~n84 & n92 ;
  assign n94 = n93 ^ n88 ;
  assign n95 = ~x1 & n94 ;
  assign n102 = ~x2 & ~x6 ;
  assign n100 = x1 & x5 ;
  assign n28 = x4 & ~x5 ;
  assign n96 = x2 & ~x5 ;
  assign n97 = x1 & ~x6 ;
  assign n98 = n96 & n97 ;
  assign n99 = ~n28 & ~n98 ;
  assign n101 = n100 ^ n99 ;
  assign n103 = n102 ^ n101 ;
  assign n104 = n103 ^ n99 ;
  assign n109 = n104 ^ n101 ;
  assign n110 = n109 ^ n99 ;
  assign n111 = n110 ^ n99 ;
  assign n31 = ~x3 & x6 ;
  assign n32 = x4 & ~n31 ;
  assign n112 = x2 & ~n32 ;
  assign n113 = n112 ^ n101 ;
  assign n114 = n113 ^ n101 ;
  assign n115 = n114 ^ n99 ;
  assign n116 = ~n111 & ~n115 ;
  assign n105 = n101 ^ n31 ;
  assign n106 = n105 ^ n104 ;
  assign n107 = n106 ^ n99 ;
  assign n108 = n104 & n107 ;
  assign n117 = n116 ^ n108 ;
  assign n118 = n117 ^ n104 ;
  assign n119 = n108 ^ n99 ;
  assign n120 = n119 ^ n110 ;
  assign n121 = n99 & ~n120 ;
  assign n122 = n121 ^ n108 ;
  assign n123 = n118 & n122 ;
  assign n124 = n123 ^ n116 ;
  assign n125 = n124 ^ n121 ;
  assign n126 = n125 ^ n104 ;
  assign n127 = n126 ^ n99 ;
  assign n128 = n127 ^ n110 ;
  assign n129 = n128 ^ n100 ;
  assign n130 = ~n95 & n129 ;
  assign n8 = x3 & x5 ;
  assign n9 = ~x3 & ~x6 ;
  assign n10 = ~n8 & ~n9 ;
  assign n11 = x2 & ~x4 ;
  assign n12 = n10 & n11 ;
  assign n16 = ~x2 & ~x4 ;
  assign n13 = x4 & x6 ;
  assign n14 = ~x2 & ~x5 ;
  assign n15 = n13 & n14 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = ~x5 & ~x6 ;
  assign n20 = x1 & n19 ;
  assign n21 = n20 ^ n15 ;
  assign n22 = n21 ^ n15 ;
  assign n23 = n18 & n22 ;
  assign n24 = n23 ^ n15 ;
  assign n25 = ~x3 & n24 ;
  assign n26 = n25 ^ n15 ;
  assign n27 = ~n12 & ~n26 ;
  assign n29 = ~n8 & ~n28 ;
  assign n30 = x6 & ~n29 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = x5 & ~x6 ;
  assign n36 = n35 ^ n30 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = ~n34 & ~n37 ;
  assign n39 = n38 ^ n30 ;
  assign n40 = x2 & ~n39 ;
  assign n41 = n40 ^ n30 ;
  assign n42 = n41 ^ x1 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = x3 ^ x2 ;
  assign n45 = n44 ^ x5 ;
  assign n47 = x5 ^ x3 ;
  assign n48 = n47 ^ x3 ;
  assign n49 = n46 & n48 ;
  assign n50 = n49 ^ x3 ;
  assign n51 = ~n45 & ~n50 ;
  assign n52 = n51 ^ x3 ;
  assign n53 = n52 ^ n41 ;
  assign n54 = ~n43 & ~n53 ;
  assign n55 = n54 ^ n41 ;
  assign n56 = n27 & ~n55 ;
  assign n131 = n130 ^ n56 ;
  assign n132 = n131 ^ n56 ;
  assign n133 = ~x3 & n16 ;
  assign n134 = x6 & n133 ;
  assign n135 = n134 ^ n56 ;
  assign n136 = n135 ^ n56 ;
  assign n137 = n132 & ~n136 ;
  assign n138 = n137 ^ n56 ;
  assign n139 = x0 & n138 ;
  assign n140 = n139 ^ n56 ;
  assign n141 = ~n19 & n133 ;
  assign n142 = n141 ^ x1 ;
  assign n143 = n142 ^ n141 ;
  assign n144 = n143 ^ n140 ;
  assign n145 = ~n13 & ~n96 ;
  assign n146 = x3 & ~n145 ;
  assign n147 = x2 & n28 ;
  assign n148 = n147 ^ n146 ;
  assign n149 = n146 & ~n148 ;
  assign n150 = n149 ^ n141 ;
  assign n151 = n150 ^ n146 ;
  assign n152 = n144 & n151 ;
  assign n153 = n152 ^ n149 ;
  assign n154 = n153 ^ n146 ;
  assign n155 = n140 & n154 ;
  assign n156 = n155 ^ n140 ;
  assign y0 = ~n156 ;
endmodule
