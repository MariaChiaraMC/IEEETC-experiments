module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 ;
  assign n9 = ~x2 & ~x3 ;
  assign n10 = ~x1 & n9 ;
  assign n11 = x5 & ~n10 ;
  assign n12 = n11 ^ x6 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n13 ^ x7 ;
  assign n15 = ~x2 & x3 ;
  assign n16 = x5 & ~n15 ;
  assign n17 = x1 & n16 ;
  assign n18 = n17 ^ x4 ;
  assign n19 = x4 & ~n18 ;
  assign n20 = n19 ^ n11 ;
  assign n21 = n20 ^ x4 ;
  assign n22 = ~n14 & n21 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n23 ^ x4 ;
  assign n25 = x7 & n24 ;
  assign n26 = n25 ^ x7 ;
  assign n27 = ~x0 & ~n26 ;
  assign y0 = n27 ;
endmodule
