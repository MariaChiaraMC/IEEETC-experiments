module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 ;
  assign n12 = x6 ^ x3 ;
  assign n24 = n12 ^ x3 ;
  assign n11 = x3 ^ x2 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n14 ^ x3 ;
  assign n16 = x7 & x8 ;
  assign n17 = ~x6 & n16 ;
  assign n18 = ~x9 & n17 ;
  assign n19 = x1 & ~n18 ;
  assign n20 = n19 ^ n13 ;
  assign n21 = n20 ^ n13 ;
  assign n22 = n21 ^ n15 ;
  assign n23 = n15 & ~n22 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ n15 ;
  assign n27 = x5 ^ x3 ;
  assign n28 = n23 ^ n15 ;
  assign n29 = n27 & n28 ;
  assign n30 = n29 ^ x3 ;
  assign n31 = n26 & ~n30 ;
  assign n32 = n31 ^ x3 ;
  assign n33 = n32 ^ x6 ;
  assign n34 = n33 ^ x3 ;
  assign n35 = ~x4 & n34 ;
  assign n36 = x5 & x9 ;
  assign n37 = n16 & n36 ;
  assign n38 = x3 & ~n37 ;
  assign n39 = ~n35 & ~n38 ;
  assign n40 = ~x0 & ~n39 ;
  assign y0 = n40 ;
endmodule
