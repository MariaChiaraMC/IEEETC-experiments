module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
  assign n13 = x5 & ~x7 ;
  assign n14 = x5 & ~x6 ;
  assign n15 = ~x8 & ~x9 ;
  assign n16 = n14 & n15 ;
  assign n17 = x11 ^ x10 ;
  assign n18 = n16 & n17 ;
  assign n19 = ~n13 & ~n18 ;
  assign n20 = x6 ^ x5 ;
  assign n21 = x7 ^ x6 ;
  assign n22 = n21 ^ x7 ;
  assign n23 = ~x10 & ~x11 ;
  assign n24 = n23 ^ x7 ;
  assign n25 = ~n22 & n24 ;
  assign n26 = n25 ^ x7 ;
  assign n27 = n20 & n26 ;
  assign n28 = x9 ^ x8 ;
  assign n29 = n27 & n28 ;
  assign n30 = n19 & ~n29 ;
  assign n31 = ~x0 & ~x3 ;
  assign n32 = ~x2 & n31 ;
  assign n33 = ~x1 & n32 ;
  assign n34 = ~x4 & n33 ;
  assign n35 = ~n30 & n34 ;
  assign y0 = n35 ;
endmodule
