module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n15 = x2 & x5 ;
  assign n16 = ~x0 & n15 ;
  assign n17 = x4 ^ x3 ;
  assign n18 = n17 ^ x4 ;
  assign n19 = x4 & x8 ;
  assign n20 = ~x11 & n19 ;
  assign n21 = x6 & ~x7 ;
  assign n22 = x1 & ~x9 ;
  assign n23 = n21 & n22 ;
  assign n24 = ~x10 & ~x13 ;
  assign n25 = ~x12 & n24 ;
  assign n26 = n23 & n25 ;
  assign n27 = n20 & n26 ;
  assign n28 = n27 ^ x4 ;
  assign n29 = n18 & ~n28 ;
  assign n30 = n29 ^ x4 ;
  assign n31 = n16 & ~n30 ;
  assign y0 = n31 ;
endmodule
