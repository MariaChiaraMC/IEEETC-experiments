module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 ;
  assign n17 = x6 & x7 ;
  assign n18 = ~x5 & n17 ;
  assign n19 = ~x4 & ~x10 ;
  assign n20 = x0 & n19 ;
  assign n21 = ~x8 & ~x9 ;
  assign n22 = ~x14 & n21 ;
  assign n23 = n20 & n22 ;
  assign n24 = x3 ^ x2 ;
  assign n25 = ~x3 & n24 ;
  assign n26 = x1 & n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = ~x15 & ~n27 ;
  assign n29 = n23 & n28 ;
  assign n30 = n18 & n29 ;
  assign n31 = n30 ^ x13 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = ~x14 & x15 ;
  assign n34 = x3 & x4 ;
  assign n35 = n33 & n34 ;
  assign n36 = x2 & n35 ;
  assign n37 = x5 & x7 ;
  assign n38 = x1 & x9 ;
  assign n39 = ~n37 & n38 ;
  assign n40 = ~x8 & n39 ;
  assign n41 = n36 & n40 ;
  assign n42 = x10 ^ x7 ;
  assign n43 = x6 & n42 ;
  assign n44 = n41 & ~n43 ;
  assign n45 = x2 & ~x14 ;
  assign n46 = ~x9 & n45 ;
  assign n50 = x3 & x10 ;
  assign n47 = ~x7 & ~x10 ;
  assign n48 = ~x3 & x6 ;
  assign n49 = n47 & n48 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = n49 ^ x6 ;
  assign n54 = n53 ^ x7 ;
  assign n55 = n54 ^ n49 ;
  assign n56 = n52 & ~n55 ;
  assign n57 = n56 ^ n49 ;
  assign n58 = x8 & n57 ;
  assign n59 = n58 ^ n49 ;
  assign n60 = n46 & n59 ;
  assign n61 = x4 & ~n60 ;
  assign n62 = ~x1 & ~x15 ;
  assign n63 = x5 ^ x4 ;
  assign n64 = n63 ^ x5 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = ~x6 & x7 ;
  assign n67 = n50 & n66 ;
  assign n72 = ~n49 & ~n67 ;
  assign n73 = n45 & ~n72 ;
  assign n74 = ~x2 & ~x3 ;
  assign n75 = x14 & n74 ;
  assign n76 = n47 & n75 ;
  assign n77 = ~x6 & n76 ;
  assign n78 = ~n73 & ~n77 ;
  assign n79 = n21 & ~n78 ;
  assign n68 = x8 & x9 ;
  assign n80 = x6 & ~x7 ;
  assign n81 = x10 & n80 ;
  assign n82 = n68 & n81 ;
  assign n83 = n75 & n82 ;
  assign n84 = x11 & n83 ;
  assign n85 = ~n79 & ~n84 ;
  assign n69 = ~x2 & ~x14 ;
  assign n70 = n68 & n69 ;
  assign n71 = n67 & n70 ;
  assign n86 = n85 ^ n71 ;
  assign n87 = x5 & n86 ;
  assign n88 = n87 ^ n85 ;
  assign n89 = ~n65 & ~n88 ;
  assign n90 = n89 ^ n87 ;
  assign n91 = n90 ^ n85 ;
  assign n92 = n91 ^ x5 ;
  assign n93 = n62 & ~n92 ;
  assign n94 = ~n61 & n93 ;
  assign n95 = ~n44 & ~n94 ;
  assign n98 = n95 ^ x1 ;
  assign n99 = n98 ^ n95 ;
  assign n96 = n95 ^ n18 ;
  assign n97 = n96 ^ n95 ;
  assign n100 = n99 ^ n97 ;
  assign n101 = ~x2 & n35 ;
  assign n102 = n101 ^ n95 ;
  assign n103 = n102 ^ n95 ;
  assign n104 = n103 ^ n99 ;
  assign n105 = n99 & n104 ;
  assign n106 = n105 ^ n99 ;
  assign n107 = n100 & n106 ;
  assign n108 = n107 ^ n105 ;
  assign n109 = n108 ^ n95 ;
  assign n110 = n109 ^ n99 ;
  assign n111 = x0 & ~n110 ;
  assign n112 = n111 ^ n95 ;
  assign n113 = n112 ^ n30 ;
  assign n114 = ~n32 & ~n113 ;
  assign n115 = n114 ^ n30 ;
  assign n116 = ~x12 & n115 ;
  assign y0 = n116 ;
endmodule
