module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 ;
  assign n10 = ~x0 & x7 ;
  assign n11 = x6 ^ x5 ;
  assign n13 = n11 ^ x4 ;
  assign n14 = n13 ^ x6 ;
  assign n12 = n11 ^ x1 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n15 ^ n11 ;
  assign n17 = n16 ^ n15 ;
  assign n26 = n15 ^ n14 ;
  assign n24 = n15 ^ n13 ;
  assign n18 = n11 ^ x3 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = n19 ^ n14 ;
  assign n21 = n20 ^ n14 ;
  assign n22 = n21 ^ n11 ;
  assign n23 = n22 ^ n16 ;
  assign n25 = n24 ^ n23 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = n17 & ~n27 ;
  assign n29 = n28 ^ n22 ;
  assign n30 = n29 ^ n15 ;
  assign n31 = n20 ^ x2 ;
  assign n32 = n31 ^ n20 ;
  assign n33 = n32 ^ n13 ;
  assign n34 = n33 ^ n15 ;
  assign n35 = n34 ^ n16 ;
  assign n36 = ~n24 & ~n35 ;
  assign n37 = n36 ^ n22 ;
  assign n38 = n37 ^ n33 ;
  assign n39 = n38 ^ n15 ;
  assign n40 = n39 ^ n16 ;
  assign n41 = n40 ^ n26 ;
  assign n42 = n22 ^ n15 ;
  assign n43 = n42 ^ n16 ;
  assign n44 = n43 ^ n26 ;
  assign n45 = n26 ^ n22 ;
  assign n46 = n44 & n45 ;
  assign n47 = n46 ^ n22 ;
  assign n48 = ~n41 & ~n47 ;
  assign n49 = n48 ^ n22 ;
  assign n50 = n49 ^ n16 ;
  assign n51 = ~n30 & ~n50 ;
  assign n52 = n51 ^ n46 ;
  assign n53 = n52 ^ n28 ;
  assign n54 = n53 ^ n48 ;
  assign n55 = n54 ^ n15 ;
  assign n56 = n55 ^ n26 ;
  assign n57 = n56 ^ n11 ;
  assign n58 = n10 & ~n57 ;
  assign y0 = n58 ;
endmodule
