module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 ;
  assign n17 = ~x3 & x13 ;
  assign n18 = x4 & ~x14 ;
  assign n19 = x5 & ~x15 ;
  assign n20 = n18 & n19 ;
  assign n21 = n17 & ~n20 ;
  assign n22 = n21 ^ x0 ;
  assign n23 = x7 & ~x15 ;
  assign n24 = x9 & x10 ;
  assign n25 = ~x8 & ~n24 ;
  assign n26 = x1 & ~x13 ;
  assign n27 = n25 & n26 ;
  assign n28 = n23 & n27 ;
  assign n29 = ~x12 & ~n28 ;
  assign n30 = ~x4 & x14 ;
  assign n31 = ~n18 & ~n30 ;
  assign n32 = x6 ^ x5 ;
  assign n33 = x15 ^ x6 ;
  assign n34 = n32 & n33 ;
  assign n35 = n34 ^ x5 ;
  assign n36 = n31 & ~n35 ;
  assign n37 = x3 & ~n30 ;
  assign n38 = n19 & ~n37 ;
  assign n39 = ~n36 & ~n38 ;
  assign n40 = ~x2 & ~x7 ;
  assign n41 = ~n39 & n40 ;
  assign n42 = n41 ^ x13 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = x4 & ~x7 ;
  assign n45 = n35 & n44 ;
  assign n46 = ~x5 & n30 ;
  assign n47 = ~x2 & ~n18 ;
  assign n48 = ~n46 & n47 ;
  assign n49 = ~x3 & n48 ;
  assign n50 = ~x7 & ~n49 ;
  assign n52 = x5 & x6 ;
  assign n53 = ~x7 & n52 ;
  assign n51 = x14 ^ x12 ;
  assign n54 = n53 ^ n51 ;
  assign n55 = n54 ^ x14 ;
  assign n62 = n55 ^ n54 ;
  assign n56 = n55 ^ x15 ;
  assign n57 = n56 ^ n54 ;
  assign n58 = n54 ^ n53 ;
  assign n59 = n58 ^ x15 ;
  assign n60 = n59 ^ n57 ;
  assign n61 = ~n57 & ~n60 ;
  assign n63 = n62 ^ n61 ;
  assign n64 = n63 ^ n57 ;
  assign n65 = n54 ^ n44 ;
  assign n66 = n61 ^ n57 ;
  assign n67 = ~n65 & ~n66 ;
  assign n68 = n67 ^ n54 ;
  assign n69 = n64 & n68 ;
  assign n70 = n69 ^ n54 ;
  assign n71 = n70 ^ n51 ;
  assign n72 = n71 ^ n54 ;
  assign n73 = ~n50 & ~n72 ;
  assign n74 = ~n45 & n73 ;
  assign n75 = n74 ^ n41 ;
  assign n76 = ~n43 & n75 ;
  assign n77 = n76 ^ n41 ;
  assign n78 = ~n29 & n77 ;
  assign n79 = n78 ^ x11 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = x13 ^ x3 ;
  assign n82 = n19 & n30 ;
  assign n83 = n82 ^ x13 ;
  assign n84 = n83 ^ x13 ;
  assign n85 = ~x5 & x15 ;
  assign n86 = n31 & n85 ;
  assign n87 = n86 ^ x13 ;
  assign n88 = n87 ^ x13 ;
  assign n89 = ~n84 & ~n88 ;
  assign n90 = n89 ^ x13 ;
  assign n91 = ~n81 & n90 ;
  assign n92 = n91 ^ x3 ;
  assign n93 = ~x12 & ~n92 ;
  assign n94 = n93 ^ n78 ;
  assign n95 = n80 & n94 ;
  assign n96 = n95 ^ n78 ;
  assign n97 = n96 ^ n21 ;
  assign n98 = n22 & ~n97 ;
  assign n99 = n98 ^ n95 ;
  assign n100 = n99 ^ n78 ;
  assign n101 = n100 ^ x0 ;
  assign n102 = ~n21 & ~n101 ;
  assign n103 = n102 ^ n21 ;
  assign y0 = ~n103 ;
endmodule
