module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 ;
  assign n11 = ~x1 & ~x2 ;
  assign n64 = x6 & x7 ;
  assign n65 = n11 & n64 ;
  assign n66 = n65 ^ x1 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = ~x6 & ~x7 ;
  assign n69 = n68 ^ n65 ;
  assign n70 = n69 ^ n65 ;
  assign n71 = n67 & n70 ;
  assign n72 = n71 ^ n65 ;
  assign n73 = ~x5 & n72 ;
  assign n74 = n73 ^ n65 ;
  assign n75 = x0 & n74 ;
  assign n76 = x4 & x7 ;
  assign n77 = ~x3 & ~x5 ;
  assign n78 = ~n68 & n77 ;
  assign n79 = ~n76 & n78 ;
  assign n80 = x4 & x5 ;
  assign n33 = ~x4 & ~x5 ;
  assign n81 = n80 ^ n33 ;
  assign n82 = n81 ^ x3 ;
  assign n83 = n33 ^ x6 ;
  assign n84 = n33 ^ x7 ;
  assign n85 = n84 ^ n83 ;
  assign n86 = ~n83 & n85 ;
  assign n87 = n86 ^ n33 ;
  assign n88 = n87 ^ n83 ;
  assign n89 = n82 & ~n88 ;
  assign n90 = n89 ^ n86 ;
  assign n91 = n90 ^ n83 ;
  assign n92 = x3 & ~n91 ;
  assign n93 = x1 & ~n92 ;
  assign n94 = ~n79 & n93 ;
  assign n95 = ~x0 & ~x2 ;
  assign n96 = x6 ^ x1 ;
  assign n97 = n96 ^ n95 ;
  assign n99 = x5 & x7 ;
  assign n98 = ~x3 & ~x4 ;
  assign n100 = n99 ^ n98 ;
  assign n101 = ~x6 & n100 ;
  assign n102 = n101 ^ n98 ;
  assign n103 = ~n97 & ~n102 ;
  assign n104 = n103 ^ n101 ;
  assign n105 = n104 ^ n98 ;
  assign n106 = n105 ^ x6 ;
  assign n107 = n95 & n106 ;
  assign n108 = ~n94 & n107 ;
  assign n109 = ~x1 & x4 ;
  assign n111 = ~x6 & ~n98 ;
  assign n116 = ~x3 & x6 ;
  assign n124 = ~n111 & ~n116 ;
  assign n125 = ~n109 & ~n124 ;
  assign n110 = ~x0 & ~n109 ;
  assign n112 = ~x0 & n77 ;
  assign n113 = n112 ^ x5 ;
  assign n114 = n111 & ~n113 ;
  assign n115 = ~n110 & n114 ;
  assign n117 = ~x0 & x5 ;
  assign n118 = x4 ^ x1 ;
  assign n119 = n117 & ~n118 ;
  assign n120 = n116 & n119 ;
  assign n121 = ~n115 & ~n120 ;
  assign n126 = n125 ^ n121 ;
  assign n127 = n126 ^ n121 ;
  assign n122 = n121 ^ n117 ;
  assign n123 = n122 ^ n121 ;
  assign n128 = n127 ^ n123 ;
  assign n129 = ~x1 & ~n116 ;
  assign n130 = n129 ^ n121 ;
  assign n131 = n130 ^ n121 ;
  assign n132 = n131 ^ n127 ;
  assign n133 = ~n127 & n132 ;
  assign n134 = n133 ^ n127 ;
  assign n135 = ~n128 & ~n134 ;
  assign n136 = n135 ^ n133 ;
  assign n137 = n136 ^ n121 ;
  assign n138 = n137 ^ n127 ;
  assign n139 = x7 & n138 ;
  assign n140 = n139 ^ n121 ;
  assign n141 = x2 & ~n140 ;
  assign n142 = ~n108 & ~n141 ;
  assign n143 = ~n75 & n142 ;
  assign n144 = x8 & ~n143 ;
  assign n12 = ~x7 & n11 ;
  assign n14 = x6 & x8 ;
  assign n13 = ~x6 & ~x8 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = ~x5 & n15 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = n12 & n17 ;
  assign n22 = x5 & n14 ;
  assign n23 = x1 & x7 ;
  assign n24 = n22 & n23 ;
  assign n25 = x4 & n24 ;
  assign n26 = x7 ^ x1 ;
  assign n27 = x5 ^ x4 ;
  assign n28 = n26 & n27 ;
  assign n29 = n17 & n28 ;
  assign n30 = ~n25 & ~n29 ;
  assign n19 = x1 & ~x5 ;
  assign n20 = n15 & ~n19 ;
  assign n21 = n20 ^ n14 ;
  assign n31 = n30 ^ n21 ;
  assign n32 = n31 ^ x2 ;
  assign n42 = n32 ^ n31 ;
  assign n34 = ~x1 & ~x7 ;
  assign n35 = n33 & n34 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ n31 ;
  assign n38 = n35 ^ n21 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n39 ^ n37 ;
  assign n41 = ~n37 & ~n40 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = n43 ^ n37 ;
  assign n45 = x7 ^ x4 ;
  assign n46 = x1 & ~n45 ;
  assign n47 = n46 ^ n31 ;
  assign n48 = n41 ^ n37 ;
  assign n49 = n47 & ~n48 ;
  assign n50 = n49 ^ n31 ;
  assign n51 = ~n44 & ~n50 ;
  assign n52 = n51 ^ n31 ;
  assign n53 = n52 ^ n21 ;
  assign n54 = n53 ^ n31 ;
  assign n55 = ~x3 & n54 ;
  assign n56 = x2 & ~x5 ;
  assign n57 = x3 & ~x4 ;
  assign n58 = n56 & n57 ;
  assign n59 = n13 & n58 ;
  assign n60 = n23 & n59 ;
  assign n61 = ~n55 & ~n60 ;
  assign n62 = ~n18 & n61 ;
  assign n63 = ~x0 & ~n62 ;
  assign n145 = n144 ^ n63 ;
  assign n146 = n145 ^ x9 ;
  assign n153 = n146 ^ n145 ;
  assign n147 = n146 ^ n13 ;
  assign n148 = n147 ^ n145 ;
  assign n149 = n63 ^ n13 ;
  assign n150 = n149 ^ n13 ;
  assign n151 = n150 ^ n148 ;
  assign n152 = n148 & ~n151 ;
  assign n154 = n153 ^ n152 ;
  assign n155 = n154 ^ n148 ;
  assign n156 = ~x2 & n46 ;
  assign n157 = n117 & n156 ;
  assign n158 = ~x0 & ~n118 ;
  assign n159 = n158 ^ n110 ;
  assign n160 = ~x7 & ~n159 ;
  assign n161 = n160 ^ n110 ;
  assign n162 = n56 & ~n161 ;
  assign n163 = ~n157 & ~n162 ;
  assign n164 = x3 & ~n163 ;
  assign n165 = n76 ^ n34 ;
  assign n166 = n34 ^ x2 ;
  assign n167 = n166 ^ n34 ;
  assign n168 = n167 ^ n165 ;
  assign n169 = n165 & n168 ;
  assign n170 = n169 ^ n34 ;
  assign n171 = n170 ^ n165 ;
  assign n172 = n171 ^ x5 ;
  assign n173 = n23 ^ x5 ;
  assign n174 = n98 ^ n34 ;
  assign n175 = n173 & n174 ;
  assign n176 = n175 ^ n98 ;
  assign n177 = n176 ^ n34 ;
  assign n178 = n177 ^ x5 ;
  assign n179 = n34 ^ n23 ;
  assign n180 = ~n23 & ~n179 ;
  assign n181 = n180 ^ x5 ;
  assign n182 = ~n178 & ~n181 ;
  assign n183 = n182 ^ x5 ;
  assign n184 = ~n172 & ~n183 ;
  assign n185 = n184 ^ x5 ;
  assign n186 = x0 & ~n185 ;
  assign n187 = ~n164 & ~n186 ;
  assign n188 = ~n14 & ~n187 ;
  assign n189 = n188 ^ n145 ;
  assign n190 = n152 ^ n148 ;
  assign n191 = n189 & n190 ;
  assign n192 = n191 ^ n145 ;
  assign n193 = ~n155 & n192 ;
  assign n194 = n193 ^ n145 ;
  assign n195 = n194 ^ n63 ;
  assign n196 = n195 ^ n145 ;
  assign y0 = n196 ;
endmodule
