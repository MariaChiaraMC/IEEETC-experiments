module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 ;
  assign n8 = ~x0 & x3 ;
  assign y0 = ~n8 ;
endmodule
