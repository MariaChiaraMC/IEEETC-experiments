// Benchmark "./dk27.pla" written by ABC on Thu Apr 23 10:59:50 2020

module \./dk27.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8,
    z8  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8;
  output z8;
  assign z8 = 1'b1;
endmodule


