module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 ;
  assign n17 = ~x9 & ~x13 ;
  assign n18 = x12 & x14 ;
  assign n19 = n17 & n18 ;
  assign n20 = x15 & n19 ;
  assign n21 = ~x5 & ~n20 ;
  assign n22 = x7 & ~n21 ;
  assign n23 = ~x10 & x11 ;
  assign n24 = x13 & n23 ;
  assign n25 = x10 & ~x11 ;
  assign n26 = ~x13 & n25 ;
  assign n27 = ~n24 & ~n26 ;
  assign n28 = x12 & ~n27 ;
  assign n29 = n28 ^ x14 ;
  assign n30 = n25 ^ n23 ;
  assign n31 = n23 ^ x15 ;
  assign n32 = n31 ^ n23 ;
  assign n33 = n30 & ~n32 ;
  assign n34 = n33 ^ n23 ;
  assign n35 = n34 ^ n28 ;
  assign n36 = ~n29 & ~n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ n23 ;
  assign n39 = n38 ^ x14 ;
  assign n40 = ~n28 & n39 ;
  assign n41 = n40 ^ n28 ;
  assign n42 = n41 ^ n28 ;
  assign n43 = ~x9 & ~n42 ;
  assign n44 = ~x5 & ~x6 ;
  assign n45 = n26 ^ n24 ;
  assign n46 = ~x15 & n45 ;
  assign n47 = n46 ^ n24 ;
  assign n48 = n18 & n47 ;
  assign n49 = ~n44 & ~n48 ;
  assign n50 = ~n43 & n49 ;
  assign n51 = x6 ^ x5 ;
  assign n52 = ~n50 & ~n51 ;
  assign n53 = ~n22 & ~n52 ;
  assign n54 = x4 & ~n53 ;
  assign n56 = x14 & ~x15 ;
  assign n57 = ~x12 & n56 ;
  assign n58 = ~x13 & n57 ;
  assign n59 = ~x7 & ~n58 ;
  assign n60 = ~x6 & ~x9 ;
  assign n61 = ~n59 & n60 ;
  assign n55 = ~x4 & n51 ;
  assign n62 = n61 ^ n55 ;
  assign n63 = n62 ^ x5 ;
  assign n70 = n63 ^ n62 ;
  assign n64 = n63 ^ x7 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = n63 ^ n61 ;
  assign n67 = n66 ^ x7 ;
  assign n68 = n67 ^ n65 ;
  assign n69 = n65 & ~n68 ;
  assign n71 = n70 ^ n69 ;
  assign n72 = n71 ^ n65 ;
  assign n73 = ~x10 & ~x11 ;
  assign n74 = ~x9 & n73 ;
  assign n75 = n74 ^ n62 ;
  assign n76 = n69 ^ n65 ;
  assign n77 = ~n75 & n76 ;
  assign n78 = n77 ^ n62 ;
  assign n79 = n72 & n78 ;
  assign n80 = n79 ^ n62 ;
  assign n81 = n80 ^ n55 ;
  assign n82 = n81 ^ n62 ;
  assign n83 = ~n54 & ~n82 ;
  assign n84 = ~x0 & ~x2 ;
  assign n85 = ~x3 & n84 ;
  assign n86 = x8 & n85 ;
  assign n87 = ~x1 & n86 ;
  assign n88 = ~n83 & n87 ;
  assign y0 = n88 ;
endmodule
