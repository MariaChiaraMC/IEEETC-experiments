// Benchmark "./pla/dc2.pla_res_6NonExact" written by ABC on Fri Nov 20 10:20:13 2020

module \./pla/dc2.pla_res_6NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = x0;
endmodule


