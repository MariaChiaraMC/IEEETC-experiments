module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 ;
  assign n11 = x2 & x3 ;
  assign n12 = x5 ^ x1 ;
  assign n13 = n12 ^ x5 ;
  assign n14 = n13 ^ x4 ;
  assign n15 = ~x8 & ~x9 ;
  assign n16 = n15 ^ x8 ;
  assign n17 = ~x5 & n16 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = ~n14 & n18 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n20 ^ n15 ;
  assign n22 = n21 ^ x5 ;
  assign n23 = x4 & ~n22 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n11 & ~n24 ;
  assign n26 = x3 & ~x4 ;
  assign n27 = n15 ^ x5 ;
  assign n28 = n15 ^ x2 ;
  assign n29 = n15 ^ n12 ;
  assign n30 = n15 & n29 ;
  assign n31 = n30 ^ n15 ;
  assign n32 = ~n28 & n31 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ n15 ;
  assign n35 = n34 ^ n12 ;
  assign n36 = ~n27 & n35 ;
  assign n37 = n36 ^ x5 ;
  assign n38 = n26 & ~n37 ;
  assign n39 = x5 & ~x8 ;
  assign n40 = x3 & ~x5 ;
  assign n41 = ~x2 & n40 ;
  assign n42 = ~n39 & ~n41 ;
  assign n43 = x1 & x4 ;
  assign n44 = ~n42 & n43 ;
  assign n45 = n12 ^ x4 ;
  assign n46 = n45 ^ n12 ;
  assign n47 = ~x1 & x9 ;
  assign n48 = n47 ^ n12 ;
  assign n49 = n48 ^ n12 ;
  assign n50 = ~n46 & n49 ;
  assign n51 = n50 ^ n12 ;
  assign n52 = x3 & ~n51 ;
  assign n53 = n52 ^ n12 ;
  assign n57 = n53 ^ x8 ;
  assign n58 = n57 ^ n53 ;
  assign n54 = x4 & x5 ;
  assign n55 = n54 ^ n53 ;
  assign n56 = n55 ^ n53 ;
  assign n59 = n58 ^ n56 ;
  assign n60 = x3 & x9 ;
  assign n61 = n60 ^ n53 ;
  assign n62 = n61 ^ n53 ;
  assign n63 = n62 ^ n58 ;
  assign n64 = n58 & ~n63 ;
  assign n65 = n64 ^ n58 ;
  assign n66 = n59 & n65 ;
  assign n67 = n66 ^ n64 ;
  assign n68 = n67 ^ n53 ;
  assign n69 = n68 ^ n58 ;
  assign n70 = x2 & ~n69 ;
  assign n71 = n70 ^ n53 ;
  assign n72 = ~n44 & n71 ;
  assign n73 = ~n38 & n72 ;
  assign n74 = ~x0 & ~n73 ;
  assign n75 = x1 & ~x3 ;
  assign n76 = n39 & n75 ;
  assign n77 = ~x2 & n76 ;
  assign n78 = ~n74 & ~n77 ;
  assign n79 = ~n25 & n78 ;
  assign n80 = ~x7 & ~n79 ;
  assign n81 = x2 & x9 ;
  assign n82 = x1 & ~n81 ;
  assign n83 = ~x4 & ~x7 ;
  assign n84 = ~x3 & n83 ;
  assign n85 = ~n82 & n84 ;
  assign n86 = ~x1 & ~x5 ;
  assign n87 = x3 ^ x2 ;
  assign n88 = ~x7 & ~x8 ;
  assign n89 = n88 ^ x4 ;
  assign n90 = x4 ^ x3 ;
  assign n91 = n90 ^ x4 ;
  assign n92 = n89 & ~n91 ;
  assign n93 = n92 ^ x4 ;
  assign n94 = n87 & n93 ;
  assign n95 = n86 & n94 ;
  assign n96 = ~n85 & ~n95 ;
  assign n97 = x0 & ~n96 ;
  assign n98 = ~x3 & x7 ;
  assign n99 = x4 & x8 ;
  assign n100 = ~x3 & ~x5 ;
  assign n101 = n99 & ~n100 ;
  assign n102 = ~n98 & n101 ;
  assign n103 = x3 & x4 ;
  assign n104 = x5 & x9 ;
  assign n105 = n103 & n104 ;
  assign n106 = ~x1 & x5 ;
  assign n107 = ~x3 & x8 ;
  assign n108 = ~n83 & ~n107 ;
  assign n109 = n106 & ~n108 ;
  assign n110 = ~n105 & ~n109 ;
  assign n111 = ~n102 & n110 ;
  assign n112 = n111 ^ x4 ;
  assign n113 = n112 ^ n111 ;
  assign n114 = x5 & x8 ;
  assign n115 = x3 & n114 ;
  assign n116 = ~x5 & ~x8 ;
  assign n117 = ~x1 & n116 ;
  assign n118 = ~n115 & ~n117 ;
  assign n119 = n118 ^ n111 ;
  assign n120 = n119 ^ n111 ;
  assign n121 = ~n113 & ~n120 ;
  assign n122 = n121 ^ n111 ;
  assign n123 = ~x0 & ~n122 ;
  assign n124 = n123 ^ n111 ;
  assign n125 = ~x2 & ~n124 ;
  assign n126 = x0 & ~x5 ;
  assign n127 = x1 & ~x9 ;
  assign n128 = x2 & n127 ;
  assign n129 = x8 ^ x3 ;
  assign n130 = x1 & ~x7 ;
  assign n131 = n130 ^ x8 ;
  assign n132 = n131 ^ n130 ;
  assign n133 = x7 & x9 ;
  assign n134 = n133 ^ n130 ;
  assign n135 = n132 & ~n134 ;
  assign n136 = n135 ^ n130 ;
  assign n137 = n129 & n136 ;
  assign n138 = ~n128 & ~n137 ;
  assign n139 = n138 ^ n11 ;
  assign n140 = n139 ^ x4 ;
  assign n147 = n140 ^ n139 ;
  assign n141 = n140 ^ n130 ;
  assign n142 = n141 ^ n139 ;
  assign n143 = n140 ^ n138 ;
  assign n144 = n143 ^ n130 ;
  assign n145 = n144 ^ n142 ;
  assign n146 = n142 & ~n145 ;
  assign n148 = n147 ^ n146 ;
  assign n149 = n148 ^ n142 ;
  assign n150 = ~x8 & x9 ;
  assign n151 = n150 ^ n139 ;
  assign n152 = n146 ^ n142 ;
  assign n153 = n151 & n152 ;
  assign n154 = n153 ^ n139 ;
  assign n155 = ~n149 & ~n154 ;
  assign n156 = n155 ^ n139 ;
  assign n157 = n156 ^ n11 ;
  assign n158 = n157 ^ n139 ;
  assign n159 = n126 & n158 ;
  assign n160 = ~n125 & ~n159 ;
  assign n161 = ~n97 & n160 ;
  assign n162 = ~n80 & n161 ;
  assign n163 = ~x6 & ~n162 ;
  assign n164 = x8 & x9 ;
  assign n165 = ~x3 & n164 ;
  assign n166 = ~x8 & n11 ;
  assign n167 = ~n165 & ~n166 ;
  assign n168 = n106 & ~n167 ;
  assign n169 = x2 & x8 ;
  assign n170 = x0 & x5 ;
  assign n171 = ~n169 & n170 ;
  assign n172 = ~x0 & ~x5 ;
  assign n173 = x2 & ~x3 ;
  assign n174 = ~n172 & ~n173 ;
  assign n175 = n15 & ~n174 ;
  assign n176 = ~n41 & ~n175 ;
  assign n177 = ~n171 & n176 ;
  assign n178 = x1 & ~n177 ;
  assign n179 = x3 & n106 ;
  assign n180 = ~n173 & ~n179 ;
  assign n181 = ~x0 & ~n180 ;
  assign n182 = ~n178 & ~n181 ;
  assign n183 = ~n168 & n182 ;
  assign n184 = ~x4 & ~n183 ;
  assign n185 = x1 & ~x5 ;
  assign n186 = x4 & ~x9 ;
  assign n187 = ~n185 & ~n186 ;
  assign n188 = ~x2 & ~x8 ;
  assign n189 = x0 & x3 ;
  assign n190 = n188 & n189 ;
  assign n191 = ~n187 & n190 ;
  assign n199 = ~x3 & n126 ;
  assign n194 = x0 & ~x1 ;
  assign n200 = n39 & n194 ;
  assign n201 = ~n199 & ~n200 ;
  assign n202 = ~n115 & n201 ;
  assign n203 = x4 & ~n202 ;
  assign n192 = n116 & n186 ;
  assign n193 = n75 & n192 ;
  assign n195 = ~n164 & ~n194 ;
  assign n196 = ~x3 & x5 ;
  assign n197 = ~n195 & n196 ;
  assign n198 = ~n193 & ~n197 ;
  assign n204 = n203 ^ n198 ;
  assign n205 = n204 ^ n198 ;
  assign n206 = x8 & ~x9 ;
  assign n207 = n179 & n206 ;
  assign n208 = n207 ^ n198 ;
  assign n209 = n208 ^ n198 ;
  assign n210 = ~n205 & ~n209 ;
  assign n211 = n210 ^ n198 ;
  assign n212 = x2 & n211 ;
  assign n213 = n212 ^ n198 ;
  assign n214 = ~n191 & n213 ;
  assign n215 = ~n184 & n214 ;
  assign n216 = x6 & ~n215 ;
  assign n217 = ~x4 & x8 ;
  assign n218 = ~x9 & n170 ;
  assign n219 = n75 & n218 ;
  assign n220 = ~x1 & n81 ;
  assign n221 = n40 & n220 ;
  assign n222 = ~n219 & ~n221 ;
  assign n223 = n217 & ~n222 ;
  assign n224 = ~n103 & ~n114 ;
  assign n225 = ~x1 & x6 ;
  assign n226 = n225 ^ x8 ;
  assign n227 = n226 ^ n225 ;
  assign n228 = n225 ^ n105 ;
  assign n229 = n228 ^ n225 ;
  assign n230 = ~n227 & n229 ;
  assign n231 = n230 ^ n225 ;
  assign n232 = x2 & n231 ;
  assign n233 = n232 ^ n225 ;
  assign n234 = ~n224 & n233 ;
  assign n235 = ~x5 & x8 ;
  assign n236 = x1 & n235 ;
  assign n237 = x4 & n60 ;
  assign n238 = n236 & n237 ;
  assign n239 = x4 & x6 ;
  assign n240 = n100 & ~n127 ;
  assign n241 = ~n164 & n240 ;
  assign n242 = ~n115 & ~n241 ;
  assign n243 = n239 & ~n242 ;
  assign n244 = x1 & x6 ;
  assign n245 = n235 & n244 ;
  assign n246 = x2 & n245 ;
  assign n247 = ~n243 & ~n246 ;
  assign n248 = ~n238 & n247 ;
  assign n249 = ~n234 & n248 ;
  assign n250 = ~x0 & ~n249 ;
  assign n251 = ~n223 & ~n250 ;
  assign n252 = ~n216 & n251 ;
  assign n253 = ~x7 & ~n252 ;
  assign n254 = x5 & x6 ;
  assign n255 = ~x0 & n254 ;
  assign n256 = ~x3 & ~x9 ;
  assign n257 = n256 ^ n47 ;
  assign n258 = n257 ^ n47 ;
  assign n259 = n47 ^ x8 ;
  assign n260 = n259 ^ n47 ;
  assign n261 = n258 & n260 ;
  assign n262 = n261 ^ n47 ;
  assign n263 = ~x4 & n262 ;
  assign n264 = n263 ^ n47 ;
  assign n265 = n255 & n264 ;
  assign n266 = ~x2 & n265 ;
  assign n267 = ~x2 & ~x4 ;
  assign n268 = ~x1 & n199 ;
  assign n269 = n267 & n268 ;
  assign n270 = ~n266 & ~n269 ;
  assign n271 = n103 & n255 ;
  assign n272 = n150 & n271 ;
  assign n273 = n270 & ~n272 ;
  assign n274 = ~n253 & n273 ;
  assign n275 = ~n163 & n274 ;
  assign n276 = ~x0 & x3 ;
  assign n277 = n116 & n276 ;
  assign n278 = ~x4 & n196 ;
  assign n279 = ~n170 & ~n278 ;
  assign n280 = x0 & ~n26 ;
  assign n281 = ~n99 & n280 ;
  assign n282 = ~n279 & ~n281 ;
  assign n283 = ~n277 & ~n282 ;
  assign n284 = n244 & ~n283 ;
  assign n285 = x0 & ~x4 ;
  assign n286 = ~n75 & ~n115 ;
  assign n287 = n285 & ~n286 ;
  assign n288 = ~x0 & ~x4 ;
  assign n289 = n165 & n288 ;
  assign n290 = ~n47 & n116 ;
  assign n291 = n290 ^ x1 ;
  assign n294 = n291 ^ n290 ;
  assign n292 = n291 ^ n54 ;
  assign n293 = n292 ^ n291 ;
  assign n295 = n294 ^ n293 ;
  assign n296 = ~x0 & n114 ;
  assign n297 = n296 ^ n291 ;
  assign n298 = n297 ^ n291 ;
  assign n299 = n298 ^ n293 ;
  assign n300 = ~n293 & n299 ;
  assign n301 = n300 ^ n293 ;
  assign n302 = n295 & ~n301 ;
  assign n303 = n302 ^ n300 ;
  assign n304 = n303 ^ n291 ;
  assign n305 = n304 ^ n293 ;
  assign n306 = ~x3 & n305 ;
  assign n307 = n306 ^ n290 ;
  assign n308 = ~n289 & ~n307 ;
  assign n309 = ~n287 & n308 ;
  assign n310 = ~x6 & ~n309 ;
  assign n324 = ~x4 & ~x5 ;
  assign n325 = ~x0 & ~n324 ;
  assign n326 = n225 & ~n325 ;
  assign n311 = n235 & n276 ;
  assign n312 = x5 ^ x0 ;
  assign n313 = n256 ^ x0 ;
  assign n314 = n256 ^ n244 ;
  assign n315 = n256 & n314 ;
  assign n316 = n315 ^ n256 ;
  assign n317 = n313 & n316 ;
  assign n318 = n317 ^ n315 ;
  assign n319 = n318 ^ n256 ;
  assign n320 = n319 ^ n244 ;
  assign n321 = n312 & n320 ;
  assign n322 = n321 ^ n244 ;
  assign n323 = ~n311 & ~n322 ;
  assign n327 = n326 ^ n323 ;
  assign n328 = n327 ^ x4 ;
  assign n335 = n328 ^ n327 ;
  assign n329 = n328 ^ n40 ;
  assign n330 = n329 ^ n327 ;
  assign n331 = n328 ^ n323 ;
  assign n332 = n331 ^ n40 ;
  assign n333 = n332 ^ n330 ;
  assign n334 = ~n330 & ~n333 ;
  assign n336 = n335 ^ n334 ;
  assign n337 = n336 ^ n330 ;
  assign n338 = n327 ^ n196 ;
  assign n339 = n334 ^ n330 ;
  assign n340 = n338 & ~n339 ;
  assign n341 = n340 ^ n327 ;
  assign n342 = ~n337 & ~n341 ;
  assign n343 = n342 ^ n327 ;
  assign n344 = n343 ^ n326 ;
  assign n345 = n344 ^ n327 ;
  assign n346 = ~n310 & ~n345 ;
  assign n347 = x7 & ~n346 ;
  assign n348 = x4 & n116 ;
  assign n349 = x0 & n348 ;
  assign n350 = ~n114 & n288 ;
  assign n351 = ~n164 & n350 ;
  assign n352 = ~n349 & ~n351 ;
  assign n353 = x6 & ~n352 ;
  assign n356 = n353 ^ n54 ;
  assign n357 = n356 ^ n353 ;
  assign n354 = n353 ^ x0 ;
  assign n355 = n354 ^ n353 ;
  assign n358 = n357 ^ n355 ;
  assign n359 = n353 ^ x1 ;
  assign n360 = n359 ^ n353 ;
  assign n361 = n360 ^ n357 ;
  assign n362 = n357 & n361 ;
  assign n363 = n362 ^ n357 ;
  assign n364 = ~n358 & n363 ;
  assign n365 = n364 ^ n362 ;
  assign n366 = n365 ^ n353 ;
  assign n367 = n366 ^ n357 ;
  assign n368 = x3 & n367 ;
  assign n369 = n368 ^ n353 ;
  assign n370 = ~n347 & ~n369 ;
  assign n371 = ~n284 & n370 ;
  assign n372 = x2 & ~n371 ;
  assign n381 = n235 & n285 ;
  assign n373 = n99 ^ x5 ;
  assign n374 = n373 ^ n99 ;
  assign n375 = x4 & n164 ;
  assign n376 = ~n188 & ~n375 ;
  assign n377 = n376 ^ n99 ;
  assign n378 = n374 & ~n377 ;
  assign n379 = n378 ^ n99 ;
  assign n380 = ~n312 & n379 ;
  assign n382 = n381 ^ n380 ;
  assign n383 = x6 & n382 ;
  assign n384 = n383 ^ n380 ;
  assign n385 = ~x1 & n384 ;
  assign n386 = n385 ^ x7 ;
  assign n387 = x8 & n47 ;
  assign n388 = ~x0 & ~n387 ;
  assign n389 = n324 ^ x4 ;
  assign n390 = n389 ^ x4 ;
  assign n391 = x8 ^ x4 ;
  assign n392 = n391 ^ x4 ;
  assign n393 = n390 & ~n392 ;
  assign n394 = n393 ^ x4 ;
  assign n395 = x6 & n394 ;
  assign n396 = n395 ^ x4 ;
  assign n397 = ~n388 & n396 ;
  assign n398 = ~x0 & x6 ;
  assign n399 = n186 & n398 ;
  assign n400 = ~x4 & ~x6 ;
  assign n401 = n400 ^ x0 ;
  assign n402 = n400 ^ n206 ;
  assign n403 = n402 ^ n206 ;
  assign n404 = n403 ^ n401 ;
  assign n405 = n244 ^ x8 ;
  assign n406 = n244 & n405 ;
  assign n407 = n406 ^ n206 ;
  assign n408 = n407 ^ n244 ;
  assign n409 = n404 & ~n408 ;
  assign n410 = n409 ^ n406 ;
  assign n411 = n410 ^ n244 ;
  assign n412 = ~n401 & n411 ;
  assign n413 = n412 ^ n400 ;
  assign n414 = x5 & n413 ;
  assign n415 = ~n399 & ~n414 ;
  assign n416 = ~n397 & n415 ;
  assign n417 = ~x2 & ~n416 ;
  assign n418 = ~x1 & ~n39 ;
  assign n419 = n239 & ~n418 ;
  assign n420 = n400 ^ n47 ;
  assign n421 = n420 ^ n236 ;
  assign n422 = n421 ^ n400 ;
  assign n423 = n422 ^ n421 ;
  assign n424 = n421 ^ n348 ;
  assign n425 = n424 ^ n420 ;
  assign n426 = n423 & ~n425 ;
  assign n427 = n426 ^ n348 ;
  assign n428 = ~n114 & ~n348 ;
  assign n429 = n428 ^ n420 ;
  assign n430 = ~n427 & ~n429 ;
  assign n431 = n430 ^ n428 ;
  assign n432 = ~n420 & n431 ;
  assign n433 = n432 ^ n426 ;
  assign n434 = n433 ^ n47 ;
  assign n435 = n434 ^ n348 ;
  assign n436 = ~n419 & n435 ;
  assign n437 = ~x0 & ~n436 ;
  assign n438 = n104 & n285 ;
  assign n439 = ~n192 & ~n438 ;
  assign n440 = x1 & ~x6 ;
  assign n441 = ~n439 & n440 ;
  assign n442 = ~n437 & ~n441 ;
  assign n443 = ~n417 & n442 ;
  assign n444 = n443 ^ x3 ;
  assign n445 = n444 ^ n443 ;
  assign n446 = ~x0 & x8 ;
  assign n447 = ~x5 & ~x6 ;
  assign n448 = n446 & n447 ;
  assign n449 = ~n254 & ~n448 ;
  assign n450 = ~x2 & ~n449 ;
  assign n451 = x8 & n255 ;
  assign n452 = x6 & n164 ;
  assign n453 = ~x0 & ~x6 ;
  assign n454 = ~n452 & ~n453 ;
  assign n455 = x6 ^ x5 ;
  assign n456 = ~n454 & ~n455 ;
  assign n457 = ~n451 & ~n456 ;
  assign n458 = ~x1 & ~n457 ;
  assign n459 = ~n450 & ~n458 ;
  assign n460 = x4 & ~n459 ;
  assign n461 = n106 & n398 ;
  assign n462 = n150 & n453 ;
  assign n463 = n462 ^ x1 ;
  assign n464 = n463 ^ x5 ;
  assign n471 = n464 ^ n463 ;
  assign n466 = n324 & ~n454 ;
  assign n465 = n464 ^ n462 ;
  assign n467 = n466 ^ n465 ;
  assign n468 = n466 ^ n464 ;
  assign n469 = n468 ^ n463 ;
  assign n470 = ~n467 & n469 ;
  assign n472 = n471 ^ n470 ;
  assign n473 = ~x6 & ~n186 ;
  assign n474 = ~x8 & ~n473 ;
  assign n475 = n474 ^ n464 ;
  assign n476 = ~n471 & ~n475 ;
  assign n477 = n476 ^ n474 ;
  assign n478 = ~n472 & n477 ;
  assign n479 = n478 ^ n470 ;
  assign n480 = n479 ^ n464 ;
  assign n481 = n480 ^ x1 ;
  assign n482 = n481 ^ n463 ;
  assign n483 = ~n461 & n482 ;
  assign n484 = ~x2 & ~n483 ;
  assign n485 = x4 & ~x6 ;
  assign n486 = ~x2 & n452 ;
  assign n487 = ~n485 & ~n486 ;
  assign n488 = x1 & ~n487 ;
  assign n489 = ~x8 & n400 ;
  assign n490 = x9 ^ x8 ;
  assign n491 = n267 & n490 ;
  assign n492 = ~n489 & ~n491 ;
  assign n493 = ~n488 & n492 ;
  assign n494 = n126 & ~n493 ;
  assign n495 = n15 & n106 ;
  assign n496 = n285 & n495 ;
  assign n497 = ~n494 & ~n496 ;
  assign n498 = ~n484 & n497 ;
  assign n499 = ~n460 & n498 ;
  assign n500 = n499 ^ n443 ;
  assign n501 = ~n445 & n500 ;
  assign n502 = n501 ^ n443 ;
  assign n503 = n502 ^ n385 ;
  assign n504 = ~n386 & ~n503 ;
  assign n505 = n504 ^ n501 ;
  assign n506 = n505 ^ n443 ;
  assign n507 = n506 ^ x7 ;
  assign n508 = ~n385 & n507 ;
  assign n509 = n508 ^ n385 ;
  assign n510 = n509 ^ x7 ;
  assign n511 = ~n372 & n510 ;
  assign n512 = n275 & n511 ;
  assign y0 = ~n512 ;
endmodule
