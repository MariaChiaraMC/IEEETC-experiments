module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 ;
  assign n7 = ~x2 & ~x5 ;
  assign n8 = ~x3 & n7 ;
  assign n9 = x1 & ~n8 ;
  assign n10 = x0 & ~n9 ;
  assign n11 = x3 ^ x2 ;
  assign n12 = n11 ^ x4 ;
  assign n13 = n12 ^ x1 ;
  assign n14 = x5 ^ x4 ;
  assign n15 = n14 ^ x4 ;
  assign n16 = x4 ^ x3 ;
  assign n17 = n16 ^ x4 ;
  assign n18 = n15 & ~n17 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = n19 ^ n12 ;
  assign n21 = n13 & n20 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = n22 ^ x4 ;
  assign n24 = n23 ^ x1 ;
  assign n25 = ~n12 & n24 ;
  assign n26 = n25 ^ n12 ;
  assign n27 = n10 & n26 ;
  assign y0 = n27 ;
endmodule
