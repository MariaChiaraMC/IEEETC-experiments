module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n10 = x5 ^ x3 ;
  assign n11 = n10 ^ x3 ;
  assign n12 = n11 ^ x4 ;
  assign n13 = x2 ^ x0 ;
  assign n14 = ~x0 & n13 ;
  assign n15 = n14 ^ x3 ;
  assign n16 = n15 ^ x0 ;
  assign n17 = n12 & ~n16 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = n18 ^ x0 ;
  assign n20 = x4 & ~n19 ;
  assign n21 = n20 ^ x4 ;
  assign n22 = x6 & ~n21 ;
  assign n23 = ~x2 & x5 ;
  assign n24 = x3 & n23 ;
  assign n25 = ~x4 & ~n24 ;
  assign n26 = x1 & ~n25 ;
  assign n27 = ~x0 & n26 ;
  assign n28 = n22 & ~n27 ;
  assign y0 = n28 ;
endmodule
