module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 ;
  assign n15 = x2 & ~x3 ;
  assign n16 = ~x1 & n15 ;
  assign n17 = x0 & n16 ;
  assign n18 = ~x4 & n15 ;
  assign n19 = x7 & x8 ;
  assign n20 = ~x11 & ~n19 ;
  assign n21 = x6 & ~n20 ;
  assign n22 = ~x12 & ~x13 ;
  assign n23 = ~x6 & ~x11 ;
  assign n24 = ~n22 & ~n23 ;
  assign n25 = ~x10 & ~n24 ;
  assign n26 = ~x12 & x13 ;
  assign n27 = ~x11 & ~n26 ;
  assign n28 = ~x6 & n22 ;
  assign n29 = n28 ^ x13 ;
  assign n30 = n27 & n29 ;
  assign n31 = x8 & ~x9 ;
  assign n32 = x7 & ~x9 ;
  assign n33 = ~n31 & ~n32 ;
  assign n34 = ~n30 & ~n33 ;
  assign n35 = n25 & n34 ;
  assign n36 = ~n21 & n35 ;
  assign n37 = ~x5 & ~n36 ;
  assign n38 = n18 & ~n37 ;
  assign n39 = n38 ^ x1 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = n40 ^ x0 ;
  assign n42 = x6 & ~x7 ;
  assign n43 = ~x3 & n42 ;
  assign n44 = ~x2 & x5 ;
  assign n45 = x4 & n44 ;
  assign n46 = n43 & n45 ;
  assign n47 = ~x8 & ~x9 ;
  assign n48 = ~x6 & x7 ;
  assign n49 = ~n42 & ~n48 ;
  assign n50 = n47 & ~n49 ;
  assign n51 = x5 & ~n50 ;
  assign n52 = n15 & ~n51 ;
  assign n53 = ~n18 & ~n52 ;
  assign n54 = x5 ^ x2 ;
  assign n55 = n54 ^ x3 ;
  assign n65 = x9 ^ x8 ;
  assign n56 = x8 ^ x4 ;
  assign n57 = n56 ^ x9 ;
  assign n58 = n57 ^ x9 ;
  assign n59 = n58 ^ x8 ;
  assign n60 = n57 ^ x7 ;
  assign n61 = n60 ^ x6 ;
  assign n62 = n61 ^ n57 ;
  assign n63 = n62 ^ n59 ;
  assign n64 = ~n59 & n63 ;
  assign n66 = n65 ^ n64 ;
  assign n67 = n66 ^ n59 ;
  assign n68 = x8 ^ x6 ;
  assign n69 = n64 ^ n59 ;
  assign n70 = n68 & ~n69 ;
  assign n71 = n70 ^ x8 ;
  assign n72 = n67 & ~n71 ;
  assign n73 = n72 ^ x8 ;
  assign n74 = n73 ^ x8 ;
  assign n75 = n74 ^ x5 ;
  assign n76 = n75 ^ n74 ;
  assign n77 = x4 & x12 ;
  assign n78 = n31 ^ x13 ;
  assign n79 = n78 ^ n31 ;
  assign n80 = ~x8 & x9 ;
  assign n81 = n80 ^ n31 ;
  assign n82 = n79 & n81 ;
  assign n83 = n82 ^ n31 ;
  assign n84 = n77 & n83 ;
  assign n85 = n84 ^ n74 ;
  assign n86 = ~n76 & n85 ;
  assign n87 = n86 ^ n74 ;
  assign n88 = n87 ^ n54 ;
  assign n89 = n55 & ~n88 ;
  assign n90 = n89 ^ n86 ;
  assign n91 = n90 ^ n74 ;
  assign n92 = n91 ^ x3 ;
  assign n93 = n54 & ~n92 ;
  assign n94 = n93 ^ n54 ;
  assign n95 = n94 ^ x3 ;
  assign n96 = n53 & ~n95 ;
  assign n97 = ~x10 & ~n27 ;
  assign n98 = ~n96 & n97 ;
  assign n99 = ~n46 & ~n98 ;
  assign n100 = ~x4 & ~x6 ;
  assign n101 = ~n31 & ~n80 ;
  assign n102 = n100 & ~n101 ;
  assign n103 = ~x7 & n102 ;
  assign n104 = x4 & n47 ;
  assign n105 = ~x2 & ~n104 ;
  assign n106 = ~n103 & n105 ;
  assign n107 = x2 & ~x5 ;
  assign n108 = x11 & n81 ;
  assign n109 = n108 ^ n31 ;
  assign n110 = x4 & n109 ;
  assign n111 = n107 & ~n110 ;
  assign n112 = x3 & ~n111 ;
  assign n113 = ~n106 & n112 ;
  assign n114 = x3 ^ x2 ;
  assign n115 = ~n51 & n114 ;
  assign n116 = ~n18 & n115 ;
  assign n117 = n116 ^ n18 ;
  assign n118 = ~n113 & ~n117 ;
  assign n119 = x10 & ~n118 ;
  assign n120 = n26 & n119 ;
  assign n121 = n120 ^ n99 ;
  assign n122 = n99 & ~n121 ;
  assign n123 = n122 ^ n38 ;
  assign n124 = n123 ^ n99 ;
  assign n125 = n41 & ~n124 ;
  assign n126 = n125 ^ n122 ;
  assign n127 = n126 ^ n99 ;
  assign n128 = ~x0 & n127 ;
  assign n129 = n128 ^ x0 ;
  assign n130 = ~n17 & n129 ;
  assign y0 = ~n130 ;
endmodule
