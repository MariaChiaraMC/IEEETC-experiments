module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 ;
  assign n10 = x6 ^ x5 ;
  assign n9 = x7 ^ x2 ;
  assign n15 = n10 ^ n9 ;
  assign n16 = n15 ^ x4 ;
  assign n17 = n16 ^ x4 ;
  assign n18 = x7 ^ x6 ;
  assign n19 = n18 ^ n10 ;
  assign n20 = n19 ^ x4 ;
  assign n21 = n17 & ~n20 ;
  assign n11 = n10 ^ x7 ;
  assign n12 = n11 ^ n9 ;
  assign n13 = n12 ^ x4 ;
  assign n14 = n9 & n13 ;
  assign n22 = n21 ^ n14 ;
  assign n23 = n22 ^ n9 ;
  assign n24 = n14 ^ x4 ;
  assign n25 = n24 ^ n16 ;
  assign n26 = x4 & n25 ;
  assign n27 = n26 ^ n14 ;
  assign n28 = n23 & n27 ;
  assign n29 = n28 ^ n21 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n30 ^ n9 ;
  assign n32 = n31 ^ x4 ;
  assign n33 = n32 ^ n16 ;
  assign n34 = ~x3 & n33 ;
  assign n35 = x6 ^ x4 ;
  assign n36 = x6 ^ x3 ;
  assign n37 = ~x2 & ~x5 ;
  assign n38 = ~x7 & n37 ;
  assign n39 = n38 ^ x3 ;
  assign n40 = ~x3 & ~n39 ;
  assign n41 = n40 ^ x3 ;
  assign n42 = n36 & ~n41 ;
  assign n43 = n42 ^ n40 ;
  assign n44 = n43 ^ x3 ;
  assign n45 = n44 ^ n38 ;
  assign n46 = ~n35 & ~n45 ;
  assign n47 = ~n34 & ~n46 ;
  assign n48 = ~x0 & ~x1 ;
  assign n49 = ~n47 & n48 ;
  assign y0 = n49 ;
endmodule
