module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n9 = x3 ^ x2 ;
  assign n10 = n9 ^ x3 ;
  assign n11 = n10 ^ x0 ;
  assign n12 = x5 ^ x4 ;
  assign n13 = n12 ^ x6 ;
  assign n14 = n13 ^ x1 ;
  assign n15 = x7 ^ x6 ;
  assign n16 = x6 ^ x5 ;
  assign n17 = n16 ^ x6 ;
  assign n18 = ~n15 & n17 ;
  assign n19 = n18 ^ x6 ;
  assign n20 = n19 ^ n13 ;
  assign n21 = ~n14 & n20 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = n22 ^ x6 ;
  assign n24 = n23 ^ x1 ;
  assign n25 = n13 & ~n24 ;
  assign n26 = n25 ^ n13 ;
  assign n27 = n26 ^ x1 ;
  assign n28 = ~x3 & ~n27 ;
  assign n29 = n28 ^ x1 ;
  assign n30 = n11 & n29 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n31 ^ x1 ;
  assign n33 = n32 ^ x3 ;
  assign n34 = ~x0 & ~n33 ;
  assign y0 = n34 ;
endmodule
