module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 ;
  assign n8 = x3 & x6 ;
  assign n9 = n8 ^ x5 ;
  assign n10 = x0 & ~n9 ;
  assign n11 = n10 ^ x5 ;
  assign n12 = n11 ^ x2 ;
  assign n20 = n12 ^ n11 ;
  assign n21 = n20 ^ x3 ;
  assign n22 = n21 ^ x3 ;
  assign n23 = n12 ^ x5 ;
  assign n24 = n23 ^ x3 ;
  assign n25 = n22 & ~n24 ;
  assign n13 = x4 & x6 ;
  assign n14 = x0 & n13 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = n16 ^ n11 ;
  assign n18 = n17 ^ x3 ;
  assign n19 = n11 & n18 ;
  assign n26 = n25 ^ n19 ;
  assign n27 = n26 ^ n11 ;
  assign n28 = n19 ^ x3 ;
  assign n29 = n28 ^ n21 ;
  assign n30 = ~x3 & n29 ;
  assign n31 = n30 ^ n19 ;
  assign n32 = n27 & n31 ;
  assign n33 = n32 ^ n25 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ n11 ;
  assign n36 = n35 ^ x3 ;
  assign n37 = n36 ^ n21 ;
  assign n38 = n37 ^ x2 ;
  assign n39 = ~x1 & n38 ;
  assign n40 = ~x4 & x6 ;
  assign n41 = x2 & n40 ;
  assign n42 = ~x3 & ~n41 ;
  assign n43 = n42 ^ x2 ;
  assign n44 = n42 ^ x1 ;
  assign n45 = n44 ^ n42 ;
  assign n46 = n45 ^ n43 ;
  assign n47 = ~x5 & ~x6 ;
  assign n48 = n47 ^ n8 ;
  assign n49 = ~n42 & ~n48 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = n46 & ~n50 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = n52 ^ n47 ;
  assign n54 = n53 ^ n42 ;
  assign n55 = n43 & n54 ;
  assign n56 = n55 ^ x2 ;
  assign n57 = ~x0 & n56 ;
  assign n58 = ~n39 & ~n57 ;
  assign y0 = ~n58 ;
endmodule
