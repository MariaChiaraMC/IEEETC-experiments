module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 ;
  assign n22 = x1 ^ x0 ;
  assign n23 = x2 ^ x1 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = x5 ^ x3 ;
  assign n27 = x5 ^ x1 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = ~n26 & ~n28 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = n30 ^ n26 ;
  assign n32 = n25 & ~n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ n26 ;
  assign n35 = n22 & ~n34 ;
  assign n36 = ~x4 & n35 ;
  assign n37 = x14 & ~n36 ;
  assign n215 = ~x19 & ~x20 ;
  assign n38 = ~x12 & ~x13 ;
  assign n39 = x8 & x9 ;
  assign n40 = ~x0 & ~x2 ;
  assign n41 = x1 & n40 ;
  assign n42 = ~x6 & ~x7 ;
  assign n43 = ~x10 & x11 ;
  assign n44 = ~x4 & n43 ;
  assign n45 = n42 & n44 ;
  assign n46 = n41 & n45 ;
  assign n47 = ~x1 & x3 ;
  assign n48 = n45 ^ x0 ;
  assign n49 = n48 ^ x2 ;
  assign n58 = n49 ^ n48 ;
  assign n50 = n42 & n43 ;
  assign n51 = ~x5 & n50 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = n52 ^ n48 ;
  assign n54 = n49 ^ n45 ;
  assign n55 = n54 ^ n51 ;
  assign n56 = n55 ^ n53 ;
  assign n57 = ~n53 & ~n56 ;
  assign n59 = n58 ^ n57 ;
  assign n60 = n59 ^ n53 ;
  assign n61 = x10 & ~x11 ;
  assign n62 = n61 ^ n48 ;
  assign n63 = n57 ^ n53 ;
  assign n64 = ~n62 & ~n63 ;
  assign n65 = n64 ^ n48 ;
  assign n66 = ~n60 & n65 ;
  assign n67 = n66 ^ n48 ;
  assign n68 = n67 ^ x0 ;
  assign n69 = n68 ^ n48 ;
  assign n70 = n47 & n69 ;
  assign n71 = ~n46 & ~n70 ;
  assign n72 = n39 & ~n71 ;
  assign n73 = x2 & x5 ;
  assign n74 = ~n40 & ~n73 ;
  assign n75 = x9 & ~n74 ;
  assign n76 = ~x11 & n75 ;
  assign n77 = x5 & ~x9 ;
  assign n78 = ~x1 & ~x2 ;
  assign n79 = ~x0 & n78 ;
  assign n80 = ~n77 & ~n79 ;
  assign n81 = n61 & ~n80 ;
  assign n82 = ~n76 & ~n81 ;
  assign n83 = ~x8 & n42 ;
  assign n84 = ~x4 & n83 ;
  assign n85 = ~n82 & n84 ;
  assign n86 = ~n72 & ~n85 ;
  assign n87 = n38 & ~n86 ;
  assign n88 = x5 & ~x8 ;
  assign n89 = x13 & n88 ;
  assign n90 = ~x9 & n43 ;
  assign n91 = ~x4 & n90 ;
  assign n92 = n89 & n91 ;
  assign n93 = ~x0 & x4 ;
  assign n94 = ~x5 & ~n93 ;
  assign n95 = x2 & ~n94 ;
  assign n96 = x1 & n95 ;
  assign n97 = ~n92 & ~n96 ;
  assign n98 = ~x8 & ~x9 ;
  assign n99 = x5 & ~x12 ;
  assign n100 = n45 & n99 ;
  assign n101 = n98 & n100 ;
  assign n102 = n97 & ~n101 ;
  assign n103 = n78 ^ x5 ;
  assign n104 = n103 ^ n78 ;
  assign n105 = ~x0 & ~x1 ;
  assign n106 = x4 & ~n105 ;
  assign n107 = n106 ^ n78 ;
  assign n108 = ~n104 & n107 ;
  assign n109 = n108 ^ n78 ;
  assign n110 = x3 & n109 ;
  assign n111 = n102 & ~n110 ;
  assign n112 = ~x0 & ~x4 ;
  assign n113 = x1 & n112 ;
  assign n114 = n38 & n113 ;
  assign n115 = n42 ^ x10 ;
  assign n116 = ~x8 & n115 ;
  assign n117 = n116 ^ x10 ;
  assign n118 = n114 & n117 ;
  assign n119 = n118 ^ x11 ;
  assign n120 = n119 ^ n118 ;
  assign n121 = x12 ^ x5 ;
  assign n122 = n121 ^ n118 ;
  assign n123 = ~n120 & n122 ;
  assign n124 = n123 ^ x12 ;
  assign n125 = n124 ^ x5 ;
  assign n126 = n125 ^ n120 ;
  assign n127 = n119 ^ x10 ;
  assign n128 = n127 ^ n118 ;
  assign n129 = n128 ^ n126 ;
  assign n130 = n128 ^ n120 ;
  assign n131 = n89 ^ x12 ;
  assign n132 = ~n130 & ~n131 ;
  assign n133 = n132 ^ x12 ;
  assign n134 = ~n129 & ~n133 ;
  assign n135 = n134 ^ n120 ;
  assign n136 = ~n126 & ~n135 ;
  assign n137 = n136 ^ x11 ;
  assign n138 = x9 & ~n137 ;
  assign n139 = x0 & ~x13 ;
  assign n140 = x1 & ~n139 ;
  assign n141 = x4 & ~n140 ;
  assign n142 = x5 & ~n141 ;
  assign n143 = x11 & ~x12 ;
  assign n144 = ~x1 & x9 ;
  assign n145 = n143 & n144 ;
  assign n146 = n88 & n145 ;
  assign n147 = ~n142 & ~n146 ;
  assign n148 = x0 & ~x1 ;
  assign n149 = x4 & n148 ;
  assign n150 = n149 ^ n147 ;
  assign n151 = x13 & n99 ;
  assign n152 = ~n112 & ~n151 ;
  assign n153 = n152 ^ x2 ;
  assign n154 = n153 ^ n152 ;
  assign n155 = ~x8 & n148 ;
  assign n156 = n90 & n155 ;
  assign n157 = x13 ^ x5 ;
  assign n158 = x1 & n98 ;
  assign n159 = ~x4 & n158 ;
  assign n160 = ~n155 & ~n159 ;
  assign n161 = n61 & ~n160 ;
  assign n162 = n39 & n44 ;
  assign n163 = ~n105 & n162 ;
  assign n164 = ~n161 & ~n163 ;
  assign n165 = n42 & ~n164 ;
  assign n166 = ~x12 & n165 ;
  assign n167 = n166 ^ n157 ;
  assign n168 = n167 ^ x13 ;
  assign n169 = n168 ^ n167 ;
  assign n170 = ~x6 & ~x10 ;
  assign n171 = ~x17 & n170 ;
  assign n172 = x13 & x15 ;
  assign n173 = n171 & ~n172 ;
  assign n174 = n173 ^ n98 ;
  assign n175 = ~x7 & x16 ;
  assign n176 = n175 ^ x11 ;
  assign n177 = n176 ^ n175 ;
  assign n178 = n175 ^ x12 ;
  assign n179 = ~n177 & ~n178 ;
  assign n180 = n179 ^ n175 ;
  assign n181 = n180 ^ n173 ;
  assign n182 = n174 & n181 ;
  assign n183 = n182 ^ n179 ;
  assign n184 = n183 ^ n175 ;
  assign n185 = n184 ^ n98 ;
  assign n186 = n173 & n185 ;
  assign n187 = n186 ^ n173 ;
  assign n188 = n187 ^ n167 ;
  assign n189 = n188 ^ n157 ;
  assign n190 = ~n169 & n189 ;
  assign n191 = n190 ^ n187 ;
  assign n192 = n143 & n187 ;
  assign n193 = n192 ^ n157 ;
  assign n194 = n191 & n193 ;
  assign n195 = n194 ^ n192 ;
  assign n196 = n157 & n195 ;
  assign n197 = n196 ^ n190 ;
  assign n198 = n197 ^ x5 ;
  assign n199 = n198 ^ n187 ;
  assign n200 = ~n156 & ~n199 ;
  assign n201 = n200 ^ n152 ;
  assign n202 = n154 & n201 ;
  assign n203 = n202 ^ n152 ;
  assign n204 = n203 ^ n147 ;
  assign n205 = ~n150 & n204 ;
  assign n206 = n205 ^ n202 ;
  assign n207 = n206 ^ n152 ;
  assign n208 = n207 ^ n149 ;
  assign n209 = n147 & ~n208 ;
  assign n210 = n209 ^ n147 ;
  assign n211 = ~n138 & n210 ;
  assign n212 = ~x3 & ~n211 ;
  assign n213 = n111 & ~n212 ;
  assign n214 = ~n87 & n213 ;
  assign n216 = n215 ^ n214 ;
  assign n217 = n216 ^ n214 ;
  assign n218 = n214 ^ x18 ;
  assign n219 = ~n217 & n218 ;
  assign n220 = n219 ^ n214 ;
  assign n221 = n37 & n220 ;
  assign y0 = ~n221 ;
endmodule
