module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 ;
  assign n9 = ~x1 & x2 ;
  assign n10 = ~x5 & ~x6 ;
  assign n11 = x7 ^ x4 ;
  assign n12 = n11 ^ x4 ;
  assign n13 = n12 ^ n10 ;
  assign n14 = x3 ^ x0 ;
  assign n15 = x4 & ~n14 ;
  assign n16 = n15 ^ x3 ;
  assign n17 = ~n13 & ~n16 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n18 ^ x3 ;
  assign n20 = n19 ^ x4 ;
  assign n21 = n10 & ~n20 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = n9 & ~n22 ;
  assign n24 = x7 ^ x3 ;
  assign n25 = n24 ^ n14 ;
  assign n26 = x7 ^ x5 ;
  assign n27 = n26 ^ x5 ;
  assign n28 = x5 & x6 ;
  assign n29 = n28 ^ x5 ;
  assign n30 = n27 & ~n29 ;
  assign n31 = n30 ^ x5 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = ~n25 & ~n32 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ x5 ;
  assign n36 = n35 ^ n14 ;
  assign n37 = n24 & n36 ;
  assign n38 = n37 ^ n24 ;
  assign n39 = n38 ^ x3 ;
  assign n40 = n23 & ~n39 ;
  assign y0 = n40 ;
endmodule
