module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 ;
  assign n16 = ~x11 & ~x12 ;
  assign n17 = ~x2 & x3 ;
  assign n18 = ~x4 & ~n17 ;
  assign n19 = x8 & x9 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = n19 ^ x9 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = ~n21 & ~n23 ;
  assign n25 = n24 ^ n19 ;
  assign n26 = x7 & n25 ;
  assign n27 = n26 ^ n19 ;
  assign n28 = x6 & n27 ;
  assign n29 = n18 & n28 ;
  assign n30 = x1 & ~n29 ;
  assign n31 = x2 & x3 ;
  assign n32 = ~x0 & ~x13 ;
  assign n33 = n31 & n32 ;
  assign n34 = x7 & n33 ;
  assign n35 = x10 & ~n34 ;
  assign n36 = ~x14 & ~n35 ;
  assign n37 = ~n30 & n36 ;
  assign n38 = ~x2 & ~x7 ;
  assign n39 = ~x3 & x13 ;
  assign n40 = n38 & n39 ;
  assign n41 = ~x9 & n40 ;
  assign n42 = ~x10 & ~n41 ;
  assign n43 = ~x6 & ~x8 ;
  assign n44 = ~n42 & n43 ;
  assign n45 = ~x4 & n44 ;
  assign n46 = n45 ^ x13 ;
  assign n49 = n46 ^ n45 ;
  assign n47 = n46 ^ x1 ;
  assign n48 = n47 ^ n46 ;
  assign n50 = n49 ^ n48 ;
  assign n51 = x4 & x7 ;
  assign n52 = x6 & n51 ;
  assign n53 = x9 ^ x8 ;
  assign n54 = n52 & ~n53 ;
  assign n55 = n31 & n54 ;
  assign n56 = n55 ^ n46 ;
  assign n57 = n56 ^ n46 ;
  assign n58 = n57 ^ n48 ;
  assign n59 = ~n48 & n58 ;
  assign n60 = n59 ^ n48 ;
  assign n61 = n50 & ~n60 ;
  assign n62 = n61 ^ n59 ;
  assign n63 = n62 ^ n46 ;
  assign n64 = n63 ^ n48 ;
  assign n65 = x0 & n64 ;
  assign n66 = n65 ^ n45 ;
  assign n67 = n37 & n66 ;
  assign n68 = x1 & n17 ;
  assign n69 = x0 & x13 ;
  assign n70 = n52 & n69 ;
  assign n71 = n68 & n70 ;
  assign n72 = ~n67 & ~n71 ;
  assign n73 = n72 ^ x5 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = ~x0 & ~x1 ;
  assign n76 = x2 & x13 ;
  assign n77 = ~x8 & n76 ;
  assign n78 = n75 & n77 ;
  assign n79 = x10 & x14 ;
  assign n80 = ~x3 & x4 ;
  assign n81 = x9 & n80 ;
  assign n82 = n79 & n81 ;
  assign n83 = n82 ^ x6 ;
  assign n84 = n83 ^ n82 ;
  assign n85 = x7 & ~x9 ;
  assign n86 = x3 & ~x14 ;
  assign n87 = n85 & n86 ;
  assign n88 = ~x4 & n87 ;
  assign n89 = n88 ^ n82 ;
  assign n90 = n84 & n89 ;
  assign n91 = n90 ^ n82 ;
  assign n92 = n78 & n91 ;
  assign n93 = n92 ^ n72 ;
  assign n94 = n74 & ~n93 ;
  assign n95 = n94 ^ n72 ;
  assign n96 = n16 & ~n95 ;
  assign y0 = n96 ;
endmodule
