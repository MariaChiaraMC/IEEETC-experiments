module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 ;
  assign n9 = ~x0 & x3 ;
  assign n10 = x4 & ~n9 ;
  assign n11 = x0 & ~x5 ;
  assign n12 = ~x2 & ~n11 ;
  assign n13 = n10 & ~n12 ;
  assign n14 = x2 & ~x4 ;
  assign n15 = x6 & x7 ;
  assign n16 = ~x3 & n15 ;
  assign n17 = n16 ^ x1 ;
  assign n18 = n14 & ~n17 ;
  assign n19 = n18 ^ x1 ;
  assign n20 = ~n13 & ~n19 ;
  assign n21 = x6 ^ x3 ;
  assign n22 = x0 & n21 ;
  assign n23 = n22 ^ x3 ;
  assign n24 = ~x2 & n23 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = n24 ^ n9 ;
  assign n27 = n26 ^ n9 ;
  assign n28 = ~x5 & x6 ;
  assign n29 = ~x7 & n28 ;
  assign n30 = ~n11 & ~n29 ;
  assign n31 = n30 ^ n9 ;
  assign n32 = ~n27 & ~n31 ;
  assign n33 = n32 ^ n9 ;
  assign n34 = ~n25 & n33 ;
  assign n35 = n34 ^ x4 ;
  assign n36 = n20 & n35 ;
  assign y0 = ~n36 ;
endmodule
