module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n12 = ~x2 & ~x3 ;
  assign n13 = x6 & x7 ;
  assign n14 = x5 & x8 ;
  assign n15 = n13 & n14 ;
  assign n16 = x4 & n15 ;
  assign n17 = ~n12 & n16 ;
  assign n18 = ~x9 & ~n17 ;
  assign n19 = ~x10 & n18 ;
  assign n20 = ~x7 & ~x8 ;
  assign n21 = x6 ^ x5 ;
  assign n22 = n20 & ~n21 ;
  assign n23 = x2 & x4 ;
  assign n24 = x3 & n23 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = x0 & x1 ;
  assign n28 = ~x5 & ~n27 ;
  assign n29 = n28 ^ n22 ;
  assign n30 = ~n26 & n29 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n22 & n31 ;
  assign n33 = n32 ^ n20 ;
  assign n34 = n19 & ~n33 ;
  assign y0 = ~n34 ;
endmodule
