module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 ;
  assign n12 = x6 ^ x5 ;
  assign n13 = n12 ^ x5 ;
  assign n16 = ~x0 & ~x10 ;
  assign n14 = ~x7 & ~x9 ;
  assign n15 = n14 ^ n12 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = ~n13 & n17 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = n12 ^ x8 ;
  assign n22 = n21 ^ n15 ;
  assign n23 = x3 & x4 ;
  assign n24 = x1 & ~x2 ;
  assign n25 = n23 & n24 ;
  assign n26 = n25 ^ n12 ;
  assign n27 = ~n22 & n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n28 ^ n12 ;
  assign n30 = n29 ^ n15 ;
  assign n31 = n30 ^ n21 ;
  assign n32 = n31 ^ n16 ;
  assign n33 = n15 ^ n12 ;
  assign n34 = n16 & ~n33 ;
  assign n35 = n34 ^ n15 ;
  assign n36 = n35 ^ n21 ;
  assign n37 = n36 ^ n16 ;
  assign n38 = ~n32 & ~n37 ;
  assign n39 = n38 ^ n21 ;
  assign n40 = ~n20 & ~n39 ;
  assign n41 = n40 ^ n34 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = n42 ^ n15 ;
  assign n44 = n43 ^ n21 ;
  assign n45 = n44 ^ n16 ;
  assign y0 = ~n45 ;
endmodule
