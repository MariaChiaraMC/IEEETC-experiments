module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ;
  assign n21 = x0 & ~x2 ;
  assign n22 = ~x1 & x3 ;
  assign n23 = x4 & n22 ;
  assign n24 = ~n21 & n23 ;
  assign n9 = x3 ^ x0 ;
  assign n10 = n9 ^ x2 ;
  assign n11 = n10 ^ x4 ;
  assign n12 = x1 ^ x0 ;
  assign n13 = ~x1 & ~n12 ;
  assign n14 = n13 ^ x2 ;
  assign n15 = n14 ^ x1 ;
  assign n16 = n11 & n15 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n17 ^ x1 ;
  assign n19 = ~x4 & ~n18 ;
  assign n20 = n19 ^ x3 ;
  assign n25 = n24 ^ n20 ;
  assign n26 = ~x6 & ~x7 ;
  assign n27 = n26 ^ x5 ;
  assign n28 = n27 ^ x5 ;
  assign n29 = n28 ^ n25 ;
  assign n30 = x5 ^ x2 ;
  assign n31 = n30 ^ n24 ;
  assign n32 = n24 & ~n31 ;
  assign n33 = n32 ^ x5 ;
  assign n34 = n33 ^ n24 ;
  assign n35 = ~n29 & ~n34 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ n24 ;
  assign n38 = ~n25 & n37 ;
  assign n39 = n38 ^ n20 ;
  assign y0 = ~n39 ;
endmodule
