module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n9 = x2 & ~x3 ;
  assign n10 = x4 & x5 ;
  assign n11 = n9 & ~n10 ;
  assign n12 = x0 & ~n11 ;
  assign n13 = x1 & n12 ;
  assign n14 = x3 ^ x2 ;
  assign n15 = x7 ^ x2 ;
  assign n16 = n14 & ~n15 ;
  assign n17 = x6 & n16 ;
  assign n18 = n13 & ~n17 ;
  assign n19 = x3 & ~x5 ;
  assign n20 = ~x4 & n19 ;
  assign n21 = ~x0 & ~n20 ;
  assign n22 = n21 ^ x2 ;
  assign n23 = ~x3 & x4 ;
  assign n24 = n23 ^ x2 ;
  assign n25 = ~n22 & ~n24 ;
  assign n26 = n25 ^ x2 ;
  assign n27 = ~x1 & ~n26 ;
  assign n28 = ~n18 & ~n27 ;
  assign y0 = ~n28 ;
endmodule
