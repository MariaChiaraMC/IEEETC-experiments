module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 ;
  output y0 ;
  wire n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 ;
  assign n26 = ~x0 & ~x4 ;
  assign n27 = ~x5 & ~x20 ;
  assign n28 = ~x23 & n27 ;
  assign n29 = ~x1 & ~x2 ;
  assign n30 = ~x3 & n29 ;
  assign n31 = n28 & n30 ;
  assign n32 = n26 & n31 ;
  assign n33 = ~x22 & ~x24 ;
  assign n34 = ~x17 & ~x18 ;
  assign n35 = ~x19 & n34 ;
  assign n36 = ~x21 & n35 ;
  assign n37 = n33 & n36 ;
  assign n38 = n32 & n37 ;
  assign n39 = x14 & n38 ;
  assign n40 = x0 & x22 ;
  assign n41 = x17 & x19 ;
  assign n42 = n40 & n41 ;
  assign n43 = x2 & x24 ;
  assign n44 = x4 & n43 ;
  assign n45 = n42 & n44 ;
  assign n46 = x3 & x21 ;
  assign n47 = x1 & n46 ;
  assign n48 = n45 & n47 ;
  assign n49 = x18 & x23 ;
  assign n50 = x20 & n49 ;
  assign n51 = x5 & n50 ;
  assign n52 = n48 & n51 ;
  assign n53 = x6 & n52 ;
  assign n54 = ~n39 & ~n53 ;
  assign n55 = x9 ^ x8 ;
  assign n56 = x9 & ~n55 ;
  assign n57 = x7 & n56 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = ~n54 & ~n58 ;
  assign n60 = x15 & n38 ;
  assign n61 = x10 & n52 ;
  assign n62 = ~n60 & ~n61 ;
  assign n63 = ~x11 & ~x12 ;
  assign n64 = ~x7 & n63 ;
  assign n65 = ~n62 & n64 ;
  assign n66 = x16 & n38 ;
  assign n67 = x13 & n52 ;
  assign n68 = ~n66 & ~n67 ;
  assign n69 = ~x8 & ~x9 ;
  assign n70 = x7 & ~n69 ;
  assign n71 = ~n68 & n70 ;
  assign n72 = ~n65 & ~n71 ;
  assign n73 = ~n59 & n72 ;
  assign y0 = ~n73 ;
endmodule
