module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n9 = x4 ^ x2 ;
  assign n10 = n9 ^ x5 ;
  assign n22 = n10 ^ x4 ;
  assign n15 = x7 ^ x4 ;
  assign n11 = n10 ^ x5 ;
  assign n12 = n11 ^ x7 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = n16 ^ x4 ;
  assign n18 = n10 ^ x6 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = ~n17 & n19 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n23 ^ x1 ;
  assign n13 = n12 ^ x4 ;
  assign n14 = ~x4 & n13 ;
  assign n25 = n22 ^ n14 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = n24 & ~n26 ;
  assign n21 = n20 ^ n14 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = n28 ^ n22 ;
  assign n30 = n29 ^ x1 ;
  assign n31 = x1 & n30 ;
  assign n32 = n31 ^ n20 ;
  assign n33 = n32 ^ n14 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = n34 ^ n22 ;
  assign n36 = n35 ^ x1 ;
  assign n37 = n36 ^ x2 ;
  assign y0 = n37 ;
endmodule
