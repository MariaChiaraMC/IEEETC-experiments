module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 ;
  assign n11 = ~x6 & ~x7 ;
  assign n12 = ~x4 & ~x5 ;
  assign n13 = n11 & n12 ;
  assign n14 = x2 & ~n13 ;
  assign n15 = x4 & x5 ;
  assign n16 = ~x0 & ~x1 ;
  assign n17 = ~n15 & n16 ;
  assign n18 = ~n14 & n17 ;
  assign n19 = n12 ^ x7 ;
  assign n20 = n12 ^ x6 ;
  assign n21 = n20 ^ n12 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = x8 ^ x3 ;
  assign n24 = ~n12 & ~n23 ;
  assign n25 = n24 ^ x3 ;
  assign n26 = n22 & ~n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n27 ^ x3 ;
  assign n29 = n28 ^ n12 ;
  assign n30 = ~n19 & n29 ;
  assign n31 = n30 ^ x7 ;
  assign n32 = n18 & ~n31 ;
  assign n39 = x3 ^ x2 ;
  assign n36 = x9 ^ x3 ;
  assign n37 = n36 ^ x9 ;
  assign n40 = n39 ^ n37 ;
  assign n33 = ~x6 & ~x8 ;
  assign n34 = n33 ^ n13 ;
  assign n35 = n34 ^ x9 ;
  assign n38 = n37 ^ n35 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n39 ^ n33 ;
  assign n43 = n42 ^ n35 ;
  assign n44 = n43 ^ n40 ;
  assign n45 = n43 ^ n37 ;
  assign n46 = ~n44 & ~n45 ;
  assign n47 = n46 ^ n35 ;
  assign n48 = n47 ^ n40 ;
  assign n49 = n39 ^ x9 ;
  assign n50 = n49 ^ n42 ;
  assign n51 = n50 ^ n35 ;
  assign n52 = ~n37 & ~n51 ;
  assign n53 = n52 ^ n37 ;
  assign n54 = n53 ^ n40 ;
  assign n55 = n48 & n54 ;
  assign n56 = ~n41 & n55 ;
  assign n57 = n56 ^ n46 ;
  assign n58 = n57 ^ n52 ;
  assign n59 = n58 ^ n42 ;
  assign n60 = n59 ^ n35 ;
  assign n61 = n60 ^ n40 ;
  assign n62 = n32 & ~n61 ;
  assign y0 = n62 ;
endmodule
