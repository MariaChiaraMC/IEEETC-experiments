module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n8 = ~x2 & x5 ;
  assign n9 = x3 & ~x4 ;
  assign n10 = ~n8 & ~n9 ;
  assign n11 = ~x0 & ~n10 ;
  assign n12 = x5 ^ x1 ;
  assign n13 = n12 ^ x5 ;
  assign n14 = x6 ^ x5 ;
  assign n15 = n14 ^ x6 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n14 ^ x2 ;
  assign n18 = n16 & ~n17 ;
  assign n19 = n18 ^ n14 ;
  assign n20 = ~x3 & x4 ;
  assign n21 = ~n14 & n20 ;
  assign n22 = n21 ^ n13 ;
  assign n23 = ~n19 & n22 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n13 & n24 ;
  assign n26 = n25 ^ n12 ;
  assign n27 = n26 ^ n13 ;
  assign n28 = n11 & ~n27 ;
  assign y0 = n28 ;
endmodule
