module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 ;
  assign n13 = x9 ^ x5 ;
  assign n14 = n13 ^ x11 ;
  assign n15 = n14 ^ x1 ;
  assign n16 = x6 & ~x7 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = x11 & n18 ;
  assign n20 = n19 ^ x5 ;
  assign n21 = n20 ^ x11 ;
  assign n22 = n21 ^ n14 ;
  assign n23 = n22 ^ x1 ;
  assign n24 = n15 & ~n23 ;
  assign n25 = n24 ^ n19 ;
  assign n26 = n25 ^ x5 ;
  assign n27 = n26 ^ n14 ;
  assign n28 = ~x1 & n27 ;
  assign n29 = n28 ^ x1 ;
  assign n30 = n29 ^ x1 ;
  assign n31 = ~x3 & n30 ;
  assign n32 = ~x0 & ~n31 ;
  assign n33 = x8 ^ x0 ;
  assign n34 = x8 ^ x6 ;
  assign n35 = n34 ^ x6 ;
  assign n36 = x7 ^ x6 ;
  assign n37 = ~n35 & n36 ;
  assign n38 = n37 ^ x6 ;
  assign n39 = n33 & n38 ;
  assign n40 = n39 ^ x0 ;
  assign n41 = ~n32 & ~n40 ;
  assign y0 = n41 ;
endmodule
