module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 ;
  assign n9 = x0 & ~x1 ;
  assign n10 = n9 ^ x6 ;
  assign n11 = x5 ^ x0 ;
  assign n12 = x7 ^ x2 ;
  assign n13 = x1 & ~x4 ;
  assign n14 = n13 ^ x2 ;
  assign n15 = n12 & ~n14 ;
  assign n16 = n15 ^ x2 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = ~n11 & ~n17 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n19 ^ x2 ;
  assign n21 = n20 ^ x0 ;
  assign n22 = x5 & n21 ;
  assign n23 = n22 ^ x5 ;
  assign n24 = n23 ^ n9 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ n10 ;
  assign n27 = ~x5 & ~x7 ;
  assign n28 = x4 & ~n27 ;
  assign n29 = x2 & x7 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = n28 & ~n30 ;
  assign n32 = n31 ^ n23 ;
  assign n33 = n32 ^ n28 ;
  assign n34 = ~n26 & n33 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = n35 ^ n28 ;
  assign n37 = ~n10 & n36 ;
  assign n38 = n37 ^ n9 ;
  assign n39 = x2 & x4 ;
  assign n40 = x1 & ~x6 ;
  assign n41 = ~n39 & n40 ;
  assign n42 = n41 ^ x2 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = ~x6 & ~x7 ;
  assign n45 = ~x4 & n44 ;
  assign n46 = n45 ^ n41 ;
  assign n47 = n43 & ~n46 ;
  assign n48 = n47 ^ n41 ;
  assign n49 = x7 & ~n41 ;
  assign n50 = n49 ^ x0 ;
  assign n51 = ~n48 & ~n50 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = ~x0 & n52 ;
  assign n54 = n53 ^ x0 ;
  assign n56 = ~x2 & ~x4 ;
  assign n55 = ~x1 & ~x7 ;
  assign n57 = n56 ^ n55 ;
  assign n58 = x6 & n57 ;
  assign n59 = n58 ^ n56 ;
  assign n60 = n54 & ~n59 ;
  assign n61 = ~x5 & ~n60 ;
  assign n62 = ~x6 & x7 ;
  assign n63 = x4 & ~n62 ;
  assign n64 = x1 & ~n44 ;
  assign n65 = ~n63 & ~n64 ;
  assign n66 = ~x2 & n65 ;
  assign n67 = ~x4 & x6 ;
  assign n68 = ~x0 & x1 ;
  assign n69 = x5 & n68 ;
  assign n70 = n69 ^ x0 ;
  assign n71 = n70 ^ n69 ;
  assign n72 = x5 & x7 ;
  assign n73 = n72 ^ n69 ;
  assign n74 = n73 ^ n69 ;
  assign n75 = n71 & n74 ;
  assign n76 = n75 ^ n69 ;
  assign n77 = ~x2 & n76 ;
  assign n78 = n77 ^ n69 ;
  assign n79 = n67 & n78 ;
  assign n80 = x4 & x5 ;
  assign n81 = ~x1 & n80 ;
  assign n82 = x7 & n81 ;
  assign n83 = ~x1 & n39 ;
  assign n84 = ~n9 & ~n83 ;
  assign n85 = ~n82 & n84 ;
  assign n86 = ~n79 & n85 ;
  assign n87 = ~n66 & n86 ;
  assign n88 = ~n61 & n87 ;
  assign n89 = n88 ^ x3 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = x5 ^ x4 ;
  assign n92 = ~x6 & n91 ;
  assign n93 = n92 ^ x4 ;
  assign n94 = n93 ^ x0 ;
  assign n95 = n94 ^ x1 ;
  assign n102 = n95 ^ n94 ;
  assign n96 = n95 ^ n45 ;
  assign n97 = n96 ^ n94 ;
  assign n98 = n95 ^ n93 ;
  assign n99 = n98 ^ n45 ;
  assign n100 = n99 ^ n97 ;
  assign n101 = n97 & n100 ;
  assign n103 = n102 ^ n101 ;
  assign n104 = n103 ^ n97 ;
  assign n105 = ~n62 & ~n80 ;
  assign n106 = n105 ^ n94 ;
  assign n107 = n101 ^ n97 ;
  assign n108 = n106 & n107 ;
  assign n109 = n108 ^ n94 ;
  assign n110 = ~n104 & n109 ;
  assign n111 = n110 ^ n94 ;
  assign n112 = n111 ^ x0 ;
  assign n113 = n112 ^ n94 ;
  assign n114 = x2 & ~n113 ;
  assign n115 = ~x2 & ~x7 ;
  assign n116 = x4 & ~x5 ;
  assign n117 = ~n115 & ~n116 ;
  assign n118 = n68 & ~n117 ;
  assign n119 = ~x2 & n81 ;
  assign n120 = ~n118 & ~n119 ;
  assign n121 = n120 ^ x1 ;
  assign n122 = n121 ^ x6 ;
  assign n129 = n122 ^ n121 ;
  assign n124 = ~x4 & ~n72 ;
  assign n123 = n122 ^ n120 ;
  assign n125 = n124 ^ n123 ;
  assign n126 = n124 ^ n122 ;
  assign n127 = n126 ^ n121 ;
  assign n128 = ~n125 & ~n127 ;
  assign n130 = n129 ^ n128 ;
  assign n131 = n122 ^ n27 ;
  assign n132 = n129 & n131 ;
  assign n133 = n132 ^ n27 ;
  assign n134 = n130 & n133 ;
  assign n135 = n134 ^ n128 ;
  assign n136 = n135 ^ n122 ;
  assign n137 = n136 ^ x1 ;
  assign n138 = n137 ^ n121 ;
  assign n139 = ~n114 & n138 ;
  assign n140 = n139 ^ n88 ;
  assign n141 = n90 & n140 ;
  assign n142 = n141 ^ n88 ;
  assign n143 = ~n38 & n142 ;
  assign y0 = ~n143 ;
endmodule
