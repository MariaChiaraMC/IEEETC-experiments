module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;
  assign n9 = ~x4 & x5 ;
  assign n10 = n9 ^ x2 ;
  assign n11 = n9 ^ x0 ;
  assign n12 = x3 & ~n11 ;
  assign n13 = n12 ^ x6 ;
  assign n14 = x2 & ~n13 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n10 & n15 ;
  assign n17 = n16 ^ n9 ;
  assign n18 = n17 ^ n12 ;
  assign n19 = n18 ^ n14 ;
  assign n20 = n19 ^ x2 ;
  assign n21 = x3 ^ x0 ;
  assign n23 = ~x4 & x6 ;
  assign n24 = ~x7 & n23 ;
  assign n22 = n21 ^ x3 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = ~n21 & ~n25 ;
  assign n27 = n26 ^ x3 ;
  assign n28 = ~x1 & ~x2 ;
  assign n29 = n28 ^ n21 ;
  assign n30 = n9 ^ x1 ;
  assign n31 = n30 ^ x3 ;
  assign n32 = n30 ^ n21 ;
  assign n33 = n31 & ~n32 ;
  assign n34 = n33 ^ x1 ;
  assign n35 = n34 ^ n21 ;
  assign n36 = n35 ^ n24 ;
  assign n37 = ~n29 & n36 ;
  assign n38 = n37 ^ n21 ;
  assign n39 = n38 ^ n24 ;
  assign n40 = n27 & ~n39 ;
  assign n41 = n40 ^ n26 ;
  assign n42 = n41 ^ x3 ;
  assign n43 = ~n20 & n42 ;
  assign y0 = ~n43 ;
endmodule
