// Benchmark "./newapla1.pla" written by ABC on Thu Apr 23 10:59:57 2020

module \./newapla1.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11,
    z0  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11;
  output z0;
  assign z0 = 1'b1;
endmodule


