module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n8 = x4 ^ x3 ;
  assign n9 = ~x5 & ~x6 ;
  assign n10 = n9 ^ x1 ;
  assign n11 = x1 ^ x0 ;
  assign n12 = n11 ^ n9 ;
  assign n13 = ~n9 & ~n12 ;
  assign n14 = n13 ^ n9 ;
  assign n15 = n10 & ~n14 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = n16 ^ n9 ;
  assign n18 = n17 ^ n11 ;
  assign n19 = n8 & ~n18 ;
  assign n20 = n19 ^ x0 ;
  assign n21 = n20 ^ x0 ;
  assign n22 = x0 & ~x1 ;
  assign n23 = ~x3 & ~x4 ;
  assign n24 = n22 & n23 ;
  assign n25 = x6 ^ x5 ;
  assign n26 = n24 & n25 ;
  assign n27 = n26 ^ x0 ;
  assign n28 = n27 ^ x0 ;
  assign n29 = ~n21 & ~n28 ;
  assign n30 = n29 ^ x0 ;
  assign n31 = x2 & ~n30 ;
  assign n32 = n31 ^ x0 ;
  assign y0 = n32 ;
endmodule
