module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 ;
  assign n11 = ~x2 & x6 ;
  assign n32 = x5 & ~x9 ;
  assign n33 = ~x3 & x7 ;
  assign n34 = n32 & ~n33 ;
  assign n35 = ~n11 & n34 ;
  assign n12 = x0 & x2 ;
  assign n13 = ~x6 & ~n12 ;
  assign n14 = ~x7 & n13 ;
  assign n15 = x3 & ~n14 ;
  assign n16 = n15 ^ x8 ;
  assign n17 = n15 ^ x2 ;
  assign n18 = n15 ^ x7 ;
  assign n19 = n15 & ~n18 ;
  assign n20 = n19 ^ n15 ;
  assign n21 = n17 & n20 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ n15 ;
  assign n24 = n23 ^ x7 ;
  assign n25 = n16 & ~n24 ;
  assign n26 = n25 ^ n15 ;
  assign n27 = x9 ^ x5 ;
  assign n28 = n26 & ~n27 ;
  assign n29 = ~n11 & n28 ;
  assign n30 = ~x1 & ~n29 ;
  assign n31 = x4 & ~n30 ;
  assign n36 = n35 ^ n31 ;
  assign n37 = n31 ^ x1 ;
  assign n38 = n37 ^ x1 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = ~x3 & ~x7 ;
  assign n41 = x4 & ~n40 ;
  assign n42 = ~n14 & n41 ;
  assign n43 = n42 ^ x8 ;
  assign n44 = ~x8 & n43 ;
  assign n45 = n44 ^ x1 ;
  assign n46 = n45 ^ x8 ;
  assign n47 = ~n39 & ~n46 ;
  assign n48 = n47 ^ n44 ;
  assign n49 = n48 ^ x8 ;
  assign n50 = n36 & ~n49 ;
  assign n51 = n50 ^ n31 ;
  assign y0 = n51 ;
endmodule
