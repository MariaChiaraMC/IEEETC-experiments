module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 ;
  output y0 ;
  wire n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 ;
  assign n16 = x2 & x5 ;
  assign n17 = n16 ^ x2 ;
  assign n18 = n17 ^ x2 ;
  assign n14 = x8 ^ x2 ;
  assign n15 = n14 ^ x2 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = ~x6 & x7 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = n21 ^ x2 ;
  assign n23 = n22 ^ n18 ;
  assign n24 = n18 & n23 ;
  assign n25 = n24 ^ n18 ;
  assign n26 = n19 & n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n27 ^ x2 ;
  assign n29 = n28 ^ n18 ;
  assign n30 = x0 & ~n29 ;
  assign n31 = n30 ^ x2 ;
  assign n32 = x4 & ~n31 ;
  assign n33 = ~x4 & ~x5 ;
  assign n34 = n33 ^ n16 ;
  assign n35 = n34 ^ n16 ;
  assign n36 = n17 ^ n16 ;
  assign n37 = n35 & ~n36 ;
  assign n38 = n37 ^ n16 ;
  assign n39 = x0 & n38 ;
  assign n40 = n39 ^ n16 ;
  assign n41 = ~n20 & n40 ;
  assign n42 = ~n32 & ~n41 ;
  assign n43 = ~x1 & x9 ;
  assign n44 = x3 & x12 ;
  assign n45 = n43 & n44 ;
  assign n46 = x11 & n45 ;
  assign n47 = x10 & n46 ;
  assign n48 = ~n42 & n47 ;
  assign y0 = n48 ;
endmodule
