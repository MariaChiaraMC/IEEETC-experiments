module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n10 = ~x7 & ~x8 ;
  assign n11 = ~x1 & x2 ;
  assign n12 = n11 ^ x6 ;
  assign n13 = n12 ^ x4 ;
  assign n14 = n13 ^ n11 ;
  assign n15 = n14 ^ n12 ;
  assign n24 = n11 ^ x5 ;
  assign n25 = n24 ^ x5 ;
  assign n21 = n14 ^ x5 ;
  assign n22 = n21 ^ n12 ;
  assign n16 = n12 ^ x3 ;
  assign n17 = n16 ^ n12 ;
  assign n18 = n12 ^ x0 ;
  assign n19 = n18 ^ n12 ;
  assign n20 = n17 & ~n19 ;
  assign n23 = n22 ^ n20 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n15 & n26 ;
  assign n28 = n27 ^ n12 ;
  assign n29 = n28 ^ n22 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = ~n22 & ~n30 ;
  assign n32 = n31 ^ n15 ;
  assign n33 = ~n28 & n32 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = n34 ^ x6 ;
  assign n36 = n35 ^ n12 ;
  assign n37 = ~n10 & n36 ;
  assign y0 = n37 ;
endmodule
