module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 ;
  assign n73 = x11 & x13 ;
  assign n74 = x12 & n73 ;
  assign n21 = ~x17 & ~x18 ;
  assign n75 = ~x16 & n21 ;
  assign n76 = x3 & ~x5 ;
  assign n77 = ~x10 & n76 ;
  assign n78 = x1 & ~n77 ;
  assign n79 = n75 & n78 ;
  assign n80 = ~n74 & n79 ;
  assign n81 = x7 & ~x17 ;
  assign n57 = x8 & ~x18 ;
  assign n82 = ~x6 & x16 ;
  assign n83 = n57 & n82 ;
  assign n84 = n81 & n83 ;
  assign n58 = x17 & ~n57 ;
  assign n85 = ~x7 & n58 ;
  assign n25 = x16 ^ x6 ;
  assign n86 = ~x7 & x17 ;
  assign n87 = ~x8 & x18 ;
  assign n88 = ~n81 & n87 ;
  assign n89 = ~n86 & ~n88 ;
  assign n90 = ~n25 & ~n89 ;
  assign n91 = ~n85 & n90 ;
  assign n92 = ~n84 & ~n91 ;
  assign n93 = x4 & ~x9 ;
  assign n94 = ~n92 & n93 ;
  assign n95 = ~n80 & ~n94 ;
  assign n20 = ~x2 & ~x10 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n20 ^ x16 ;
  assign n24 = n23 ^ x16 ;
  assign n26 = n25 ^ x16 ;
  assign n27 = n24 & ~n26 ;
  assign n28 = n27 ^ x16 ;
  assign n29 = n22 & n28 ;
  assign n30 = n29 ^ n21 ;
  assign n31 = x9 & ~x18 ;
  assign n32 = x6 & ~n31 ;
  assign n33 = x16 & ~n32 ;
  assign n34 = ~x8 & n33 ;
  assign n37 = x17 ^ x9 ;
  assign n38 = n37 ^ x9 ;
  assign n35 = x16 ^ x9 ;
  assign n36 = n35 ^ x9 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = x9 ^ x7 ;
  assign n41 = n40 ^ x9 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = ~n38 & n42 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = ~n39 & ~n44 ;
  assign n46 = n45 ^ n43 ;
  assign n47 = n46 ^ x9 ;
  assign n48 = n47 ^ n38 ;
  assign n49 = ~x18 & ~n48 ;
  assign n50 = n49 ^ x9 ;
  assign n51 = x8 & n50 ;
  assign n52 = n51 ^ n34 ;
  assign n53 = x16 & n21 ;
  assign n54 = x6 & n53 ;
  assign n55 = n54 ^ n21 ;
  assign n56 = x7 & ~n55 ;
  assign n59 = n58 ^ n56 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = x7 & ~n31 ;
  assign n62 = n61 ^ n56 ;
  assign n63 = n60 & ~n62 ;
  assign n64 = n63 ^ n56 ;
  assign n65 = n64 ^ n34 ;
  assign n66 = n52 & n65 ;
  assign n67 = n66 ^ n63 ;
  assign n68 = n67 ^ n56 ;
  assign n69 = n68 ^ n51 ;
  assign n70 = ~n34 & n69 ;
  assign n71 = n70 ^ n34 ;
  assign n72 = n30 & ~n71 ;
  assign n96 = n95 ^ n72 ;
  assign n97 = n96 ^ n72 ;
  assign n98 = x3 & ~n75 ;
  assign n99 = n98 ^ n72 ;
  assign n100 = n99 ^ n72 ;
  assign n101 = n97 & ~n100 ;
  assign n102 = n101 ^ n72 ;
  assign n103 = ~x15 & n102 ;
  assign n104 = n103 ^ n72 ;
  assign y0 = ~n104 ;
endmodule
