module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n10 = ~x0 & ~x2 ;
  assign n11 = x5 & ~n10 ;
  assign n12 = ~x1 & ~n11 ;
  assign n13 = x4 & ~x8 ;
  assign n14 = x6 & n13 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = x2 & x3 ;
  assign n17 = ~x0 & n16 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = n17 ^ x3 ;
  assign n21 = n19 & ~n20 ;
  assign n22 = n21 ^ n17 ;
  assign n23 = n22 ^ n12 ;
  assign n24 = ~n15 & ~n23 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ n17 ;
  assign n27 = n26 ^ n14 ;
  assign n28 = ~n12 & n27 ;
  assign n29 = n28 ^ n12 ;
  assign y0 = ~n29 ;
endmodule
