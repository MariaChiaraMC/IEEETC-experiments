module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 ;
  assign n13 = ~x10 & ~x11 ;
  assign n14 = ~x9 & n13 ;
  assign n15 = ~x9 & ~n13 ;
  assign n16 = ~x4 & ~x5 ;
  assign n17 = ~x11 & ~n16 ;
  assign n18 = n17 ^ x10 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = x4 ^ x3 ;
  assign n21 = x10 & n20 ;
  assign n22 = n21 ^ x3 ;
  assign n23 = n19 & ~n22 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n24 ^ x3 ;
  assign n26 = n25 ^ x10 ;
  assign n27 = ~n15 & ~n26 ;
  assign n28 = x2 & ~n27 ;
  assign n29 = ~x2 & x9 ;
  assign n30 = ~x3 & x10 ;
  assign n31 = ~n29 & ~n30 ;
  assign n32 = n31 ^ x11 ;
  assign n33 = n31 ^ x4 ;
  assign n34 = n33 ^ x4 ;
  assign n35 = x3 & ~x10 ;
  assign n36 = x4 & x5 ;
  assign n37 = ~n35 & ~n36 ;
  assign n38 = n37 ^ x4 ;
  assign n39 = n34 & ~n38 ;
  assign n40 = n39 ^ x4 ;
  assign n41 = ~n32 & ~n40 ;
  assign n42 = n41 ^ x11 ;
  assign n43 = ~x1 & ~x6 ;
  assign n44 = x4 & ~x10 ;
  assign n45 = n17 & ~n44 ;
  assign n46 = n45 ^ n29 ;
  assign n47 = n29 ^ x3 ;
  assign n48 = n47 ^ n29 ;
  assign n49 = n48 ^ n43 ;
  assign n50 = n49 ^ x6 ;
  assign n51 = n46 & ~n50 ;
  assign n52 = n51 ^ n29 ;
  assign n53 = n43 & n52 ;
  assign n54 = n53 ^ n43 ;
  assign n55 = ~n42 & n54 ;
  assign n56 = ~n28 & n55 ;
  assign n57 = ~n14 & ~n56 ;
  assign n58 = ~x7 & x8 ;
  assign n59 = ~n57 & n58 ;
  assign n60 = ~x0 & ~n59 ;
  assign y0 = ~n60 ;
endmodule
