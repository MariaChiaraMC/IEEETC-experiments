module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n9 = x2 ^ x1 ;
  assign n10 = x5 ^ x4 ;
  assign n11 = x6 ^ x5 ;
  assign n12 = x6 ^ x3 ;
  assign n13 = x6 & ~n12 ;
  assign n14 = n13 ^ x6 ;
  assign n15 = ~n11 & n14 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = n16 ^ x6 ;
  assign n18 = n17 ^ x3 ;
  assign n19 = n10 & ~n18 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = x1 ^ x0 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = ~n20 & ~n23 ;
  assign n25 = n24 ^ n20 ;
  assign n26 = ~n21 & ~n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n27 ^ n20 ;
  assign n29 = n28 ^ n22 ;
  assign n30 = ~n9 & ~n29 ;
  assign y0 = n30 ;
endmodule
