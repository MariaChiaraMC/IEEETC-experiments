module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 ;
  assign n11 = ~x0 & x5 ;
  assign n12 = ~x4 & ~x6 ;
  assign n13 = ~x2 & n12 ;
  assign n14 = ~x1 & x9 ;
  assign n15 = ~x8 & n14 ;
  assign n16 = n13 & n15 ;
  assign n17 = n11 & n16 ;
  assign n18 = x1 & x4 ;
  assign n19 = x2 & n18 ;
  assign n20 = ~x5 & x6 ;
  assign n21 = x0 & n20 ;
  assign n22 = x8 & ~x9 ;
  assign n23 = n21 & n22 ;
  assign n24 = n19 & n23 ;
  assign n25 = ~n17 & ~n24 ;
  assign n26 = ~x7 & ~n25 ;
  assign n106 = ~x7 & ~x8 ;
  assign n169 = x0 & x5 ;
  assign n170 = n106 & n169 ;
  assign n171 = n12 & n170 ;
  assign n172 = ~x9 & n171 ;
  assign n69 = ~x6 & ~x7 ;
  assign n86 = ~x5 & n18 ;
  assign n173 = ~n69 & n86 ;
  assign n31 = x6 & x7 ;
  assign n59 = ~x8 & ~x9 ;
  assign n27 = x8 & x9 ;
  assign n174 = n59 ^ n27 ;
  assign n175 = n174 ^ n27 ;
  assign n176 = n27 ^ x0 ;
  assign n177 = n176 ^ n27 ;
  assign n178 = n175 & n177 ;
  assign n179 = n178 ^ n27 ;
  assign n180 = ~n31 & n179 ;
  assign n181 = n180 ^ n27 ;
  assign n182 = n173 & n181 ;
  assign n183 = ~n172 & ~n182 ;
  assign n184 = ~x0 & x4 ;
  assign n87 = ~x6 & x7 ;
  assign n135 = x5 & x8 ;
  assign n185 = n87 & n135 ;
  assign n186 = n185 ^ x5 ;
  assign n187 = n186 ^ n185 ;
  assign n188 = n185 ^ n106 ;
  assign n189 = n188 ^ n185 ;
  assign n190 = ~n187 & n189 ;
  assign n191 = n190 ^ n185 ;
  assign n192 = ~x9 & n191 ;
  assign n193 = n192 ^ n185 ;
  assign n194 = n184 & n193 ;
  assign n195 = n27 & n31 ;
  assign n196 = n195 ^ n169 ;
  assign n197 = n196 ^ n194 ;
  assign n199 = ~x4 & ~x5 ;
  assign n198 = n59 & n69 ;
  assign n200 = n199 ^ n198 ;
  assign n201 = ~n195 & ~n200 ;
  assign n202 = n201 ^ n199 ;
  assign n203 = ~n197 & ~n202 ;
  assign n204 = n203 ^ n201 ;
  assign n205 = n204 ^ n199 ;
  assign n206 = n205 ^ n195 ;
  assign n207 = ~n194 & n206 ;
  assign n208 = ~x1 & ~n207 ;
  assign n118 = x7 & x8 ;
  assign n119 = x9 & n118 ;
  assign n209 = ~x0 & ~x4 ;
  assign n210 = n20 & n209 ;
  assign n211 = n119 & n210 ;
  assign n212 = ~x2 & ~n211 ;
  assign n213 = ~n208 & n212 ;
  assign n214 = n183 & n213 ;
  assign n215 = x4 ^ x0 ;
  assign n216 = n215 ^ x8 ;
  assign n217 = n87 & ~n216 ;
  assign n218 = n217 ^ n87 ;
  assign n219 = x5 ^ x0 ;
  assign n220 = n219 ^ n217 ;
  assign n221 = n215 & ~n220 ;
  assign n222 = n221 ^ n215 ;
  assign n223 = n222 ^ x8 ;
  assign n224 = n218 & ~n223 ;
  assign n225 = ~x1 & n224 ;
  assign n226 = n225 ^ x2 ;
  assign n227 = x0 & ~x5 ;
  assign n228 = ~x8 & ~n227 ;
  assign n229 = ~x6 & ~n228 ;
  assign n77 = x1 & x6 ;
  assign n78 = ~x8 & n77 ;
  assign n230 = x4 & ~n78 ;
  assign n231 = ~x5 & ~x8 ;
  assign n232 = ~x1 & ~n231 ;
  assign n102 = ~x5 & x7 ;
  assign n233 = n106 ^ n102 ;
  assign n234 = ~x0 & n233 ;
  assign n235 = n234 ^ n106 ;
  assign n236 = ~n232 & n235 ;
  assign n237 = n230 & n236 ;
  assign n238 = ~n229 & n237 ;
  assign n239 = ~x1 & ~x4 ;
  assign n37 = ~x5 & ~x6 ;
  assign n240 = ~x0 & n37 ;
  assign n241 = n240 ^ x6 ;
  assign n242 = n239 & n241 ;
  assign n243 = ~n118 & n227 ;
  assign n244 = n243 ^ n106 ;
  assign n245 = n244 ^ n243 ;
  assign n246 = x6 & ~n11 ;
  assign n247 = n246 ^ n243 ;
  assign n248 = n245 & ~n247 ;
  assign n249 = n248 ^ n243 ;
  assign n250 = n242 & n249 ;
  assign n251 = ~n238 & ~n250 ;
  assign n252 = n251 ^ x9 ;
  assign n253 = n252 ^ n251 ;
  assign n254 = x5 & ~n31 ;
  assign n255 = ~n102 & n209 ;
  assign n256 = ~x8 & n255 ;
  assign n257 = x1 & n256 ;
  assign n258 = ~n254 & n257 ;
  assign n259 = ~n69 & ~n106 ;
  assign n260 = n259 ^ n185 ;
  assign n261 = n260 ^ n185 ;
  assign n262 = ~n187 & ~n261 ;
  assign n263 = n262 ^ n185 ;
  assign n264 = x0 & n263 ;
  assign n265 = n264 ^ n185 ;
  assign n266 = n239 & n265 ;
  assign n28 = x4 & x6 ;
  assign n267 = ~x1 & ~x5 ;
  assign n268 = n118 & n267 ;
  assign n269 = ~n170 & ~n268 ;
  assign n270 = n28 & ~n269 ;
  assign n271 = ~n266 & ~n270 ;
  assign n272 = ~n258 & n271 ;
  assign n273 = n272 ^ n251 ;
  assign n274 = n253 & n273 ;
  assign n275 = n274 ^ n251 ;
  assign n276 = n275 ^ n225 ;
  assign n277 = ~n226 & ~n276 ;
  assign n278 = n277 ^ n274 ;
  assign n279 = n278 ^ n251 ;
  assign n280 = n279 ^ x2 ;
  assign n281 = ~n225 & n280 ;
  assign n282 = n281 ^ n225 ;
  assign n283 = ~n214 & n282 ;
  assign n44 = ~x4 & ~x9 ;
  assign n103 = ~x2 & x8 ;
  assign n104 = n102 & n103 ;
  assign n105 = n44 & n104 ;
  assign n107 = ~x9 & n106 ;
  assign n49 = x4 & x5 ;
  assign n108 = ~x8 & ~n49 ;
  assign n109 = ~n107 & ~n108 ;
  assign n110 = x5 ^ x4 ;
  assign n36 = x7 & x9 ;
  assign n111 = n36 ^ x5 ;
  assign n112 = n110 & ~n111 ;
  assign n113 = n112 ^ x4 ;
  assign n114 = x2 & n113 ;
  assign n115 = ~n109 & n114 ;
  assign n116 = ~n105 & ~n115 ;
  assign n117 = x6 & ~n116 ;
  assign n38 = x4 & n37 ;
  assign n120 = ~n107 & ~n119 ;
  assign n121 = n38 & ~n120 ;
  assign n122 = ~x2 & n121 ;
  assign n123 = ~n117 & ~n122 ;
  assign n124 = ~x1 & ~n123 ;
  assign n32 = ~x4 & x5 ;
  assign n125 = n32 & n59 ;
  assign n126 = n87 & n125 ;
  assign n131 = n126 ^ x2 ;
  assign n152 = n131 ^ n126 ;
  assign n62 = ~x7 & ~x9 ;
  assign n127 = x2 & ~n12 ;
  assign n128 = ~n62 & ~n127 ;
  assign n129 = x1 & ~n128 ;
  assign n130 = n129 ^ n126 ;
  assign n132 = n131 ^ n130 ;
  assign n133 = n132 ^ n131 ;
  assign n134 = n133 ^ n126 ;
  assign n136 = x9 & ~n135 ;
  assign n137 = x7 ^ x5 ;
  assign n138 = n136 & n137 ;
  assign n139 = x6 & ~n138 ;
  assign n140 = x5 ^ x2 ;
  assign n141 = n140 ^ x8 ;
  assign n142 = x8 ^ x4 ;
  assign n143 = ~n110 & ~n142 ;
  assign n144 = n143 ^ x4 ;
  assign n145 = n141 & n144 ;
  assign n146 = n145 ^ x2 ;
  assign n147 = ~n139 & n146 ;
  assign n148 = n147 ^ n132 ;
  assign n149 = n148 ^ n132 ;
  assign n150 = n149 ^ n134 ;
  assign n151 = n134 & n150 ;
  assign n153 = n152 ^ n151 ;
  assign n154 = n153 ^ n134 ;
  assign n43 = x7 & ~x8 ;
  assign n155 = x4 & ~n43 ;
  assign n156 = ~n37 & ~n155 ;
  assign n157 = n156 ^ n126 ;
  assign n158 = n151 ^ n134 ;
  assign n159 = ~n157 & n158 ;
  assign n160 = n159 ^ n126 ;
  assign n161 = ~n154 & ~n160 ;
  assign n162 = n161 ^ n126 ;
  assign n163 = n162 ^ x2 ;
  assign n164 = n163 ^ n126 ;
  assign n165 = ~n124 & n164 ;
  assign n70 = n69 ^ n31 ;
  assign n71 = n31 ^ x5 ;
  assign n72 = n71 ^ n31 ;
  assign n73 = n70 & ~n72 ;
  assign n74 = n73 ^ n31 ;
  assign n75 = n14 & n74 ;
  assign n76 = ~x8 & n75 ;
  assign n79 = ~x5 & n62 ;
  assign n80 = n78 & n79 ;
  assign n81 = ~n76 & ~n80 ;
  assign n82 = x4 & ~n81 ;
  assign n45 = n43 & n44 ;
  assign n46 = n20 & n45 ;
  assign n29 = x5 & ~x7 ;
  assign n30 = n28 & n29 ;
  assign n33 = n31 & n32 ;
  assign n34 = ~n30 & ~n33 ;
  assign n35 = n27 & ~n34 ;
  assign n39 = x8 ^ x7 ;
  assign n40 = n38 & n39 ;
  assign n41 = ~n36 & n40 ;
  assign n42 = ~n35 & ~n41 ;
  assign n47 = n46 ^ n42 ;
  assign n48 = n47 ^ n42 ;
  assign n50 = n27 & n49 ;
  assign n51 = ~x6 & n50 ;
  assign n52 = n51 ^ n42 ;
  assign n53 = n52 ^ n42 ;
  assign n54 = ~n48 & ~n53 ;
  assign n55 = n54 ^ n42 ;
  assign n56 = x1 & n55 ;
  assign n57 = n56 ^ n42 ;
  assign n83 = n82 ^ n57 ;
  assign n84 = n83 ^ n57 ;
  assign n58 = x1 & n12 ;
  assign n60 = ~x7 & n27 ;
  assign n61 = ~n59 & ~n60 ;
  assign n63 = n62 ^ n61 ;
  assign n64 = x5 & ~n63 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = n58 & n65 ;
  assign n67 = n66 ^ n57 ;
  assign n68 = n67 ^ n57 ;
  assign n85 = n84 ^ n68 ;
  assign n88 = n22 & n87 ;
  assign n89 = ~n60 & ~n88 ;
  assign n90 = n86 & ~n89 ;
  assign n91 = n90 ^ n57 ;
  assign n92 = n91 ^ n57 ;
  assign n93 = n92 ^ n84 ;
  assign n94 = ~n84 & n93 ;
  assign n95 = n94 ^ n84 ;
  assign n96 = n85 & ~n95 ;
  assign n97 = n96 ^ n94 ;
  assign n98 = n97 ^ n57 ;
  assign n99 = n98 ^ n84 ;
  assign n100 = x2 & ~n99 ;
  assign n101 = n100 ^ n57 ;
  assign n166 = n165 ^ n101 ;
  assign n167 = x0 & n166 ;
  assign n168 = n167 ^ n101 ;
  assign n284 = n283 ^ n168 ;
  assign n285 = n284 ^ n283 ;
  assign n286 = x2 & x4 ;
  assign n287 = n267 & n286 ;
  assign n288 = n22 & n69 ;
  assign n289 = n287 & n288 ;
  assign n290 = n289 ^ n283 ;
  assign n291 = n290 ^ n283 ;
  assign n292 = n285 & ~n291 ;
  assign n293 = n292 ^ n283 ;
  assign n294 = x3 & ~n293 ;
  assign n295 = n294 ^ n283 ;
  assign n296 = ~n26 & ~n295 ;
  assign y0 = ~n296 ;
endmodule
