module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 ;
  assign n11 = ~x3 & ~x9 ;
  assign n12 = ~x0 & ~x8 ;
  assign n13 = n11 & ~n12 ;
  assign n14 = x4 & n13 ;
  assign n15 = ~x8 & x9 ;
  assign n16 = ~x3 & x7 ;
  assign n17 = ~n15 & ~n16 ;
  assign n18 = ~x1 & x4 ;
  assign n19 = ~n17 & n18 ;
  assign n20 = ~n14 & ~n19 ;
  assign n28 = ~x4 & x7 ;
  assign n29 = ~n15 & ~n28 ;
  assign n30 = ~x2 & ~n29 ;
  assign n21 = x7 & x8 ;
  assign n22 = ~x4 & n21 ;
  assign n23 = ~x7 & x8 ;
  assign n24 = x7 & ~x8 ;
  assign n25 = ~n23 & ~n24 ;
  assign n26 = x9 & ~n25 ;
  assign n27 = ~n22 & ~n26 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = x8 & ~x9 ;
  assign n34 = ~x4 & n33 ;
  assign n35 = n34 ^ n27 ;
  assign n36 = n35 ^ n27 ;
  assign n37 = ~n32 & ~n36 ;
  assign n38 = n37 ^ n27 ;
  assign n39 = x1 & n38 ;
  assign n40 = n39 ^ n27 ;
  assign n41 = n20 & n40 ;
  assign n42 = x5 & ~n41 ;
  assign n43 = x1 & ~x5 ;
  assign n44 = x0 & ~x9 ;
  assign n45 = ~n43 & ~n44 ;
  assign n46 = n21 & ~n45 ;
  assign n47 = ~x0 & ~x4 ;
  assign n48 = ~x1 & n47 ;
  assign n49 = x8 & x9 ;
  assign n50 = ~x7 & n49 ;
  assign n51 = x0 & x4 ;
  assign n52 = ~n50 & ~n51 ;
  assign n53 = x1 & ~x3 ;
  assign n54 = ~n15 & ~n33 ;
  assign n55 = ~n23 & n54 ;
  assign n56 = ~n53 & n55 ;
  assign n57 = ~n52 & ~n56 ;
  assign n58 = ~n15 & ~n44 ;
  assign n59 = ~x4 & ~n15 ;
  assign n60 = x7 & ~n59 ;
  assign n61 = ~n58 & n60 ;
  assign n62 = ~n57 & ~n61 ;
  assign n63 = ~n48 & ~n62 ;
  assign n64 = ~n46 & ~n63 ;
  assign n65 = ~x2 & ~n64 ;
  assign n66 = ~n42 & ~n65 ;
  assign n68 = x4 & ~x9 ;
  assign n67 = ~x1 & x8 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = n69 ^ x7 ;
  assign n71 = ~x5 & x9 ;
  assign n72 = n71 ^ n43 ;
  assign n73 = n68 & ~n72 ;
  assign n74 = n73 ^ n71 ;
  assign n75 = n70 & n74 ;
  assign n76 = n75 ^ n73 ;
  assign n77 = n76 ^ n71 ;
  assign n78 = n77 ^ n68 ;
  assign n79 = x7 & n78 ;
  assign n80 = n66 & ~n79 ;
  assign n81 = x6 & ~n80 ;
  assign n82 = ~x1 & ~x2 ;
  assign n83 = x0 & ~x4 ;
  assign n84 = ~n22 & ~n83 ;
  assign n85 = ~n54 & ~n84 ;
  assign n86 = x6 & n15 ;
  assign n87 = ~x4 & n86 ;
  assign n88 = ~n85 & ~n87 ;
  assign n89 = x3 & ~n88 ;
  assign n90 = ~x0 & ~x6 ;
  assign n91 = x4 & ~n90 ;
  assign n92 = ~x6 & ~x7 ;
  assign n93 = ~x5 & n92 ;
  assign n94 = x0 & ~n93 ;
  assign n95 = ~n91 & ~n94 ;
  assign n96 = ~n54 & ~n95 ;
  assign n97 = ~x0 & x6 ;
  assign n98 = x5 & n97 ;
  assign n99 = x0 & ~x7 ;
  assign n100 = n49 & n99 ;
  assign n101 = ~n98 & ~n100 ;
  assign n102 = ~n47 & ~n101 ;
  assign n103 = x5 & x6 ;
  assign n104 = ~x4 & ~x6 ;
  assign n105 = x7 & ~n104 ;
  assign n106 = ~n103 & ~n105 ;
  assign n107 = n44 & ~n106 ;
  assign n108 = n107 ^ n102 ;
  assign n109 = ~x4 & ~x5 ;
  assign n110 = n21 & ~n109 ;
  assign n111 = n110 ^ x9 ;
  assign n112 = n111 ^ n110 ;
  assign n113 = x5 & ~x8 ;
  assign n114 = x4 & n113 ;
  assign n115 = n114 ^ n110 ;
  assign n116 = n112 & n115 ;
  assign n117 = n116 ^ n110 ;
  assign n118 = n117 ^ n102 ;
  assign n119 = n108 & n118 ;
  assign n120 = n119 ^ n116 ;
  assign n121 = n120 ^ n110 ;
  assign n122 = n121 ^ n107 ;
  assign n123 = ~n102 & n122 ;
  assign n124 = n123 ^ n102 ;
  assign n125 = ~n96 & ~n124 ;
  assign n126 = n125 ^ n58 ;
  assign n127 = n126 ^ x3 ;
  assign n135 = n127 ^ n126 ;
  assign n128 = x5 & n16 ;
  assign n129 = n128 ^ n127 ;
  assign n130 = n129 ^ n126 ;
  assign n131 = n127 ^ n125 ;
  assign n132 = n131 ^ n128 ;
  assign n133 = n132 ^ n130 ;
  assign n134 = n130 & n133 ;
  assign n136 = n135 ^ n134 ;
  assign n137 = n136 ^ n130 ;
  assign n138 = ~x4 & x5 ;
  assign n139 = ~n28 & ~n138 ;
  assign n140 = n139 ^ n126 ;
  assign n141 = n134 ^ n130 ;
  assign n142 = n140 & n141 ;
  assign n143 = n142 ^ n126 ;
  assign n144 = ~n137 & n143 ;
  assign n145 = n144 ^ n126 ;
  assign n146 = n145 ^ n58 ;
  assign n147 = n146 ^ n126 ;
  assign n148 = ~n89 & n147 ;
  assign n149 = ~n82 & ~n148 ;
  assign n150 = x6 ^ x5 ;
  assign n151 = x7 & ~n150 ;
  assign n152 = n151 ^ x5 ;
  assign n153 = x1 & n152 ;
  assign n154 = ~x2 & n153 ;
  assign n156 = x0 & ~x2 ;
  assign n155 = ~x1 & x5 ;
  assign n157 = n156 ^ n155 ;
  assign n158 = ~x6 & x7 ;
  assign n159 = n158 ^ n156 ;
  assign n160 = ~n156 & ~n159 ;
  assign n161 = n160 ^ n156 ;
  assign n162 = n157 & ~n161 ;
  assign n163 = n162 ^ n160 ;
  assign n164 = n163 ^ n156 ;
  assign n165 = n164 ^ n158 ;
  assign n166 = ~n154 & ~n165 ;
  assign n167 = n166 ^ n154 ;
  assign n168 = n49 & n167 ;
  assign n169 = n67 & n152 ;
  assign n170 = ~n43 & ~n156 ;
  assign n171 = ~n128 & n170 ;
  assign n172 = ~n25 & ~n171 ;
  assign n173 = ~n169 & ~n172 ;
  assign n174 = n173 ^ x9 ;
  assign n175 = n174 ^ n173 ;
  assign n176 = n21 & n155 ;
  assign n177 = n21 & n156 ;
  assign n178 = x1 & ~x6 ;
  assign n179 = ~n12 & n178 ;
  assign n180 = x5 & n179 ;
  assign n181 = ~n177 & ~n180 ;
  assign n182 = ~n176 & n181 ;
  assign n183 = n182 ^ n173 ;
  assign n184 = ~n175 & n183 ;
  assign n185 = n184 ^ n173 ;
  assign n186 = x4 & ~n185 ;
  assign n187 = ~n168 & ~n186 ;
  assign n188 = ~x3 & ~x5 ;
  assign n189 = ~n59 & ~n91 ;
  assign n190 = x1 & x2 ;
  assign n191 = n189 & n190 ;
  assign n192 = ~x7 & ~x8 ;
  assign n193 = n156 ^ x4 ;
  assign n194 = n156 ^ x6 ;
  assign n195 = n194 ^ x6 ;
  assign n196 = ~x1 & x2 ;
  assign n197 = n196 ^ x6 ;
  assign n198 = ~n195 & ~n197 ;
  assign n199 = n198 ^ x6 ;
  assign n200 = n193 & n199 ;
  assign n201 = n200 ^ x4 ;
  assign n202 = ~n192 & n201 ;
  assign n203 = ~x2 & x4 ;
  assign n204 = x7 & n203 ;
  assign n205 = x1 & n204 ;
  assign n206 = ~n177 & ~n205 ;
  assign n207 = ~n202 & n206 ;
  assign n208 = n207 ^ x9 ;
  assign n209 = n208 ^ n207 ;
  assign n210 = n209 ^ n191 ;
  assign n211 = ~x4 & ~x8 ;
  assign n212 = ~n21 & ~n211 ;
  assign n213 = ~x8 & ~n92 ;
  assign n214 = ~n212 & ~n213 ;
  assign n215 = n214 ^ n156 ;
  assign n216 = n156 & ~n215 ;
  assign n217 = n216 ^ n207 ;
  assign n218 = n217 ^ n156 ;
  assign n219 = ~n210 & ~n218 ;
  assign n220 = n219 ^ n216 ;
  assign n221 = n220 ^ n156 ;
  assign n222 = ~n191 & n221 ;
  assign n223 = n222 ^ n191 ;
  assign n224 = ~n188 & n223 ;
  assign n225 = n187 & ~n224 ;
  assign n226 = ~n149 & n225 ;
  assign n227 = ~n81 & n226 ;
  assign n228 = x5 & ~x9 ;
  assign n229 = n158 & n228 ;
  assign n230 = x9 ^ x8 ;
  assign n231 = n230 ^ x9 ;
  assign n232 = n231 ^ x5 ;
  assign n233 = n232 ^ x9 ;
  assign n234 = n233 ^ n232 ;
  assign n238 = n231 ^ x6 ;
  assign n239 = n238 ^ n232 ;
  assign n240 = n232 & ~n239 ;
  assign n235 = n230 ^ x4 ;
  assign n236 = ~n231 & n235 ;
  assign n243 = n240 ^ n236 ;
  assign n237 = n236 ^ n234 ;
  assign n241 = n240 ^ n232 ;
  assign n242 = n237 & n241 ;
  assign n244 = n243 ^ n242 ;
  assign n245 = n234 & n244 ;
  assign n246 = n245 ^ n240 ;
  assign n247 = n246 ^ n242 ;
  assign n248 = n247 ^ n230 ;
  assign n249 = ~x2 & n248 ;
  assign n250 = x6 & ~x9 ;
  assign n251 = n156 & n250 ;
  assign n252 = ~x5 & x6 ;
  assign n253 = n28 & n252 ;
  assign n254 = ~n251 & ~n253 ;
  assign n257 = ~x0 & x2 ;
  assign n255 = x6 & ~x7 ;
  assign n256 = ~n33 & ~n255 ;
  assign n258 = n257 ^ n256 ;
  assign n259 = n258 ^ n254 ;
  assign n260 = n203 ^ n24 ;
  assign n261 = ~n257 & ~n260 ;
  assign n262 = n261 ^ n24 ;
  assign n263 = ~n259 & ~n262 ;
  assign n264 = n263 ^ n261 ;
  assign n265 = n264 ^ n24 ;
  assign n266 = n265 ^ n257 ;
  assign n267 = n254 & n266 ;
  assign n268 = ~n249 & n267 ;
  assign n269 = x2 & n228 ;
  assign n270 = ~n50 & ~n269 ;
  assign n271 = n270 ^ x0 ;
  assign n272 = n271 ^ x4 ;
  assign n280 = n272 ^ n271 ;
  assign n274 = x2 & ~x5 ;
  assign n275 = ~x8 & n274 ;
  assign n273 = n272 ^ n270 ;
  assign n276 = n275 ^ n273 ;
  assign n277 = n275 ^ n272 ;
  assign n278 = n277 ^ n271 ;
  assign n279 = ~n276 & n278 ;
  assign n281 = n280 ^ n279 ;
  assign n282 = ~x5 & ~x6 ;
  assign n283 = n282 ^ n272 ;
  assign n284 = ~n280 & n283 ;
  assign n285 = n284 ^ n282 ;
  assign n286 = ~n281 & n285 ;
  assign n287 = n286 ^ n279 ;
  assign n288 = n287 ^ n272 ;
  assign n289 = n288 ^ x0 ;
  assign n290 = n289 ^ n271 ;
  assign n291 = n268 & n290 ;
  assign n292 = ~n229 & n291 ;
  assign n293 = x1 & ~n292 ;
  assign n294 = ~x9 & ~n192 ;
  assign n295 = ~n257 & ~n294 ;
  assign n296 = n155 & ~n295 ;
  assign n297 = ~x5 & ~x9 ;
  assign n298 = n21 & n297 ;
  assign n299 = ~n44 & ~n97 ;
  assign n300 = n274 & ~n299 ;
  assign n301 = ~n298 & ~n300 ;
  assign n302 = ~n296 & n301 ;
  assign n303 = x4 & ~n302 ;
  assign n304 = ~x2 & x5 ;
  assign n305 = n21 & n304 ;
  assign n306 = ~x9 & n305 ;
  assign n307 = ~n303 & ~n306 ;
  assign n308 = ~n97 & ~n294 ;
  assign n309 = x2 & n138 ;
  assign n310 = ~n308 & n309 ;
  assign n311 = x2 & n99 ;
  assign n312 = ~n22 & ~n311 ;
  assign n313 = n250 & ~n312 ;
  assign n314 = ~n310 & ~n313 ;
  assign n315 = n307 & n314 ;
  assign n316 = n212 & n274 ;
  assign n317 = ~n22 & ~n114 ;
  assign n318 = ~x6 & ~n317 ;
  assign n319 = n113 & n156 ;
  assign n320 = ~n318 & ~n319 ;
  assign n321 = ~n103 & n192 ;
  assign n322 = ~n282 & ~n321 ;
  assign n323 = ~x4 & ~n21 ;
  assign n324 = n322 & n323 ;
  assign n325 = x4 & ~x5 ;
  assign n326 = ~n23 & ~n213 ;
  assign n327 = n325 & ~n326 ;
  assign n328 = ~n324 & ~n327 ;
  assign n329 = n320 & n328 ;
  assign n330 = ~n316 & n329 ;
  assign n331 = x9 & ~n330 ;
  assign n332 = n250 ^ x0 ;
  assign n333 = n250 ^ n155 ;
  assign n334 = n333 ^ n155 ;
  assign n335 = n192 ^ n155 ;
  assign n336 = n334 & n335 ;
  assign n337 = n336 ^ n155 ;
  assign n338 = n332 & ~n337 ;
  assign n339 = n338 ^ x0 ;
  assign n340 = ~n98 & ~n339 ;
  assign n341 = n203 & ~n340 ;
  assign n342 = x5 & n251 ;
  assign n343 = n304 ^ x6 ;
  assign n344 = n343 ^ n294 ;
  assign n345 = n196 ^ x0 ;
  assign n346 = x6 & ~n345 ;
  assign n347 = n346 ^ x0 ;
  assign n348 = n344 & n347 ;
  assign n349 = n348 ^ n346 ;
  assign n350 = n349 ^ x0 ;
  assign n351 = n350 ^ x6 ;
  assign n352 = n294 & n351 ;
  assign n353 = ~n342 & ~n352 ;
  assign n354 = ~n341 & n353 ;
  assign n355 = ~n331 & n354 ;
  assign n356 = n315 & n355 ;
  assign n357 = ~n293 & n356 ;
  assign n358 = x3 & ~n357 ;
  assign n359 = ~x6 & ~x8 ;
  assign n360 = ~n49 & n99 ;
  assign n361 = ~n359 & n360 ;
  assign n362 = ~n298 & ~n361 ;
  assign n363 = ~n68 & ~n252 ;
  assign n364 = n16 & ~n363 ;
  assign n365 = ~x4 & n50 ;
  assign n366 = ~n364 & ~n365 ;
  assign n367 = ~x3 & ~n92 ;
  assign n368 = ~n83 & ~n325 ;
  assign n369 = ~n367 & n368 ;
  assign n370 = n15 & ~n369 ;
  assign n371 = ~n24 & ~n325 ;
  assign n372 = n44 & ~n371 ;
  assign n373 = ~n211 & ~n359 ;
  assign n374 = n11 & ~n104 ;
  assign n375 = n373 & n374 ;
  assign n376 = ~n372 & ~n375 ;
  assign n377 = ~n370 & n376 ;
  assign n378 = n366 & n377 ;
  assign n379 = n362 & n378 ;
  assign n380 = x1 & ~n379 ;
  assign n381 = ~x6 & n16 ;
  assign n382 = n49 & n381 ;
  assign n383 = ~n380 & ~n382 ;
  assign n384 = n18 & n44 ;
  assign n385 = ~n365 & ~n384 ;
  assign n386 = n28 & n53 ;
  assign n387 = n99 & n178 ;
  assign n388 = ~n386 & ~n387 ;
  assign n389 = x1 & ~n256 ;
  assign n390 = ~n192 & n250 ;
  assign n391 = ~n86 & ~n390 ;
  assign n392 = ~n389 & n391 ;
  assign n393 = ~x3 & ~n392 ;
  assign n394 = n388 & ~n393 ;
  assign n395 = n385 & n394 ;
  assign n396 = x5 & ~n395 ;
  assign n397 = n26 & ~n104 ;
  assign n398 = x7 & ~n211 ;
  assign n399 = ~n51 & ~n398 ;
  assign n400 = n250 & ~n399 ;
  assign n401 = ~n397 & ~n400 ;
  assign n402 = ~x3 & ~n401 ;
  assign n403 = ~n396 & ~n402 ;
  assign n404 = n383 & n403 ;
  assign n405 = x2 & ~n404 ;
  assign n406 = ~n358 & ~n405 ;
  assign n407 = n227 & n406 ;
  assign y0 = ~n407 ;
endmodule
