module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 ;
  assign n9 = ~x1 & ~x5 ;
  assign n10 = ~x4 & ~x7 ;
  assign n11 = ~x3 & ~n10 ;
  assign n12 = x6 ^ x4 ;
  assign n13 = x2 & n12 ;
  assign n14 = ~n11 & ~n13 ;
  assign n15 = n9 & ~n14 ;
  assign n16 = ~x1 & ~x4 ;
  assign n17 = ~x3 & ~n16 ;
  assign n18 = x5 & ~x7 ;
  assign n19 = x6 & n18 ;
  assign n20 = ~n17 & n19 ;
  assign n21 = x3 & x7 ;
  assign n22 = ~n18 & ~n21 ;
  assign n23 = ~x6 & ~n22 ;
  assign n24 = x6 & x7 ;
  assign n25 = ~x3 & n24 ;
  assign n26 = ~x1 & ~n25 ;
  assign n27 = ~n23 & n26 ;
  assign n28 = x4 & ~n27 ;
  assign n34 = x7 ^ x3 ;
  assign n32 = x3 ^ x1 ;
  assign n33 = n32 ^ x3 ;
  assign n35 = n34 ^ n33 ;
  assign n36 = n35 ^ x3 ;
  assign n29 = x5 ^ x3 ;
  assign n30 = n29 ^ x6 ;
  assign n31 = n30 ^ x3 ;
  assign n37 = n36 ^ n31 ;
  assign n38 = n30 ^ x6 ;
  assign n39 = n38 ^ n33 ;
  assign n40 = n39 ^ n31 ;
  assign n41 = n37 & ~n40 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = n39 ^ n30 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = n40 ^ n38 ;
  assign n46 = ~n44 & ~n45 ;
  assign n47 = n46 ^ n39 ;
  assign n48 = n47 ^ n36 ;
  assign n49 = n38 ^ n36 ;
  assign n50 = x4 ^ x3 ;
  assign n51 = n50 ^ x3 ;
  assign n52 = n51 ^ x3 ;
  assign n53 = n52 ^ n39 ;
  assign n54 = n49 & ~n53 ;
  assign n55 = n54 ^ n51 ;
  assign n56 = n55 ^ n30 ;
  assign n57 = ~n48 & n56 ;
  assign n58 = n57 ^ n30 ;
  assign n59 = ~n42 & n58 ;
  assign n60 = n59 ^ n46 ;
  assign n61 = n60 ^ n41 ;
  assign n62 = n61 ^ n57 ;
  assign n63 = n62 ^ n30 ;
  assign n64 = n63 ^ n39 ;
  assign n65 = n64 ^ n32 ;
  assign n66 = n65 ^ x3 ;
  assign n67 = ~n28 & ~n66 ;
  assign n68 = ~n20 & n67 ;
  assign n69 = n68 ^ x2 ;
  assign n70 = n69 ^ n68 ;
  assign n71 = x3 & x5 ;
  assign n72 = n16 & n71 ;
  assign n73 = n72 ^ n68 ;
  assign n74 = n70 & ~n73 ;
  assign n75 = n74 ^ n68 ;
  assign n76 = ~n15 & n75 ;
  assign y0 = ~n76 ;
endmodule
