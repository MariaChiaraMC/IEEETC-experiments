module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n10 = ~x6 & x7 ;
  assign n29 = ~x4 & n10 ;
  assign n9 = x4 & x5 ;
  assign n11 = ~x2 & n10 ;
  assign n12 = n9 & n11 ;
  assign n13 = ~x1 & ~n12 ;
  assign n14 = x6 & ~n9 ;
  assign n15 = x7 ^ x5 ;
  assign n16 = n15 ^ x2 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = x4 ^ x2 ;
  assign n20 = x4 & n19 ;
  assign n21 = n20 ^ x5 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = ~n18 & n22 ;
  assign n24 = n23 ^ n20 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = n14 & n25 ;
  assign n27 = n13 & ~n26 ;
  assign n28 = x0 & ~n27 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = n28 ^ x5 ;
  assign n32 = n31 ^ x5 ;
  assign n33 = x5 ^ x1 ;
  assign n34 = n32 & ~n33 ;
  assign n35 = n34 ^ x5 ;
  assign n36 = n30 & n35 ;
  assign n37 = n36 ^ n29 ;
  assign n38 = ~x3 & n37 ;
  assign y0 = n38 ;
endmodule
