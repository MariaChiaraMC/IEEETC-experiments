module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 ;
  assign n9 = ~x0 & x7 ;
  assign n10 = x5 & ~x6 ;
  assign n11 = x5 ^ x4 ;
  assign n12 = x4 ^ x2 ;
  assign n13 = ~n11 & n12 ;
  assign n14 = n13 ^ x4 ;
  assign n15 = ~n10 & ~n14 ;
  assign n16 = ~x1 & n15 ;
  assign n17 = ~x4 & ~x6 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = x4 & x6 ;
  assign n21 = x1 & ~n20 ;
  assign n22 = ~n17 & n21 ;
  assign n23 = n22 ^ n17 ;
  assign n24 = ~n19 & n23 ;
  assign n25 = n24 ^ n17 ;
  assign n26 = x2 & n25 ;
  assign n27 = ~n16 & ~n26 ;
  assign n28 = n9 & ~n27 ;
  assign n29 = x4 & ~x6 ;
  assign n30 = ~x0 & ~x7 ;
  assign n31 = n29 & n30 ;
  assign n32 = x0 & x6 ;
  assign n33 = n12 & n32 ;
  assign n34 = ~n31 & ~n33 ;
  assign n35 = x1 & x5 ;
  assign n36 = ~n34 & n35 ;
  assign n37 = ~x3 & ~n36 ;
  assign n38 = ~n28 & n37 ;
  assign n53 = x0 & x7 ;
  assign n54 = ~x4 & x5 ;
  assign n55 = ~x1 & ~n29 ;
  assign n56 = ~n22 & ~n55 ;
  assign n57 = ~n54 & ~n56 ;
  assign n58 = n53 & ~n57 ;
  assign n39 = x6 ^ x5 ;
  assign n40 = n39 ^ x0 ;
  assign n41 = n40 ^ x7 ;
  assign n42 = n41 ^ x4 ;
  assign n43 = x6 ^ x4 ;
  assign n44 = x0 & ~n43 ;
  assign n45 = x7 ^ x4 ;
  assign n46 = n41 & ~n45 ;
  assign n47 = n46 ^ n42 ;
  assign n48 = n44 & ~n47 ;
  assign n49 = n48 ^ n46 ;
  assign n50 = ~n42 & n49 ;
  assign n51 = n50 ^ n46 ;
  assign n52 = ~x1 & n51 ;
  assign n59 = n58 ^ n52 ;
  assign n60 = n59 ^ x2 ;
  assign n67 = n60 ^ n59 ;
  assign n61 = n60 ^ x1 ;
  assign n62 = n61 ^ n59 ;
  assign n63 = n60 ^ n52 ;
  assign n64 = n63 ^ x1 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = ~n62 & n65 ;
  assign n68 = n67 ^ n66 ;
  assign n69 = n68 ^ n62 ;
  assign n70 = x5 & ~x7 ;
  assign n71 = n43 ^ x6 ;
  assign n72 = x6 ^ x0 ;
  assign n73 = ~n71 & n72 ;
  assign n74 = n73 ^ x6 ;
  assign n75 = n70 & ~n74 ;
  assign n76 = n75 ^ n59 ;
  assign n77 = n66 ^ n62 ;
  assign n78 = n76 & ~n77 ;
  assign n79 = n78 ^ n59 ;
  assign n80 = ~n69 & n79 ;
  assign n81 = n80 ^ n59 ;
  assign n82 = n81 ^ n58 ;
  assign n83 = n82 ^ n59 ;
  assign n84 = n38 & ~n83 ;
  assign n85 = ~x1 & x4 ;
  assign n86 = x0 & ~n85 ;
  assign n87 = x2 & ~n86 ;
  assign n88 = ~x5 & x6 ;
  assign n89 = ~x2 & ~n30 ;
  assign n90 = ~n85 & ~n89 ;
  assign n91 = n90 ^ x1 ;
  assign n92 = n91 ^ n88 ;
  assign n93 = x2 & ~x4 ;
  assign n94 = x2 & x7 ;
  assign n95 = ~n93 & ~n94 ;
  assign n96 = n95 ^ n53 ;
  assign n97 = ~x1 & ~n96 ;
  assign n98 = n97 ^ n95 ;
  assign n99 = ~n92 & n98 ;
  assign n100 = n99 ^ n97 ;
  assign n101 = n100 ^ n95 ;
  assign n102 = n101 ^ x1 ;
  assign n103 = n88 & ~n102 ;
  assign n104 = ~n87 & n103 ;
  assign n105 = ~x1 & x2 ;
  assign n106 = ~x4 & ~x5 ;
  assign n107 = n9 & n106 ;
  assign n108 = ~n105 & n107 ;
  assign n109 = ~x2 & ~n85 ;
  assign n110 = n70 ^ x1 ;
  assign n111 = n110 ^ n70 ;
  assign n112 = x4 & ~x5 ;
  assign n113 = x7 & n112 ;
  assign n114 = n113 ^ n70 ;
  assign n115 = n111 & n114 ;
  assign n116 = n115 ^ n70 ;
  assign n117 = n109 & n116 ;
  assign n118 = n117 ^ n95 ;
  assign n119 = n118 ^ x0 ;
  assign n128 = n119 ^ n118 ;
  assign n120 = ~n30 & ~n112 ;
  assign n121 = ~x1 & ~n120 ;
  assign n122 = n121 ^ n119 ;
  assign n123 = n122 ^ n118 ;
  assign n124 = n119 ^ n117 ;
  assign n125 = n124 ^ n121 ;
  assign n126 = n125 ^ n123 ;
  assign n127 = ~n123 & n126 ;
  assign n129 = n128 ^ n127 ;
  assign n130 = n129 ^ n123 ;
  assign n131 = ~x4 & x7 ;
  assign n132 = x5 & ~n131 ;
  assign n133 = n132 ^ n118 ;
  assign n134 = n127 ^ n123 ;
  assign n135 = n133 & ~n134 ;
  assign n136 = n135 ^ n118 ;
  assign n137 = ~n130 & ~n136 ;
  assign n138 = n137 ^ n118 ;
  assign n139 = n138 ^ n95 ;
  assign n140 = n139 ^ n118 ;
  assign n141 = ~n108 & n140 ;
  assign n142 = ~x6 & ~n141 ;
  assign n143 = x3 & ~n142 ;
  assign n144 = ~n104 & n143 ;
  assign n145 = ~n84 & ~n144 ;
  assign n146 = ~x1 & n53 ;
  assign n147 = ~x2 & x4 ;
  assign n148 = n147 ^ n93 ;
  assign n149 = x5 & n148 ;
  assign n150 = n149 ^ n93 ;
  assign n151 = n146 & n150 ;
  assign n152 = ~x6 & n151 ;
  assign n153 = ~n145 & ~n152 ;
  assign y0 = ~n153 ;
endmodule
