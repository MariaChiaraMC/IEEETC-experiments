module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 ;
  assign n20 = x5 ^ x4 ;
  assign n16 = x5 ^ x3 ;
  assign n17 = n16 ^ x4 ;
  assign n18 = n17 ^ x6 ;
  assign n19 = n18 ^ x6 ;
  assign n21 = n20 ^ n19 ;
  assign n29 = n21 ^ n18 ;
  assign n30 = n29 ^ n20 ;
  assign n31 = n30 ^ n20 ;
  assign n23 = n18 ^ x5 ;
  assign n32 = n23 ^ n18 ;
  assign n33 = n32 ^ n20 ;
  assign n34 = ~n31 & ~n33 ;
  assign n22 = n18 ^ x2 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ n18 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = n26 ^ n20 ;
  assign n28 = n21 & n27 ;
  assign n35 = n34 ^ n28 ;
  assign n36 = n35 ^ n21 ;
  assign n37 = n28 ^ n20 ;
  assign n38 = n37 ^ n30 ;
  assign n39 = n20 & ~n38 ;
  assign n40 = n39 ^ n28 ;
  assign n41 = n36 & n40 ;
  assign n42 = n41 ^ n34 ;
  assign n43 = n42 ^ n39 ;
  assign n44 = n43 ^ n21 ;
  assign n45 = n44 ^ n20 ;
  assign n46 = n45 ^ n30 ;
  assign n47 = n46 ^ n16 ;
  assign n48 = x1 & n47 ;
  assign n49 = x6 & ~x11 ;
  assign n50 = ~x1 & ~x4 ;
  assign n51 = ~n49 & n50 ;
  assign n52 = x4 & x6 ;
  assign n53 = x5 & n52 ;
  assign n54 = ~x8 & ~x10 ;
  assign n55 = x2 & ~x14 ;
  assign n56 = n54 & n55 ;
  assign n57 = ~x7 & ~x9 ;
  assign n58 = ~x12 & ~x13 ;
  assign n59 = ~n57 & n58 ;
  assign n60 = n56 & n59 ;
  assign n61 = n53 & n60 ;
  assign n62 = ~x2 & ~x5 ;
  assign n63 = ~x1 & n62 ;
  assign n64 = ~n61 & ~n63 ;
  assign n65 = ~n51 & n64 ;
  assign n66 = x3 & ~n65 ;
  assign n67 = ~x3 & x4 ;
  assign n68 = ~n53 & ~n67 ;
  assign n69 = ~x1 & ~n68 ;
  assign n70 = x5 ^ x2 ;
  assign n71 = n50 & n70 ;
  assign n72 = ~x3 & x6 ;
  assign n73 = ~x2 & n72 ;
  assign n74 = n73 ^ n69 ;
  assign n75 = n71 & ~n74 ;
  assign n76 = n75 ^ n73 ;
  assign n77 = ~n69 & n76 ;
  assign n78 = n77 ^ n69 ;
  assign n79 = ~n66 & ~n78 ;
  assign n80 = ~n48 & n79 ;
  assign n81 = ~x0 & ~n80 ;
  assign y0 = n81 ;
endmodule
