module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 ;
  assign n17 = ~x8 & ~x9 ;
  assign n18 = x8 & x9 ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = ~x10 & ~n19 ;
  assign n21 = ~x11 & n20 ;
  assign n22 = x11 ^ x10 ;
  assign n23 = n17 ^ x11 ;
  assign n24 = n22 & n23 ;
  assign n25 = n24 ^ x10 ;
  assign n26 = ~n21 & ~n25 ;
  assign n27 = x7 & n26 ;
  assign n28 = ~x6 & n27 ;
  assign n29 = x7 ^ x4 ;
  assign n30 = x7 ^ x6 ;
  assign n31 = n30 ^ x7 ;
  assign n32 = n31 ^ n29 ;
  assign n34 = ~x10 & ~x11 ;
  assign n33 = ~x10 & x11 ;
  assign n35 = n34 ^ n33 ;
  assign n36 = x7 & n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n32 & n37 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n39 ^ n33 ;
  assign n41 = n40 ^ x7 ;
  assign n42 = n29 & n41 ;
  assign n43 = n42 ^ x4 ;
  assign n44 = ~n28 & n43 ;
  assign n45 = x12 & x13 ;
  assign n46 = x15 & ~n45 ;
  assign n47 = ~n44 & n46 ;
  assign n48 = x10 & ~x11 ;
  assign n49 = ~x6 & ~n34 ;
  assign n50 = n17 & ~n49 ;
  assign n51 = ~n25 & ~n50 ;
  assign n52 = ~n18 & n51 ;
  assign n53 = x15 & ~n52 ;
  assign n54 = ~x12 & n53 ;
  assign n55 = x13 ^ x6 ;
  assign n56 = n55 ^ x6 ;
  assign n57 = n56 ^ x12 ;
  assign n58 = ~x11 & ~n20 ;
  assign n59 = n58 ^ n26 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = x6 & n60 ;
  assign n62 = n61 ^ n26 ;
  assign n63 = n62 ^ x6 ;
  assign n64 = n63 ^ n56 ;
  assign n65 = n64 ^ x12 ;
  assign n66 = ~n57 & n65 ;
  assign n67 = n66 ^ n61 ;
  assign n68 = n67 ^ n26 ;
  assign n69 = n68 ^ n56 ;
  assign n70 = x12 & n69 ;
  assign n71 = n70 ^ x12 ;
  assign n72 = n71 ^ x12 ;
  assign n73 = n72 ^ x12 ;
  assign n74 = ~n54 & ~n73 ;
  assign n75 = ~x13 & ~x15 ;
  assign n76 = x4 & x7 ;
  assign n77 = ~n75 & n76 ;
  assign n78 = ~n74 & n77 ;
  assign n79 = n78 ^ x15 ;
  assign n89 = n79 ^ x15 ;
  assign n90 = n89 ^ x15 ;
  assign n91 = n89 & n90 ;
  assign n81 = x4 & x6 ;
  assign n82 = x12 & n81 ;
  assign n80 = n79 ^ x13 ;
  assign n83 = n82 ^ n80 ;
  assign n84 = n83 ^ n80 ;
  assign n85 = n80 ^ n79 ;
  assign n86 = n85 ^ x15 ;
  assign n87 = n84 & n86 ;
  assign n94 = n91 ^ n87 ;
  assign n88 = n87 ^ n48 ;
  assign n92 = n91 ^ n89 ;
  assign n93 = ~n88 & n92 ;
  assign n95 = n94 ^ n93 ;
  assign n96 = ~n48 & n95 ;
  assign n97 = n96 ^ n87 ;
  assign n98 = n97 ^ n91 ;
  assign n99 = n98 ^ n93 ;
  assign n100 = n99 ^ n78 ;
  assign n101 = ~n47 & ~n100 ;
  assign n102 = x14 & ~n101 ;
  assign n103 = x5 & n102 ;
  assign n104 = x5 & n45 ;
  assign n129 = n19 & n34 ;
  assign n130 = x6 & x7 ;
  assign n131 = ~n129 & n130 ;
  assign n132 = x5 & ~n81 ;
  assign n133 = n132 ^ n45 ;
  assign n134 = x14 & x15 ;
  assign n135 = n134 ^ n132 ;
  assign n136 = n134 ^ x4 ;
  assign n137 = n134 & n136 ;
  assign n138 = n137 ^ n134 ;
  assign n139 = ~n135 & n138 ;
  assign n140 = n139 ^ n137 ;
  assign n141 = n140 ^ n134 ;
  assign n142 = n141 ^ x4 ;
  assign n143 = ~n133 & n142 ;
  assign n144 = n143 ^ n132 ;
  assign n145 = ~n131 & ~n144 ;
  assign n122 = ~x4 & ~x6 ;
  assign n123 = ~x5 & ~n122 ;
  assign n124 = ~x7 & ~n123 ;
  assign n125 = ~x4 & ~n33 ;
  assign n126 = ~n124 & ~n125 ;
  assign n127 = n126 ^ n104 ;
  assign n105 = x6 ^ x4 ;
  assign n106 = n105 ^ n43 ;
  assign n107 = n26 ^ x4 ;
  assign n108 = n107 ^ n26 ;
  assign n109 = x7 & ~x14 ;
  assign n110 = n109 ^ n26 ;
  assign n111 = n108 & n110 ;
  assign n112 = n111 ^ n26 ;
  assign n113 = n112 ^ n105 ;
  assign n114 = ~n106 & ~n113 ;
  assign n115 = n114 ^ n111 ;
  assign n116 = n115 ^ n26 ;
  assign n117 = n116 ^ n43 ;
  assign n118 = ~n105 & n117 ;
  assign n119 = n118 ^ n105 ;
  assign n120 = n119 ^ n43 ;
  assign n121 = n120 ^ n104 ;
  assign n128 = n127 ^ n121 ;
  assign n146 = n145 ^ n128 ;
  assign n147 = n146 ^ n128 ;
  assign n148 = n128 ^ n121 ;
  assign n149 = n148 ^ n104 ;
  assign n150 = n147 & n149 ;
  assign n151 = n150 ^ n121 ;
  assign n152 = ~x6 & n121 ;
  assign n153 = n152 ^ n104 ;
  assign n154 = n151 & n153 ;
  assign n155 = n154 ^ n152 ;
  assign n156 = n104 & n155 ;
  assign n157 = n156 ^ n150 ;
  assign n158 = n157 ^ n120 ;
  assign n159 = n158 ^ n121 ;
  assign n160 = ~n103 & ~n159 ;
  assign n161 = ~x0 & ~x3 ;
  assign n162 = ~x1 & n161 ;
  assign n163 = ~x2 & n162 ;
  assign n164 = ~n160 & n163 ;
  assign y0 = n164 ;
endmodule
