module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 ;
  assign n17 = ~x1 & ~x4 ;
  assign n18 = ~x0 & ~x3 ;
  assign n19 = ~x5 & ~x7 ;
  assign n20 = ~x2 & ~n19 ;
  assign n21 = n18 & n20 ;
  assign n22 = n17 & n21 ;
  assign n23 = x6 ^ x5 ;
  assign n24 = ~x10 & ~x11 ;
  assign n25 = ~x6 & ~n24 ;
  assign n26 = n23 & n25 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = n27 ^ x9 ;
  assign n29 = n28 ^ x8 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n30 ^ x7 ;
  assign n32 = x5 & ~x6 ;
  assign n33 = x11 ^ x10 ;
  assign n34 = n32 & n33 ;
  assign n35 = n34 ^ x8 ;
  assign n36 = n34 & ~n35 ;
  assign n37 = n36 ^ n27 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = ~n31 & n38 ;
  assign n40 = n39 ^ n36 ;
  assign n41 = n40 ^ n34 ;
  assign n42 = x7 & n41 ;
  assign n43 = n42 ^ x7 ;
  assign n44 = n22 & ~n43 ;
  assign y0 = n44 ;
endmodule
