module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 ;
  assign n17 = x1 & ~x3 ;
  assign n18 = x4 & x5 ;
  assign n19 = n17 & n18 ;
  assign n20 = x8 ^ x5 ;
  assign n21 = x12 & ~x13 ;
  assign n22 = x10 & ~x11 ;
  assign n23 = ~n21 & ~n22 ;
  assign n24 = x3 & ~n23 ;
  assign n25 = n24 ^ x8 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n26 ^ n20 ;
  assign n28 = x7 ^ x6 ;
  assign n29 = ~x3 & n28 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = n29 & ~n30 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = ~n27 & n33 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = n35 ^ n29 ;
  assign n37 = n20 & n36 ;
  assign n38 = ~x1 & n37 ;
  assign n39 = ~x7 & ~x8 ;
  assign n40 = ~x6 & n39 ;
  assign n41 = ~x10 & n17 ;
  assign n42 = ~n40 & n41 ;
  assign n43 = x11 & x13 ;
  assign n44 = ~x5 & ~n43 ;
  assign n45 = ~x11 & ~x13 ;
  assign n46 = n45 ^ x12 ;
  assign n47 = x8 ^ x7 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = x12 ^ x6 ;
  assign n50 = n49 ^ n45 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = n47 & ~n51 ;
  assign n53 = n52 ^ n47 ;
  assign n54 = n48 & n53 ;
  assign n55 = n54 ^ n52 ;
  assign n56 = n55 ^ n47 ;
  assign n57 = n56 ^ n50 ;
  assign n58 = n46 & ~n57 ;
  assign n59 = n58 ^ n50 ;
  assign n60 = n44 & ~n59 ;
  assign n61 = n42 & n60 ;
  assign n62 = ~n38 & ~n61 ;
  assign n63 = x4 & ~x9 ;
  assign n64 = ~n62 & n63 ;
  assign n65 = ~n19 & ~n64 ;
  assign n66 = x2 & ~n65 ;
  assign n15 = x2 & x3 ;
  assign n67 = ~x5 & n15 ;
  assign n68 = x4 & ~n45 ;
  assign n69 = n67 & n68 ;
  assign n70 = x10 & x12 ;
  assign n71 = ~x8 & x9 ;
  assign n72 = ~n43 & n71 ;
  assign n73 = n70 & n72 ;
  assign n74 = n69 & n73 ;
  assign n75 = x2 & ~n18 ;
  assign n76 = ~x3 & ~n75 ;
  assign n77 = n15 ^ x5 ;
  assign n78 = n77 ^ n15 ;
  assign n79 = n78 ^ n23 ;
  assign n80 = ~x6 & ~x7 ;
  assign n81 = ~x4 & n71 ;
  assign n82 = n80 & n81 ;
  assign n83 = n82 ^ x2 ;
  assign n84 = ~x2 & n83 ;
  assign n85 = n84 ^ n15 ;
  assign n86 = n85 ^ x2 ;
  assign n87 = ~n79 & ~n86 ;
  assign n88 = n87 ^ n84 ;
  assign n89 = n88 ^ x2 ;
  assign n90 = ~n23 & ~n89 ;
  assign n91 = n90 ^ n23 ;
  assign n92 = ~n76 & ~n91 ;
  assign n93 = ~n74 & ~n92 ;
  assign n94 = ~x2 & ~x9 ;
  assign n95 = ~x3 & x8 ;
  assign n96 = x8 & ~n80 ;
  assign n97 = n24 & ~n96 ;
  assign n98 = x6 & x7 ;
  assign n99 = ~n40 & ~n98 ;
  assign n100 = n97 & n99 ;
  assign n101 = ~n95 & ~n100 ;
  assign n102 = x5 & ~n101 ;
  assign n103 = n102 ^ x4 ;
  assign n104 = n103 ^ n102 ;
  assign n105 = x5 & ~n23 ;
  assign n106 = ~x8 & n105 ;
  assign n107 = n106 ^ x5 ;
  assign n108 = n107 ^ n106 ;
  assign n109 = n106 ^ x8 ;
  assign n110 = n109 ^ n106 ;
  assign n111 = ~n108 & n110 ;
  assign n112 = n111 ^ n106 ;
  assign n113 = ~x3 & n112 ;
  assign n114 = n113 ^ n106 ;
  assign n115 = n114 ^ n102 ;
  assign n116 = n104 & n115 ;
  assign n117 = n116 ^ n102 ;
  assign n118 = n94 & n117 ;
  assign n119 = n93 & ~n118 ;
  assign n120 = ~x1 & ~n119 ;
  assign n121 = ~n66 & ~n120 ;
  assign n16 = ~x1 & n15 ;
  assign n122 = n121 ^ n16 ;
  assign n123 = x0 & ~n122 ;
  assign n124 = n123 ^ n121 ;
  assign y0 = ~n124 ;
endmodule
