module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 ;
  assign n11 = x1 & ~x2 ;
  assign n12 = ~x0 & n11 ;
  assign n13 = x5 & n12 ;
  assign n14 = x8 ^ x4 ;
  assign n15 = n14 ^ x9 ;
  assign n16 = x9 ^ x6 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = x9 ^ x8 ;
  assign n19 = n18 ^ x8 ;
  assign n20 = x8 ^ x3 ;
  assign n21 = n20 ^ x8 ;
  assign n22 = ~n19 & ~n21 ;
  assign n23 = n22 ^ x8 ;
  assign n24 = n23 ^ n15 ;
  assign n25 = n17 & n24 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = n26 ^ x8 ;
  assign n28 = n27 ^ n16 ;
  assign n29 = n15 & n28 ;
  assign n30 = n29 ^ n15 ;
  assign n31 = n13 & n30 ;
  assign n32 = x4 & x6 ;
  assign n33 = ~x5 & ~x9 ;
  assign n34 = n32 & n33 ;
  assign n35 = ~x1 & ~x2 ;
  assign n36 = x0 & x8 ;
  assign n37 = n35 & n36 ;
  assign n38 = n34 & n37 ;
  assign n39 = ~x2 & ~x4 ;
  assign n40 = n33 & n39 ;
  assign n41 = ~x4 & x9 ;
  assign n42 = n35 & n41 ;
  assign n43 = x5 & x9 ;
  assign n44 = n35 & n43 ;
  assign n45 = ~n42 & ~n44 ;
  assign n46 = x1 & x4 ;
  assign n47 = x5 & n46 ;
  assign n48 = n47 ^ x1 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = x4 & ~x5 ;
  assign n51 = x2 & n50 ;
  assign n52 = n51 ^ n47 ;
  assign n53 = n52 ^ n47 ;
  assign n54 = ~n49 & n53 ;
  assign n55 = n54 ^ n47 ;
  assign n56 = x9 & n55 ;
  assign n57 = n56 ^ n47 ;
  assign n58 = n45 & ~n57 ;
  assign n59 = ~n40 & n58 ;
  assign n60 = x0 & ~x6 ;
  assign n61 = ~n59 & n60 ;
  assign n62 = x5 & x6 ;
  assign n63 = ~x1 & x9 ;
  assign n64 = ~x0 & ~n63 ;
  assign n65 = ~n11 & ~n39 ;
  assign n66 = x9 ^ x4 ;
  assign n67 = x1 & ~n66 ;
  assign n68 = n65 & ~n67 ;
  assign n69 = n64 & n68 ;
  assign n70 = ~n42 & ~n69 ;
  assign n71 = n62 & ~n70 ;
  assign n72 = x8 & ~n71 ;
  assign n73 = ~n61 & n72 ;
  assign n74 = ~x4 & ~x6 ;
  assign n75 = n13 & n74 ;
  assign n76 = ~x5 & n74 ;
  assign n77 = ~x0 & ~x1 ;
  assign n78 = ~x5 & ~n77 ;
  assign n79 = n32 & ~n78 ;
  assign n80 = ~n76 & ~n79 ;
  assign n81 = x2 & ~n80 ;
  assign n82 = ~x1 & x5 ;
  assign n83 = x1 ^ x0 ;
  assign n84 = n82 & ~n83 ;
  assign n85 = n84 ^ n83 ;
  assign n86 = n81 & ~n85 ;
  assign n87 = ~n75 & ~n86 ;
  assign n88 = n87 ^ x9 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = x2 & ~x6 ;
  assign n91 = ~x4 & x5 ;
  assign n92 = n77 & n91 ;
  assign n93 = n90 & n92 ;
  assign n94 = x0 & x1 ;
  assign n95 = ~x5 & n94 ;
  assign n96 = n32 & n95 ;
  assign n97 = ~n93 & ~n96 ;
  assign n98 = n97 ^ n87 ;
  assign n99 = ~n89 & n98 ;
  assign n100 = n99 ^ n87 ;
  assign n101 = ~x8 & n100 ;
  assign n102 = ~n73 & ~n101 ;
  assign n103 = n102 ^ x3 ;
  assign n104 = n103 ^ n102 ;
  assign n105 = ~x4 & ~x9 ;
  assign n106 = x2 & ~x8 ;
  assign n107 = n105 & n106 ;
  assign n108 = x0 & ~x2 ;
  assign n109 = ~x8 & x9 ;
  assign n110 = n109 ^ x1 ;
  assign n111 = n110 ^ n109 ;
  assign n112 = x8 & ~x9 ;
  assign n113 = n112 ^ n109 ;
  assign n114 = n113 ^ n109 ;
  assign n115 = ~n111 & n114 ;
  assign n116 = n115 ^ n109 ;
  assign n117 = ~x4 & n116 ;
  assign n118 = n117 ^ n109 ;
  assign n119 = n108 & n118 ;
  assign n120 = x4 & x9 ;
  assign n121 = ~n106 & ~n120 ;
  assign n122 = x2 & x4 ;
  assign n123 = x0 & ~n122 ;
  assign n124 = ~n121 & n123 ;
  assign n125 = ~x0 & ~n41 ;
  assign n126 = x2 & n125 ;
  assign n127 = ~n109 & n126 ;
  assign n128 = ~n124 & ~n127 ;
  assign n129 = x1 & ~n128 ;
  assign n130 = ~n119 & ~n129 ;
  assign n131 = ~n107 & n130 ;
  assign n132 = n62 & ~n131 ;
  assign n158 = x2 ^ x1 ;
  assign n159 = ~x5 & n158 ;
  assign n147 = ~x1 & ~x4 ;
  assign n148 = x2 & x8 ;
  assign n149 = n147 & n148 ;
  assign n133 = x5 ^ x4 ;
  assign n134 = n133 ^ x8 ;
  assign n135 = x8 ^ x1 ;
  assign n136 = n135 ^ x2 ;
  assign n137 = n136 ^ n134 ;
  assign n138 = x5 ^ x2 ;
  assign n139 = n138 ^ x8 ;
  assign n140 = x8 & n139 ;
  assign n141 = n140 ^ x2 ;
  assign n142 = n141 ^ x8 ;
  assign n143 = n137 & ~n142 ;
  assign n144 = n143 ^ n140 ;
  assign n145 = n144 ^ x8 ;
  assign n146 = n134 & n145 ;
  assign n150 = n149 ^ n146 ;
  assign n151 = n150 ^ n146 ;
  assign n152 = n146 ^ x5 ;
  assign n153 = n152 ^ n146 ;
  assign n154 = n151 & n153 ;
  assign n155 = n154 ^ n146 ;
  assign n156 = x9 & n155 ;
  assign n157 = n156 ^ n146 ;
  assign n160 = n159 ^ n157 ;
  assign n161 = n160 ^ x0 ;
  assign n170 = n161 ^ n160 ;
  assign n162 = ~x2 & n105 ;
  assign n163 = ~x8 & n162 ;
  assign n164 = n163 ^ n161 ;
  assign n165 = n164 ^ n160 ;
  assign n166 = n163 ^ n159 ;
  assign n167 = n166 ^ n163 ;
  assign n168 = n167 ^ n165 ;
  assign n169 = n165 & n168 ;
  assign n171 = n170 ^ n169 ;
  assign n172 = n171 ^ n165 ;
  assign n173 = n160 ^ n109 ;
  assign n174 = n169 ^ n165 ;
  assign n175 = ~n173 & n174 ;
  assign n176 = n175 ^ n160 ;
  assign n177 = ~n172 & n176 ;
  assign n178 = n177 ^ n160 ;
  assign n179 = n178 ^ n159 ;
  assign n180 = n179 ^ n160 ;
  assign n181 = ~x6 & n180 ;
  assign n182 = ~x5 & x6 ;
  assign n183 = n148 & n182 ;
  assign n184 = n67 & n183 ;
  assign n185 = n147 ^ n109 ;
  assign n186 = n185 ^ n109 ;
  assign n187 = x5 & x8 ;
  assign n188 = ~n46 & n187 ;
  assign n189 = n188 ^ n109 ;
  assign n190 = ~n186 & n189 ;
  assign n191 = n190 ^ n109 ;
  assign n192 = n90 & n191 ;
  assign n193 = ~n184 & ~n192 ;
  assign n194 = x0 & ~n193 ;
  assign n195 = ~n181 & ~n194 ;
  assign n196 = ~n132 & n195 ;
  assign n197 = n196 ^ n102 ;
  assign n198 = n104 & ~n197 ;
  assign n199 = n198 ^ n102 ;
  assign n200 = ~n38 & ~n199 ;
  assign n201 = n200 ^ x7 ;
  assign n202 = n201 ^ n200 ;
  assign n205 = ~x2 & ~x6 ;
  assign n206 = x4 ^ x3 ;
  assign n207 = ~n205 & ~n206 ;
  assign n203 = ~x6 & x9 ;
  assign n208 = n207 ^ n203 ;
  assign n204 = n203 ^ x2 ;
  assign n209 = n208 ^ n204 ;
  assign n210 = n209 ^ n208 ;
  assign n211 = n210 ^ n203 ;
  assign n212 = x3 & ~x6 ;
  assign n213 = n212 ^ n209 ;
  assign n214 = n41 & n213 ;
  assign n215 = n208 ^ n203 ;
  assign n216 = n210 & n215 ;
  assign n217 = n216 ^ n211 ;
  assign n218 = n214 & ~n217 ;
  assign n219 = n218 ^ n216 ;
  assign n220 = ~n211 & n219 ;
  assign n221 = n220 ^ n216 ;
  assign n222 = n221 ^ n207 ;
  assign n223 = n82 & n222 ;
  assign n224 = x2 & ~x9 ;
  assign n225 = x3 & x4 ;
  assign n226 = n182 & n225 ;
  assign n227 = n224 & n226 ;
  assign n228 = ~n223 & ~n227 ;
  assign n229 = ~x8 & ~n228 ;
  assign n230 = x0 & n229 ;
  assign n238 = ~x3 & x6 ;
  assign n236 = ~x8 & ~n212 ;
  assign n237 = n122 & ~n236 ;
  assign n239 = n238 ^ n237 ;
  assign n240 = n239 ^ n237 ;
  assign n241 = n237 ^ x8 ;
  assign n242 = ~n240 & ~n241 ;
  assign n243 = n242 ^ n237 ;
  assign n244 = ~n39 & ~n237 ;
  assign n245 = n244 ^ x9 ;
  assign n246 = ~n243 & n245 ;
  assign n247 = n246 ^ n244 ;
  assign n248 = x9 & n247 ;
  assign n249 = n248 ^ x9 ;
  assign n250 = ~x3 & ~n39 ;
  assign n251 = n250 ^ n112 ;
  assign n252 = n74 ^ x2 ;
  assign n253 = n252 ^ n74 ;
  assign n254 = n74 ^ x6 ;
  assign n255 = ~n253 & n254 ;
  assign n256 = n255 ^ n74 ;
  assign n257 = n256 ^ n250 ;
  assign n258 = n251 & n257 ;
  assign n259 = n258 ^ n255 ;
  assign n260 = n259 ^ n74 ;
  assign n261 = n260 ^ n112 ;
  assign n262 = n250 & n261 ;
  assign n263 = n262 ^ n250 ;
  assign n264 = ~n249 & ~n263 ;
  assign n231 = ~x3 & x4 ;
  assign n232 = ~x2 & n231 ;
  assign n233 = n109 & n232 ;
  assign n234 = n105 & n148 ;
  assign n235 = ~n233 & ~n234 ;
  assign n265 = n264 ^ n235 ;
  assign n266 = n265 ^ n264 ;
  assign n267 = n264 ^ x6 ;
  assign n268 = n267 ^ n264 ;
  assign n269 = ~n266 & n268 ;
  assign n270 = n269 ^ n264 ;
  assign n271 = x5 & ~n270 ;
  assign n272 = n271 ^ n264 ;
  assign n273 = n94 & ~n272 ;
  assign n274 = ~n230 & ~n273 ;
  assign n275 = n76 & n224 ;
  assign n276 = n275 ^ n43 ;
  assign n277 = n276 ^ x1 ;
  assign n285 = n277 ^ n276 ;
  assign n278 = ~x4 & n158 ;
  assign n279 = n278 ^ n277 ;
  assign n280 = n279 ^ n276 ;
  assign n281 = n277 ^ n275 ;
  assign n282 = n281 ^ n278 ;
  assign n283 = n282 ^ n280 ;
  assign n284 = n280 & ~n283 ;
  assign n286 = n285 ^ n284 ;
  assign n287 = n286 ^ n280 ;
  assign n288 = n276 ^ x6 ;
  assign n289 = n284 ^ n280 ;
  assign n290 = n288 & n289 ;
  assign n291 = n290 ^ n276 ;
  assign n292 = ~n287 & n291 ;
  assign n293 = n292 ^ n276 ;
  assign n294 = n293 ^ n43 ;
  assign n295 = n294 ^ n276 ;
  assign n296 = ~x3 & n295 ;
  assign n297 = x6 & ~n33 ;
  assign n298 = n225 & n297 ;
  assign n299 = n35 & n298 ;
  assign n300 = ~n296 & ~n299 ;
  assign n301 = n300 ^ x8 ;
  assign n302 = n301 ^ n300 ;
  assign n303 = n203 & n232 ;
  assign n304 = x5 & ~n224 ;
  assign n305 = ~x3 & ~x4 ;
  assign n306 = n297 & n305 ;
  assign n307 = ~n304 & n306 ;
  assign n308 = ~x2 & x3 ;
  assign n309 = n43 & n74 ;
  assign n310 = ~n34 & ~n309 ;
  assign n311 = n308 & ~n310 ;
  assign n312 = ~n307 & ~n311 ;
  assign n313 = ~n303 & n312 ;
  assign n314 = x1 & ~n313 ;
  assign n315 = ~x3 & ~x5 ;
  assign n318 = x6 & ~x9 ;
  assign n316 = x5 & ~n231 ;
  assign n317 = n203 & ~n316 ;
  assign n319 = n318 ^ n317 ;
  assign n320 = ~n315 & n319 ;
  assign n321 = n320 ^ n318 ;
  assign n322 = x1 & ~n308 ;
  assign n323 = n50 ^ x2 ;
  assign n324 = ~n322 & n323 ;
  assign n325 = n321 & n324 ;
  assign n326 = ~n314 & ~n325 ;
  assign n327 = n326 ^ n300 ;
  assign n328 = ~n302 & n327 ;
  assign n329 = n328 ^ n300 ;
  assign n330 = ~x0 & ~n329 ;
  assign n331 = n274 & ~n330 ;
  assign n332 = n331 ^ n200 ;
  assign n333 = ~n202 & n332 ;
  assign n334 = n333 ^ n200 ;
  assign n335 = ~n31 & n334 ;
  assign y0 = ~n335 ;
endmodule
