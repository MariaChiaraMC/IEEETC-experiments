module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 ;
  assign n9 = ~x2 & ~x3 ;
  assign n10 = x6 & x7 ;
  assign n11 = ~n9 & ~n10 ;
  assign n12 = ~x6 & ~x7 ;
  assign n15 = ~x5 & n12 ;
  assign n16 = x4 & ~n15 ;
  assign n13 = x5 & ~n12 ;
  assign n14 = ~x2 & ~n13 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = n14 ^ x3 ;
  assign n20 = ~n18 & ~n19 ;
  assign n21 = n20 ^ n14 ;
  assign n22 = n11 & n21 ;
  assign n23 = x1 & ~n22 ;
  assign n24 = x4 ^ x1 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = x5 ^ x4 ;
  assign n27 = n26 ^ x4 ;
  assign n28 = ~n25 & n27 ;
  assign n29 = n28 ^ x4 ;
  assign n30 = x7 & ~n29 ;
  assign n31 = n30 ^ x4 ;
  assign n32 = ~x6 & ~n31 ;
  assign n33 = ~x0 & ~n32 ;
  assign n34 = ~x5 & x6 ;
  assign n35 = n34 ^ x1 ;
  assign n36 = n34 ^ x4 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = ~x4 & ~x7 ;
  assign n41 = x2 & n40 ;
  assign n42 = n41 ^ x3 ;
  assign n43 = n42 ^ n41 ;
  assign n48 = n41 ^ n36 ;
  assign n44 = n38 ^ n36 ;
  assign n45 = n44 ^ n35 ;
  assign n46 = n36 ^ x2 ;
  assign n47 = n45 & n46 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = n49 ^ n36 ;
  assign n51 = ~n43 & n50 ;
  assign n52 = n51 ^ n48 ;
  assign n53 = n52 ^ n38 ;
  assign n54 = n39 & ~n53 ;
  assign n55 = n54 ^ n51 ;
  assign n56 = n55 ^ n48 ;
  assign n57 = n56 ^ n36 ;
  assign n58 = ~n35 & n57 ;
  assign n59 = n58 ^ x1 ;
  assign n60 = n33 & n59 ;
  assign n61 = ~n23 & n60 ;
  assign n62 = ~x1 & ~x4 ;
  assign n63 = x0 & ~x5 ;
  assign n64 = n9 & n63 ;
  assign n65 = n62 & n64 ;
  assign n66 = n10 & n65 ;
  assign n67 = ~n61 & ~n66 ;
  assign y0 = ~n67 ;
endmodule
