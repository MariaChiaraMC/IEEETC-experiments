module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n10 = ~x6 & x7 ;
  assign n11 = x4 & ~x8 ;
  assign n12 = n11 ^ x2 ;
  assign n13 = n12 ^ n10 ;
  assign n14 = n11 ^ x5 ;
  assign n15 = n14 ^ x5 ;
  assign n16 = x5 ^ x3 ;
  assign n17 = ~n15 & ~n16 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = n18 ^ n10 ;
  assign n20 = ~n13 & n19 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n21 ^ x5 ;
  assign n23 = n22 ^ n12 ;
  assign n24 = n10 & ~n23 ;
  assign n25 = n24 ^ n10 ;
  assign n26 = n25 ^ n12 ;
  assign n27 = ~x0 & ~n26 ;
  assign n28 = x4 & ~x5 ;
  assign n29 = n28 ^ x1 ;
  assign n30 = x8 & n10 ;
  assign n31 = n30 ^ x1 ;
  assign n32 = n31 ^ x1 ;
  assign n33 = ~n29 & n32 ;
  assign n34 = n33 ^ x1 ;
  assign n35 = x3 & n34 ;
  assign n36 = n35 ^ x1 ;
  assign n37 = n27 & n36 ;
  assign y0 = n37 ;
endmodule
