module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 ;
  assign n9 = x4 ^ x1 ;
  assign n10 = n9 ^ x4 ;
  assign n11 = n10 ^ x5 ;
  assign n12 = n11 ^ x6 ;
  assign n13 = n12 ^ x7 ;
  assign n14 = n13 ^ x3 ;
  assign n27 = n14 ^ n9 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n15 ^ n9 ;
  assign n17 = n16 ^ x3 ;
  assign n28 = n27 ^ n17 ;
  assign n21 = n9 ^ x6 ;
  assign n19 = n12 ^ x5 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n23 ^ n12 ;
  assign n25 = n24 ^ n9 ;
  assign n31 = n28 ^ n25 ;
  assign n32 = n17 ^ n14 ;
  assign n33 = n32 ^ x3 ;
  assign n34 = n33 ^ n25 ;
  assign n35 = ~n31 & n34 ;
  assign n18 = n17 ^ x3 ;
  assign n20 = n19 ^ x3 ;
  assign n26 = n25 ^ n20 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = n18 & n29 ;
  assign n36 = n35 ^ n30 ;
  assign n37 = n36 ^ n17 ;
  assign n38 = n37 ^ n19 ;
  assign n39 = n38 ^ n28 ;
  assign n40 = n25 ^ n19 ;
  assign n41 = n25 & ~n40 ;
  assign n42 = n41 ^ x3 ;
  assign n43 = n42 ^ n19 ;
  assign n44 = n35 ^ n14 ;
  assign n45 = n44 ^ n17 ;
  assign n46 = n45 ^ x3 ;
  assign n47 = n46 ^ n25 ;
  assign n48 = n47 ^ n28 ;
  assign n49 = ~n43 & ~n48 ;
  assign n50 = n49 ^ n19 ;
  assign n51 = n39 & ~n50 ;
  assign n52 = n51 ^ n35 ;
  assign n53 = n52 ^ n41 ;
  assign n54 = n53 ^ n30 ;
  assign n55 = n54 ^ n49 ;
  assign n56 = n55 ^ n17 ;
  assign n57 = n56 ^ n28 ;
  assign n58 = ~x2 & n57 ;
  assign n59 = x3 ^ x2 ;
  assign n60 = x5 & x7 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = x5 & x6 ;
  assign n63 = ~x4 & ~n62 ;
  assign n64 = n63 ^ x2 ;
  assign n65 = n64 ^ n63 ;
  assign n66 = ~x4 & x5 ;
  assign n67 = n66 ^ n63 ;
  assign n68 = ~n65 & ~n67 ;
  assign n69 = n68 ^ n63 ;
  assign n70 = n69 ^ n59 ;
  assign n71 = ~n61 & n70 ;
  assign n72 = n71 ^ n68 ;
  assign n73 = n72 ^ n63 ;
  assign n74 = n73 ^ n60 ;
  assign n75 = n59 & ~n74 ;
  assign n76 = n75 ^ n59 ;
  assign n77 = n76 ^ x3 ;
  assign n78 = ~x1 & n77 ;
  assign n79 = ~n58 & ~n78 ;
  assign n80 = ~x0 & ~n79 ;
  assign y0 = n80 ;
endmodule
