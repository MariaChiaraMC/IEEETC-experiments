module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 ;
  assign n16 = x2 ^ x1 ;
  assign n17 = n16 ^ x3 ;
  assign n19 = n17 ^ x3 ;
  assign n18 = n17 ^ x2 ;
  assign n20 = n19 ^ n18 ;
  assign n25 = n20 ^ n17 ;
  assign n26 = n25 ^ n19 ;
  assign n27 = n26 ^ n19 ;
  assign n28 = x5 & x6 ;
  assign n29 = n28 ^ n17 ;
  assign n30 = n29 ^ n17 ;
  assign n31 = n30 ^ n19 ;
  assign n32 = n27 & ~n31 ;
  assign n21 = n17 ^ x4 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n20 & n23 ;
  assign n33 = n32 ^ n24 ;
  assign n34 = n33 ^ n20 ;
  assign n35 = n24 ^ n19 ;
  assign n36 = n35 ^ n26 ;
  assign n37 = n19 & n36 ;
  assign n38 = n37 ^ n24 ;
  assign n39 = n34 & n38 ;
  assign n40 = n39 ^ n32 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n41 ^ n20 ;
  assign n43 = n42 ^ n19 ;
  assign n44 = n43 ^ n26 ;
  assign n45 = n44 ^ x3 ;
  assign y0 = n45 ;
endmodule
