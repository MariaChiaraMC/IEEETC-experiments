module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 ;
  assign n10 = ~x3 & ~x4 ;
  assign n11 = ~x5 & x8 ;
  assign n12 = ~x2 & ~n11 ;
  assign n13 = ~n10 & ~n12 ;
  assign n14 = ~x3 & ~x6 ;
  assign n15 = x7 & ~n14 ;
  assign n16 = x0 & n15 ;
  assign n17 = n13 & n16 ;
  assign n18 = x3 & x6 ;
  assign n19 = x3 & x4 ;
  assign n20 = ~n18 & ~n19 ;
  assign n21 = x2 & ~x3 ;
  assign n22 = x5 & ~x8 ;
  assign n23 = x2 & ~n22 ;
  assign n24 = ~n21 & ~n23 ;
  assign n25 = n20 & n24 ;
  assign n26 = n17 & n25 ;
  assign n56 = ~x7 & ~x8 ;
  assign n57 = x5 ^ x3 ;
  assign n58 = x6 ^ x5 ;
  assign n59 = x3 ^ x2 ;
  assign n60 = n59 ^ x6 ;
  assign n61 = x6 & n60 ;
  assign n62 = n61 ^ x6 ;
  assign n63 = n58 & n62 ;
  assign n64 = n63 ^ n61 ;
  assign n65 = n64 ^ x6 ;
  assign n66 = n65 ^ n59 ;
  assign n67 = ~n57 & n66 ;
  assign n68 = n67 ^ n59 ;
  assign n69 = n56 & n68 ;
  assign n44 = ~x6 & x7 ;
  assign n70 = ~x2 & ~x3 ;
  assign n71 = n44 & n70 ;
  assign n72 = x8 & n71 ;
  assign n73 = x5 & n72 ;
  assign n74 = ~n69 & ~n73 ;
  assign n75 = x2 & x5 ;
  assign n30 = ~x6 & ~x7 ;
  assign n41 = x3 & x8 ;
  assign n76 = n30 & n41 ;
  assign n77 = x7 & ~x8 ;
  assign n78 = n18 & n77 ;
  assign n79 = ~n76 & ~n78 ;
  assign n80 = n75 & ~n79 ;
  assign n81 = ~x0 & ~n80 ;
  assign n82 = n74 & n81 ;
  assign n27 = x6 & x7 ;
  assign n83 = x8 ^ x7 ;
  assign n84 = n83 ^ x7 ;
  assign n85 = x2 & x6 ;
  assign n86 = n85 ^ x7 ;
  assign n87 = n84 & n86 ;
  assign n88 = n87 ^ x7 ;
  assign n89 = x3 & n88 ;
  assign n90 = ~n27 & n89 ;
  assign n91 = n90 ^ x5 ;
  assign n92 = n91 ^ n90 ;
  assign n93 = ~x2 & n77 ;
  assign n94 = x6 ^ x3 ;
  assign n95 = n93 & ~n94 ;
  assign n96 = ~n76 & ~n95 ;
  assign n97 = n96 ^ n90 ;
  assign n98 = ~n92 & ~n97 ;
  assign n99 = n98 ^ n90 ;
  assign n100 = x0 & ~n99 ;
  assign n101 = ~n82 & ~n100 ;
  assign n42 = ~x5 & x7 ;
  assign n43 = ~x2 & n42 ;
  assign n45 = n44 ^ x2 ;
  assign n46 = n45 ^ n44 ;
  assign n47 = n44 ^ n30 ;
  assign n48 = ~n46 & n47 ;
  assign n49 = n48 ^ n44 ;
  assign n50 = x5 & n49 ;
  assign n51 = ~n43 & ~n50 ;
  assign n52 = n41 & ~n51 ;
  assign n28 = ~n11 & ~n27 ;
  assign n29 = n21 & ~n28 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = ~x2 & x5 ;
  assign n33 = ~x8 & n32 ;
  assign n34 = n33 ^ n29 ;
  assign n35 = n34 ^ n33 ;
  assign n36 = n33 ^ n22 ;
  assign n37 = n35 & ~n36 ;
  assign n38 = n37 ^ n33 ;
  assign n39 = n31 & ~n38 ;
  assign n40 = n39 ^ n30 ;
  assign n53 = n52 ^ n40 ;
  assign n54 = ~x0 & n53 ;
  assign n55 = n54 ^ n52 ;
  assign n102 = n101 ^ n55 ;
  assign n103 = n102 ^ n101 ;
  assign n104 = x3 & n27 ;
  assign n105 = n33 & n104 ;
  assign n106 = n105 ^ n101 ;
  assign n107 = n106 ^ n101 ;
  assign n108 = ~n103 & ~n107 ;
  assign n109 = n108 ^ n101 ;
  assign n110 = x4 & ~n109 ;
  assign n111 = n110 ^ n101 ;
  assign n112 = n111 ^ x1 ;
  assign n113 = n112 ^ n111 ;
  assign n122 = ~x4 & ~x7 ;
  assign n123 = x5 & ~n122 ;
  assign n124 = x4 & n27 ;
  assign n125 = n124 ^ x6 ;
  assign n126 = n123 & n125 ;
  assign n127 = n70 & n126 ;
  assign n114 = ~n14 & ~n104 ;
  assign n115 = ~x2 & ~x4 ;
  assign n116 = ~x5 & n115 ;
  assign n117 = ~n114 & n116 ;
  assign n118 = x4 & ~x5 ;
  assign n119 = n21 & n118 ;
  assign n120 = n44 & n119 ;
  assign n121 = ~n117 & ~n120 ;
  assign n128 = n127 ^ n121 ;
  assign n129 = n128 ^ n121 ;
  assign n130 = n43 ^ x4 ;
  assign n131 = n30 ^ n27 ;
  assign n132 = n30 ^ x5 ;
  assign n133 = n132 ^ n30 ;
  assign n134 = n131 & n133 ;
  assign n135 = n134 ^ n30 ;
  assign n136 = n135 ^ n43 ;
  assign n137 = n130 & ~n136 ;
  assign n138 = n137 ^ n134 ;
  assign n139 = n138 ^ n30 ;
  assign n140 = n139 ^ x4 ;
  assign n141 = ~n43 & ~n140 ;
  assign n142 = n141 ^ n43 ;
  assign n143 = n142 ^ n43 ;
  assign n144 = x3 & ~n143 ;
  assign n145 = ~n115 & n144 ;
  assign n146 = n145 ^ n121 ;
  assign n147 = n146 ^ n121 ;
  assign n148 = ~n129 & ~n147 ;
  assign n149 = n148 ^ n121 ;
  assign n150 = x8 & n149 ;
  assign n151 = n150 ^ n121 ;
  assign n152 = ~x0 & n151 ;
  assign n153 = ~x4 & x5 ;
  assign n154 = ~n118 & ~n153 ;
  assign n155 = n71 & ~n154 ;
  assign n156 = n118 ^ x5 ;
  assign n157 = ~x7 & n156 ;
  assign n158 = n157 ^ x5 ;
  assign n159 = n18 & n158 ;
  assign n160 = x2 & n159 ;
  assign n161 = ~n155 & ~n160 ;
  assign n162 = n161 ^ x8 ;
  assign n163 = n162 ^ n161 ;
  assign n164 = n163 ^ x0 ;
  assign n165 = x7 ^ x6 ;
  assign n166 = n70 & ~n165 ;
  assign n167 = n166 ^ n123 ;
  assign n168 = n166 & ~n167 ;
  assign n169 = n168 ^ n161 ;
  assign n170 = n169 ^ n166 ;
  assign n171 = n164 & ~n170 ;
  assign n172 = n171 ^ n168 ;
  assign n173 = n172 ^ n166 ;
  assign n174 = x0 & n173 ;
  assign n175 = n174 ^ x0 ;
  assign n176 = ~n152 & ~n175 ;
  assign n177 = n176 ^ n111 ;
  assign n178 = n113 & n177 ;
  assign n179 = n178 ^ n111 ;
  assign n180 = ~n26 & ~n179 ;
  assign y0 = ~n180 ;
endmodule
