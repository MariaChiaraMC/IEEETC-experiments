module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n9 = ~x6 & x7 ;
  assign n10 = ~x4 & ~x5 ;
  assign n11 = ~x0 & n10 ;
  assign n12 = n9 & n11 ;
  assign n13 = ~x4 & n9 ;
  assign n14 = n13 ^ x1 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = x5 ^ x4 ;
  assign n17 = n16 ^ x6 ;
  assign n18 = x7 ^ x5 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = n19 ^ x7 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = x7 ^ x6 ;
  assign n23 = x7 ^ x2 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n22 & n24 ;
  assign n26 = n25 ^ x7 ;
  assign n27 = n26 ^ n22 ;
  assign n28 = n21 & n27 ;
  assign n29 = n28 ^ n25 ;
  assign n30 = n29 ^ n22 ;
  assign n31 = ~n17 & n30 ;
  assign n32 = n31 ^ n13 ;
  assign n33 = ~n15 & n32 ;
  assign n34 = n33 ^ n13 ;
  assign n35 = x0 & n34 ;
  assign n36 = ~n12 & ~n35 ;
  assign n37 = ~x3 & ~n36 ;
  assign y0 = n37 ;
endmodule
