module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 ;
  assign n10 = x0 & ~x4 ;
  assign n11 = ~x2 & n10 ;
  assign n12 = ~x0 & x1 ;
  assign n13 = x6 & n12 ;
  assign n14 = x3 & n13 ;
  assign n15 = ~n11 & ~n14 ;
  assign n16 = x5 & ~n15 ;
  assign n17 = x2 ^ x0 ;
  assign n18 = x4 ^ x2 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = x5 & x8 ;
  assign n22 = x6 & n21 ;
  assign n23 = n22 ^ x3 ;
  assign n24 = ~x3 & ~n23 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = n25 ^ x3 ;
  assign n27 = n20 & n26 ;
  assign n28 = n27 ^ n24 ;
  assign n29 = n28 ^ x3 ;
  assign n30 = n17 & ~n29 ;
  assign n31 = x7 & n30 ;
  assign n32 = x3 & x4 ;
  assign n33 = ~x2 & ~n32 ;
  assign n34 = n12 & ~n33 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = ~x3 & ~x4 ;
  assign n37 = x2 & ~n36 ;
  assign n38 = x4 & x7 ;
  assign n39 = n22 & n38 ;
  assign n40 = n37 & ~n39 ;
  assign n41 = n40 ^ x0 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = ~x1 & ~n37 ;
  assign n44 = ~x6 & ~x8 ;
  assign n45 = ~x4 & n44 ;
  assign n46 = n33 & ~n45 ;
  assign n47 = ~x7 & ~x8 ;
  assign n48 = n47 ^ x1 ;
  assign n49 = n48 ^ x1 ;
  assign n50 = x2 ^ x1 ;
  assign n51 = n50 ^ x1 ;
  assign n52 = n49 & ~n51 ;
  assign n53 = n52 ^ x1 ;
  assign n54 = x3 & ~n53 ;
  assign n55 = n54 ^ x1 ;
  assign n56 = ~x6 & ~n55 ;
  assign n57 = ~x5 & n56 ;
  assign n58 = ~n46 & ~n57 ;
  assign n59 = ~n43 & n58 ;
  assign n60 = n59 ^ n40 ;
  assign n61 = n42 & ~n60 ;
  assign n62 = n61 ^ n40 ;
  assign n63 = n62 ^ n31 ;
  assign n64 = n35 & n63 ;
  assign n65 = n64 ^ n61 ;
  assign n66 = n65 ^ n40 ;
  assign n67 = n66 ^ n34 ;
  assign n68 = ~n31 & n67 ;
  assign n69 = n68 ^ n31 ;
  assign n70 = ~n16 & ~n69 ;
  assign y0 = ~n70 ;
endmodule
