module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 ;
  assign n15 = x7 & ~x8 ;
  assign n16 = x6 & n15 ;
  assign n17 = ~x10 & ~n16 ;
  assign n18 = ~x4 & ~x10 ;
  assign n19 = x13 & ~n18 ;
  assign n20 = n19 ^ x12 ;
  assign n21 = n20 ^ x11 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n23 ^ n20 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ n20 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n20 ^ x1 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = ~n27 & n29 ;
  assign n31 = n30 ^ n20 ;
  assign n32 = n31 ^ n26 ;
  assign n33 = n32 ^ n24 ;
  assign n34 = ~x3 & ~x9 ;
  assign n35 = x2 & ~n34 ;
  assign n36 = n35 ^ n30 ;
  assign n37 = n36 ^ n20 ;
  assign n38 = n24 & n37 ;
  assign n39 = n38 ^ n26 ;
  assign n40 = n39 ^ n24 ;
  assign n41 = ~n33 & ~n40 ;
  assign n42 = n41 ^ n30 ;
  assign n43 = n42 ^ n20 ;
  assign n44 = n43 ^ n26 ;
  assign n45 = n44 ^ n24 ;
  assign n46 = n45 ^ x12 ;
  assign n47 = ~n17 & ~n46 ;
  assign n48 = x7 ^ x6 ;
  assign n49 = n48 ^ n15 ;
  assign n50 = ~x5 & ~n49 ;
  assign n51 = n50 ^ n15 ;
  assign n52 = ~x4 & n51 ;
  assign n53 = n16 ^ x10 ;
  assign n54 = x11 ^ x10 ;
  assign n55 = n54 ^ x10 ;
  assign n56 = n53 & n55 ;
  assign n57 = n56 ^ x10 ;
  assign n58 = ~x0 & n57 ;
  assign n59 = ~n52 & ~n58 ;
  assign n60 = x12 & ~n59 ;
  assign n61 = ~n47 & ~n60 ;
  assign y0 = ~n61 ;
endmodule
