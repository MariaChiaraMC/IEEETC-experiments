module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 ;
  assign n7 = x2 ^ x0 ;
  assign n10 = n7 ^ x5 ;
  assign n11 = n10 ^ n7 ;
  assign n8 = n7 ^ x4 ;
  assign n9 = n8 ^ n7 ;
  assign n12 = n11 ^ n9 ;
  assign n13 = n7 ^ x0 ;
  assign n14 = n13 ^ n7 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = n11 & n15 ;
  assign n17 = n16 ^ n11 ;
  assign n18 = ~n12 & n17 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n19 ^ n7 ;
  assign n21 = n20 ^ n11 ;
  assign n22 = ~x1 & ~n21 ;
  assign n23 = n22 ^ n7 ;
  assign n24 = x3 & ~n23 ;
  assign n25 = ~x1 & ~x3 ;
  assign n26 = ~x2 & ~x5 ;
  assign n27 = x4 & ~n26 ;
  assign n28 = ~n7 & n27 ;
  assign n29 = ~n25 & n28 ;
  assign n30 = ~n24 & ~n29 ;
  assign n31 = x3 ^ x1 ;
  assign n32 = n27 ^ x3 ;
  assign n33 = n32 ^ n27 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = ~x0 & x4 ;
  assign n36 = n35 ^ x5 ;
  assign n37 = ~n35 & n36 ;
  assign n38 = n37 ^ n27 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n34 & ~n39 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n41 ^ n35 ;
  assign n43 = n31 & ~n42 ;
  assign n44 = n43 ^ x3 ;
  assign n45 = n7 & ~n44 ;
  assign n46 = n30 & ~n45 ;
  assign y0 = ~n46 ;
endmodule
