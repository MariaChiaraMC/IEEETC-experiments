// Benchmark "./dekoder.pla" written by ABC on Thu Apr 23 10:59:49 2020

module \./dekoder.pla  ( 
    x0, x1, x2, x3,
    z4  );
  input  x0, x1, x2, x3;
  output z4;
  assign z4 = ~x1 | x2;
endmodule


