module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 ;
  assign n17 = x12 & x13 ;
  assign n18 = ~x12 & ~x13 ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = ~x8 & ~x9 ;
  assign n21 = x10 & x11 ;
  assign n22 = n20 & n21 ;
  assign n23 = ~x10 & ~x11 ;
  assign n24 = x8 & x9 ;
  assign n25 = n23 & n24 ;
  assign n26 = ~n22 & ~n25 ;
  assign n27 = ~x14 & ~x15 ;
  assign n28 = ~x2 & ~x3 ;
  assign n29 = x0 & x1 ;
  assign n30 = n28 & n29 ;
  assign n31 = x2 & x3 ;
  assign n32 = ~x0 & ~x1 ;
  assign n33 = n31 & n32 ;
  assign n34 = ~n30 & ~n33 ;
  assign n35 = ~n27 & ~n34 ;
  assign n36 = x14 & x15 ;
  assign n37 = n28 & n36 ;
  assign n38 = x1 ^ x0 ;
  assign n39 = n37 & n38 ;
  assign n40 = ~n35 & ~n39 ;
  assign n41 = ~n28 & ~n31 ;
  assign n42 = x15 ^ x14 ;
  assign n43 = n32 ^ x15 ;
  assign n44 = n42 & n43 ;
  assign n45 = n44 ^ x14 ;
  assign n46 = ~n29 & n45 ;
  assign n47 = n41 & n46 ;
  assign n48 = n40 & ~n47 ;
  assign n49 = x4 & x5 ;
  assign n50 = ~x6 & ~x7 ;
  assign n51 = n49 & n50 ;
  assign n52 = ~x4 & ~x5 ;
  assign n53 = x6 & x7 ;
  assign n54 = n52 & n53 ;
  assign n55 = ~n51 & ~n54 ;
  assign n56 = ~n48 & ~n55 ;
  assign n57 = n36 & n50 ;
  assign n58 = n31 & n38 ;
  assign n59 = n29 & n41 ;
  assign n60 = ~n58 & ~n59 ;
  assign n61 = n57 & ~n60 ;
  assign n62 = n52 & n61 ;
  assign n63 = n31 & n50 ;
  assign n64 = n29 & n52 ;
  assign n65 = n63 & n64 ;
  assign n66 = n32 & n53 ;
  assign n67 = n28 & n49 ;
  assign n68 = n66 & n67 ;
  assign n69 = ~n65 & ~n68 ;
  assign n70 = ~n27 & ~n69 ;
  assign n71 = ~n62 & ~n70 ;
  assign n72 = ~n56 & n71 ;
  assign n73 = ~n26 & ~n72 ;
  assign n74 = ~n21 & ~n23 ;
  assign n75 = ~n20 & ~n24 ;
  assign n76 = ~n50 & ~n53 ;
  assign n77 = n32 & n49 ;
  assign n78 = ~n64 & ~n77 ;
  assign n79 = ~n27 & ~n78 ;
  assign n80 = n36 & n52 ;
  assign n81 = n38 & n80 ;
  assign n82 = ~n79 & ~n81 ;
  assign n83 = n41 & ~n82 ;
  assign n84 = n31 & n52 ;
  assign n85 = ~n67 & ~n84 ;
  assign n86 = n46 & ~n85 ;
  assign n87 = n37 & n64 ;
  assign n88 = ~n86 & ~n87 ;
  assign n89 = ~n83 & n88 ;
  assign n90 = ~n49 & ~n52 ;
  assign n91 = ~n48 & n90 ;
  assign n92 = n89 & ~n91 ;
  assign n93 = n76 & ~n92 ;
  assign n94 = n29 & n50 ;
  assign n95 = ~n66 & ~n94 ;
  assign n96 = ~n27 & ~n95 ;
  assign n97 = n38 & n57 ;
  assign n98 = ~n96 & ~n97 ;
  assign n99 = n41 & ~n98 ;
  assign n100 = n30 & n57 ;
  assign n101 = n28 & n53 ;
  assign n102 = ~n63 & ~n101 ;
  assign n103 = n46 & ~n102 ;
  assign n104 = ~n100 & ~n103 ;
  assign n105 = ~n99 & n104 ;
  assign n106 = n90 & ~n105 ;
  assign n107 = n72 & ~n106 ;
  assign n108 = ~n93 & n107 ;
  assign n109 = n75 & ~n108 ;
  assign n110 = n24 & n50 ;
  assign n111 = n20 & n53 ;
  assign n112 = ~n110 & ~n111 ;
  assign n113 = ~n89 & ~n112 ;
  assign n114 = n24 & n52 ;
  assign n115 = n46 & n114 ;
  assign n116 = n101 & n115 ;
  assign n117 = ~n113 & ~n116 ;
  assign n118 = n20 & n49 ;
  assign n119 = n94 & n118 ;
  assign n120 = n24 & n66 ;
  assign n121 = n52 & n120 ;
  assign n122 = ~n119 & ~n121 ;
  assign n123 = ~n27 & ~n122 ;
  assign n124 = n20 & n36 ;
  assign n125 = n38 & n124 ;
  assign n126 = n51 & n125 ;
  assign n127 = ~n123 & ~n126 ;
  assign n128 = n41 & ~n127 ;
  assign n129 = n20 & n50 ;
  assign n130 = n31 & n49 ;
  assign n131 = n46 & n130 ;
  assign n132 = n131 ^ n50 ;
  assign n133 = n29 & ~n85 ;
  assign n134 = n36 & n133 ;
  assign n135 = n134 ^ n129 ;
  assign n136 = ~n132 & n135 ;
  assign n137 = n136 ^ n134 ;
  assign n138 = n129 & n137 ;
  assign n139 = ~n128 & ~n138 ;
  assign n140 = n117 & n139 ;
  assign n141 = n20 & n31 ;
  assign n142 = n64 & n141 ;
  assign n143 = ~n27 & n142 ;
  assign n144 = ~n114 & ~n118 ;
  assign n145 = ~n48 & ~n144 ;
  assign n146 = ~n60 & n124 ;
  assign n147 = n52 & n146 ;
  assign n148 = n24 & n32 ;
  assign n149 = ~n27 & n148 ;
  assign n150 = n67 & n149 ;
  assign n151 = ~n147 & ~n150 ;
  assign n152 = ~n145 & n151 ;
  assign n153 = ~n143 & n152 ;
  assign n154 = n41 & n90 ;
  assign n155 = n20 & n29 ;
  assign n156 = ~n27 & n155 ;
  assign n157 = ~n149 & ~n156 ;
  assign n158 = ~n125 & n157 ;
  assign n159 = n154 & ~n158 ;
  assign n160 = n153 & ~n159 ;
  assign n161 = n76 & ~n160 ;
  assign n162 = n140 & ~n161 ;
  assign n163 = ~n109 & n162 ;
  assign n164 = n74 & ~n163 ;
  assign n165 = n23 & n36 ;
  assign n166 = n38 & n165 ;
  assign n167 = ~n27 & n29 ;
  assign n168 = n23 & n167 ;
  assign n169 = ~n166 & ~n168 ;
  assign n170 = n21 & n32 ;
  assign n171 = ~n27 & n170 ;
  assign n172 = n169 & ~n171 ;
  assign n173 = n154 & ~n172 ;
  assign n174 = n67 & n170 ;
  assign n175 = ~n27 & n174 ;
  assign n176 = n84 & n168 ;
  assign n177 = ~n175 & ~n176 ;
  assign n178 = ~n60 & n165 ;
  assign n179 = n52 & n178 ;
  assign n180 = n177 & ~n179 ;
  assign n181 = n21 & n52 ;
  assign n182 = n23 & n49 ;
  assign n183 = ~n181 & ~n182 ;
  assign n184 = ~n48 & ~n183 ;
  assign n185 = n30 & n165 ;
  assign n186 = n21 & n28 ;
  assign n187 = n23 & n31 ;
  assign n188 = ~n186 & ~n187 ;
  assign n189 = n46 & ~n188 ;
  assign n190 = ~n185 & ~n189 ;
  assign n191 = n90 & ~n190 ;
  assign n192 = ~n184 & ~n191 ;
  assign n193 = n180 & n192 ;
  assign n194 = ~n173 & n193 ;
  assign n195 = n75 & ~n194 ;
  assign n196 = ~n26 & ~n89 ;
  assign n197 = n155 & n182 ;
  assign n198 = n148 & n181 ;
  assign n199 = ~n197 & ~n198 ;
  assign n200 = ~n27 & ~n199 ;
  assign n201 = n118 & n166 ;
  assign n202 = ~n200 & ~n201 ;
  assign n203 = n41 & ~n202 ;
  assign n204 = ~n85 & n165 ;
  assign n205 = n155 & n204 ;
  assign n206 = ~n203 & ~n205 ;
  assign n207 = n114 & n186 ;
  assign n208 = n118 & n187 ;
  assign n209 = ~n207 & ~n208 ;
  assign n210 = n46 & ~n209 ;
  assign n211 = n206 & ~n210 ;
  assign n212 = ~n196 & n211 ;
  assign n213 = ~n195 & n212 ;
  assign n214 = n76 & ~n213 ;
  assign n215 = n21 & n50 ;
  assign n216 = n23 & n53 ;
  assign n217 = ~n215 & ~n216 ;
  assign n218 = ~n92 & ~n217 ;
  assign n219 = n54 & n186 ;
  assign n220 = n51 & n187 ;
  assign n221 = ~n219 & ~n220 ;
  assign n222 = n46 & ~n221 ;
  assign n223 = n94 & n187 ;
  assign n224 = n66 & n186 ;
  assign n225 = ~n223 & ~n224 ;
  assign n226 = ~n27 & ~n225 ;
  assign n227 = n50 & n178 ;
  assign n228 = ~n226 & ~n227 ;
  assign n229 = n90 & ~n228 ;
  assign n230 = ~n222 & ~n229 ;
  assign n231 = n51 & ~n169 ;
  assign n232 = n54 & n171 ;
  assign n233 = ~n231 & ~n232 ;
  assign n234 = n41 & ~n233 ;
  assign n235 = n94 & n204 ;
  assign n236 = ~n234 & ~n235 ;
  assign n237 = n230 & n236 ;
  assign n238 = ~n218 & n237 ;
  assign n239 = n75 & ~n238 ;
  assign n240 = n110 & n181 ;
  assign n241 = n118 & n216 ;
  assign n242 = ~n240 & ~n241 ;
  assign n243 = ~n48 & ~n242 ;
  assign n244 = n155 & n187 ;
  assign n245 = n148 & n186 ;
  assign n246 = ~n244 & ~n245 ;
  assign n247 = ~n27 & ~n246 ;
  assign n248 = n23 & n146 ;
  assign n249 = ~n247 & ~n248 ;
  assign n250 = ~n55 & ~n249 ;
  assign n251 = ~n243 & ~n250 ;
  assign n252 = ~n239 & n251 ;
  assign n253 = ~n214 & n252 ;
  assign n254 = ~n164 & n253 ;
  assign n255 = ~n73 & n254 ;
  assign n256 = n19 & ~n255 ;
  assign n257 = n18 & n36 ;
  assign n258 = ~n17 & ~n257 ;
  assign n259 = n23 & ~n258 ;
  assign n260 = ~n21 & ~n259 ;
  assign n261 = n38 & ~n260 ;
  assign n262 = n17 & n50 ;
  assign n263 = n21 & n262 ;
  assign n264 = ~n53 & ~n263 ;
  assign n265 = n261 & ~n264 ;
  assign n266 = n171 & n262 ;
  assign n267 = ~n18 & n29 ;
  assign n268 = ~n217 & n267 ;
  assign n269 = ~n18 & n53 ;
  assign n270 = n170 & n269 ;
  assign n271 = ~n23 & n29 ;
  assign n272 = n53 & n271 ;
  assign n273 = ~n270 & ~n272 ;
  assign n274 = ~n268 & n273 ;
  assign n275 = n23 & n29 ;
  assign n276 = n18 & n53 ;
  assign n277 = n275 & n276 ;
  assign n278 = ~n27 & n277 ;
  assign n279 = n274 & ~n278 ;
  assign n280 = ~n266 & n279 ;
  assign n281 = ~n265 & n280 ;
  assign n282 = n90 & ~n281 ;
  assign n283 = n17 & n52 ;
  assign n284 = n21 & n283 ;
  assign n285 = n29 & n284 ;
  assign n286 = n50 & n285 ;
  assign n287 = n182 & n276 ;
  assign n288 = n52 & n263 ;
  assign n289 = ~n287 & ~n288 ;
  assign n290 = n46 & ~n289 ;
  assign n291 = n18 & n23 ;
  assign n292 = n38 & ~n291 ;
  assign n293 = n17 & n23 ;
  assign n294 = ~n21 & ~n293 ;
  assign n295 = n32 & ~n294 ;
  assign n296 = ~n292 & ~n295 ;
  assign n297 = n49 & n53 ;
  assign n298 = ~n296 & n297 ;
  assign n299 = ~n290 & ~n298 ;
  assign n300 = ~n286 & n299 ;
  assign n301 = ~n282 & n300 ;
  assign n302 = n41 & ~n301 ;
  assign n303 = ~n18 & n21 ;
  assign n304 = ~n29 & ~n303 ;
  assign n305 = ~n17 & n32 ;
  assign n306 = ~n260 & ~n305 ;
  assign n307 = ~n304 & n306 ;
  assign n308 = n41 & n307 ;
  assign n309 = ~n188 & n267 ;
  assign n310 = ~n308 & ~n309 ;
  assign n311 = n38 & ~n258 ;
  assign n312 = n18 & n167 ;
  assign n313 = ~n311 & ~n312 ;
  assign n314 = n187 & ~n313 ;
  assign n315 = ~x0 & n17 ;
  assign n316 = ~x1 & n315 ;
  assign n317 = ~n27 & n316 ;
  assign n318 = n186 & n317 ;
  assign n319 = n17 & n28 ;
  assign n320 = ~n31 & ~n319 ;
  assign n321 = n21 & ~n320 ;
  assign n322 = n38 & n321 ;
  assign n323 = ~n318 & ~n322 ;
  assign n324 = n318 ^ n31 ;
  assign n325 = ~n18 & n32 ;
  assign n326 = n21 & n325 ;
  assign n327 = ~n271 & ~n326 ;
  assign n328 = n327 ^ n323 ;
  assign n329 = ~n324 & n328 ;
  assign n330 = n329 ^ n327 ;
  assign n331 = n323 & n330 ;
  assign n332 = ~n314 & n331 ;
  assign n333 = n310 & n332 ;
  assign n334 = n76 & n90 ;
  assign n335 = n55 & ~n334 ;
  assign n336 = ~n333 & ~n335 ;
  assign n337 = n17 & n38 ;
  assign n338 = n84 & n215 ;
  assign n339 = n337 & n338 ;
  assign n340 = n67 & n216 ;
  assign n341 = ~n338 & ~n340 ;
  assign n342 = n267 & ~n341 ;
  assign n343 = ~n34 & n297 ;
  assign n344 = ~n23 & n343 ;
  assign n345 = ~n342 & ~n344 ;
  assign n346 = n297 & n325 ;
  assign n347 = ~n188 & n346 ;
  assign n348 = ~n40 & ~n289 ;
  assign n349 = ~n347 & ~n348 ;
  assign n350 = n53 & ~n294 ;
  assign n351 = n67 & n350 ;
  assign n352 = n38 & n351 ;
  assign n353 = n349 & ~n352 ;
  assign n354 = n345 & n353 ;
  assign n355 = ~n339 & n354 ;
  assign n356 = ~n336 & n355 ;
  assign n357 = n72 & ~n93 ;
  assign n358 = n18 & n21 ;
  assign n359 = ~n293 & ~n358 ;
  assign n360 = ~n357 & ~n359 ;
  assign n361 = n131 & n291 ;
  assign n362 = ~n85 & n307 ;
  assign n363 = ~n29 & ~n45 ;
  assign n364 = n28 & n284 ;
  assign n365 = ~n363 & n364 ;
  assign n366 = n130 & ~n296 ;
  assign n367 = ~n365 & ~n366 ;
  assign n368 = ~n362 & n367 ;
  assign n369 = ~n361 & n368 ;
  assign n370 = n181 & n317 ;
  assign n371 = ~n183 & n267 ;
  assign n372 = n18 & n49 ;
  assign n373 = n168 & n372 ;
  assign n374 = ~n371 & ~n373 ;
  assign n375 = ~n370 & n374 ;
  assign n376 = n261 ^ n49 ;
  assign n377 = n376 ^ n375 ;
  assign n378 = n327 ^ n284 ;
  assign n379 = ~n261 & n378 ;
  assign n380 = n379 ^ n284 ;
  assign n381 = n377 & ~n380 ;
  assign n382 = n381 ^ n379 ;
  assign n383 = n382 ^ n284 ;
  assign n384 = n383 ^ n261 ;
  assign n385 = n375 & n384 ;
  assign n386 = n41 & ~n385 ;
  assign n387 = n369 & ~n386 ;
  assign n388 = n76 & ~n387 ;
  assign n389 = ~n360 & ~n388 ;
  assign n390 = n356 & n389 ;
  assign n391 = ~n302 & n390 ;
  assign n392 = n75 & ~n391 ;
  assign n393 = n24 & n28 ;
  assign n394 = n53 & n393 ;
  assign n395 = n64 & ~n294 ;
  assign n396 = ~n18 & n38 ;
  assign n397 = ~n316 & ~n396 ;
  assign n398 = ~n183 & ~n397 ;
  assign n399 = ~x1 & n23 ;
  assign n400 = x0 & n49 ;
  assign n401 = ~n399 & n400 ;
  assign n402 = ~n398 & ~n401 ;
  assign n403 = ~n395 & n402 ;
  assign n404 = n394 & ~n403 ;
  assign n405 = ~n140 & ~n359 ;
  assign n406 = n17 & n20 ;
  assign n407 = n21 & n406 ;
  assign n408 = n94 & n407 ;
  assign n409 = n24 & n53 ;
  assign n410 = x11 ^ x10 ;
  assign n411 = x10 ^ x1 ;
  assign n412 = n410 & n411 ;
  assign n413 = n412 ^ x10 ;
  assign n414 = n409 & n413 ;
  assign n415 = ~n408 & ~n414 ;
  assign n416 = n67 & ~n415 ;
  assign n417 = ~n405 & ~n416 ;
  assign n418 = ~n404 & n417 ;
  assign n419 = n417 ^ n112 ;
  assign n420 = n418 ^ n387 ;
  assign n421 = ~n419 & n420 ;
  assign n422 = n421 ^ n387 ;
  assign n423 = n418 & n422 ;
  assign n424 = ~n392 & n423 ;
  assign n425 = ~n256 & n424 ;
  assign n426 = ~n262 & ~n276 ;
  assign n427 = ~n92 & ~n426 ;
  assign n428 = n18 & n31 ;
  assign n429 = ~n319 & ~n428 ;
  assign n430 = n46 & ~n429 ;
  assign n431 = ~n315 & ~n396 ;
  assign n432 = n31 & ~n431 ;
  assign n433 = n30 & ~n258 ;
  assign n434 = ~n432 & ~n433 ;
  assign n435 = ~n430 & n434 ;
  assign n436 = n90 & ~n435 ;
  assign n437 = n33 & n49 ;
  assign n438 = ~n133 & ~n437 ;
  assign n439 = ~n18 & ~n438 ;
  assign n440 = n84 & n311 ;
  assign n441 = n67 & n337 ;
  assign n442 = ~n440 & ~n441 ;
  assign n443 = n67 & n316 ;
  assign n444 = n64 & n428 ;
  assign n445 = ~n443 & ~n444 ;
  assign n446 = ~n27 & ~n445 ;
  assign n447 = n442 & ~n446 ;
  assign n448 = ~n439 & n447 ;
  assign n449 = ~n283 & ~n372 ;
  assign n450 = ~n48 & ~n449 ;
  assign n451 = n448 & ~n450 ;
  assign n452 = ~n436 & n451 ;
  assign n453 = n76 & ~n452 ;
  assign n454 = ~n267 & ~n311 ;
  assign n455 = n63 & ~n454 ;
  assign n456 = n66 & n319 ;
  assign n457 = n94 & n428 ;
  assign n458 = ~n456 & ~n457 ;
  assign n459 = ~n27 & ~n458 ;
  assign n460 = ~n34 & n269 ;
  assign n461 = n101 & n337 ;
  assign n462 = ~n460 & ~n461 ;
  assign n463 = ~n459 & n462 ;
  assign n464 = ~n455 & n463 ;
  assign n465 = n90 & ~n464 ;
  assign n466 = n130 & ~n397 ;
  assign n467 = n50 & n466 ;
  assign n468 = n85 & ~n154 ;
  assign n469 = n94 & ~n258 ;
  assign n470 = n53 & ~n431 ;
  assign n471 = ~n469 & ~n470 ;
  assign n472 = ~n468 & ~n471 ;
  assign n473 = n54 & n319 ;
  assign n474 = ~n29 & n428 ;
  assign n475 = n45 & n474 ;
  assign n476 = n51 & n475 ;
  assign n477 = ~n473 & ~n476 ;
  assign n478 = ~n363 & ~n477 ;
  assign n479 = ~n472 & ~n478 ;
  assign n480 = ~n467 & n479 ;
  assign n481 = ~n465 & n480 ;
  assign n482 = ~n453 & n481 ;
  assign n483 = ~n427 & n482 ;
  assign n484 = n75 & ~n483 ;
  assign n485 = n24 & n49 ;
  assign n486 = n325 & n485 ;
  assign n487 = n118 & ~n313 ;
  assign n488 = n267 ^ n114 ;
  assign n489 = n267 ^ n118 ;
  assign n490 = n489 ^ n118 ;
  assign n491 = ~n317 & ~n337 ;
  assign n492 = n491 ^ n118 ;
  assign n493 = ~n490 & n492 ;
  assign n494 = n493 ^ n118 ;
  assign n495 = n488 & n494 ;
  assign n496 = n495 ^ n114 ;
  assign n497 = ~n487 & ~n496 ;
  assign n498 = ~n486 & n497 ;
  assign n499 = n41 & ~n498 ;
  assign n500 = n18 & n24 ;
  assign n501 = ~n406 & ~n500 ;
  assign n502 = ~n92 & ~n501 ;
  assign n503 = n20 & n466 ;
  assign n504 = n155 & ~n258 ;
  assign n505 = n24 & ~n431 ;
  assign n506 = ~n504 & ~n505 ;
  assign n507 = ~n468 & ~n506 ;
  assign n508 = n114 & n319 ;
  assign n509 = n118 & n474 ;
  assign n510 = ~n508 & ~n509 ;
  assign n511 = ~n363 & ~n510 ;
  assign n512 = ~n507 & ~n511 ;
  assign n513 = ~n503 & n512 ;
  assign n514 = ~n502 & n513 ;
  assign n515 = ~n499 & n514 ;
  assign n516 = n76 & ~n515 ;
  assign n517 = ~n107 & ~n501 ;
  assign n518 = ~n141 & ~n393 ;
  assign n519 = n346 & ~n518 ;
  assign n520 = ~n517 & ~n519 ;
  assign n521 = ~n516 & n520 ;
  assign n522 = ~n167 & ~n317 ;
  assign n523 = n454 & n522 ;
  assign n524 = n90 & ~n523 ;
  assign n525 = n64 & ~n258 ;
  assign n526 = ~n29 & n49 ;
  assign n527 = ~n305 & n526 ;
  assign n528 = ~n18 & n527 ;
  assign n529 = ~n525 & ~n528 ;
  assign n530 = ~n524 & n529 ;
  assign n531 = n76 & ~n530 ;
  assign n532 = n94 & n372 ;
  assign n533 = n66 & n283 ;
  assign n534 = ~n532 & ~n533 ;
  assign n535 = ~n27 & ~n534 ;
  assign n536 = n54 & n337 ;
  assign n537 = ~n346 & ~n536 ;
  assign n538 = ~n535 & n537 ;
  assign n539 = n267 ^ n51 ;
  assign n540 = n267 ^ n54 ;
  assign n541 = n540 ^ n54 ;
  assign n542 = n311 ^ n54 ;
  assign n543 = ~n541 & ~n542 ;
  assign n544 = n543 ^ n54 ;
  assign n545 = n539 & n544 ;
  assign n546 = n545 ^ n51 ;
  assign n547 = n538 & ~n546 ;
  assign n548 = ~n531 & n547 ;
  assign n549 = n75 & ~n548 ;
  assign n550 = ~n55 & ~n506 ;
  assign n551 = n111 & ~n397 ;
  assign n552 = n49 & n551 ;
  assign n553 = n110 & n283 ;
  assign n554 = n111 & n372 ;
  assign n555 = ~n553 & ~n554 ;
  assign n556 = n45 ^ n29 ;
  assign n557 = n556 ^ n45 ;
  assign n558 = n553 ^ n45 ;
  assign n559 = n557 & n558 ;
  assign n560 = n559 ^ n45 ;
  assign n561 = ~n555 & n560 ;
  assign n562 = ~n552 & ~n561 ;
  assign n563 = ~n550 & n562 ;
  assign n564 = ~n549 & n563 ;
  assign n565 = n41 & ~n564 ;
  assign n566 = ~n18 & n120 ;
  assign n567 = n110 & ~n491 ;
  assign n568 = ~n566 & ~n567 ;
  assign n569 = n267 ^ n111 ;
  assign n570 = n267 ^ n110 ;
  assign n571 = n570 ^ n110 ;
  assign n572 = n313 ^ n110 ;
  assign n573 = ~n571 & n572 ;
  assign n574 = n573 ^ n110 ;
  assign n575 = n569 & n574 ;
  assign n576 = n575 ^ n111 ;
  assign n577 = n568 & ~n576 ;
  assign n578 = n41 & ~n577 ;
  assign n579 = ~n102 & ~n506 ;
  assign n580 = n31 & n551 ;
  assign n581 = n262 & n393 ;
  assign n582 = n581 ^ n29 ;
  assign n583 = n582 ^ n581 ;
  assign n584 = n581 ^ n45 ;
  assign n585 = ~n583 & n584 ;
  assign n586 = n585 ^ n581 ;
  assign n587 = n141 & n276 ;
  assign n588 = ~n581 & ~n587 ;
  assign n589 = n588 ^ n580 ;
  assign n590 = ~n586 & ~n589 ;
  assign n591 = n590 ^ n588 ;
  assign n592 = ~n580 & n591 ;
  assign n593 = n592 ^ n580 ;
  assign n594 = n593 ^ n580 ;
  assign n595 = ~n579 & n594 ;
  assign n596 = ~n578 & n595 ;
  assign n597 = n90 & ~n596 ;
  assign n598 = ~n267 & ~n337 ;
  assign n599 = n84 & n110 ;
  assign n600 = n67 & n111 ;
  assign n601 = ~n599 & ~n600 ;
  assign n602 = ~n598 & ~n601 ;
  assign n603 = ~n597 & ~n602 ;
  assign n604 = n393 & ~n598 ;
  assign n605 = n141 & ~n454 ;
  assign n606 = n24 & n31 ;
  assign n607 = n325 & n606 ;
  assign n608 = n148 & n319 ;
  assign n609 = n155 & n428 ;
  assign n610 = ~n608 & ~n609 ;
  assign n611 = ~n27 & ~n610 ;
  assign n612 = ~n607 & ~n611 ;
  assign n613 = ~n605 & n612 ;
  assign n614 = ~n604 & n613 ;
  assign n615 = ~n335 & ~n614 ;
  assign n616 = ~n40 & ~n555 ;
  assign n617 = ~n615 & ~n616 ;
  assign n618 = n603 & n617 ;
  assign n619 = ~n565 & n618 ;
  assign n620 = n521 & n619 ;
  assign n621 = ~n484 & n620 ;
  assign n622 = n74 & ~n621 ;
  assign n623 = n20 & n61 ;
  assign n624 = ~n48 & ~n112 ;
  assign n625 = n63 & n155 ;
  assign n626 = n28 & n120 ;
  assign n627 = ~n625 & ~n626 ;
  assign n628 = ~n27 & ~n627 ;
  assign n629 = ~n624 & ~n628 ;
  assign n630 = ~n623 & n629 ;
  assign n631 = n46 & ~n518 ;
  assign n632 = n30 & n124 ;
  assign n633 = ~n631 & ~n632 ;
  assign n634 = n76 & ~n633 ;
  assign n635 = n630 & ~n634 ;
  assign n636 = n74 & ~n635 ;
  assign n637 = n155 & n216 ;
  assign n638 = n110 & n170 ;
  assign n639 = ~n637 & ~n638 ;
  assign n640 = ~n27 & ~n639 ;
  assign n641 = n111 & n166 ;
  assign n642 = ~n640 & ~n641 ;
  assign n643 = n41 & ~n642 ;
  assign n644 = n124 & n275 ;
  assign n645 = ~n102 & n644 ;
  assign n646 = ~n643 & ~n645 ;
  assign n647 = ~n26 & ~n48 ;
  assign n648 = n249 & ~n647 ;
  assign n649 = n76 & ~n648 ;
  assign n650 = n215 & n393 ;
  assign n651 = n111 & n187 ;
  assign n652 = ~n650 & ~n651 ;
  assign n653 = n46 & ~n652 ;
  assign n654 = ~n26 & ~n105 ;
  assign n655 = ~n653 & ~n654 ;
  assign n656 = ~n649 & n655 ;
  assign n657 = n646 & n656 ;
  assign n658 = ~n636 & n657 ;
  assign n659 = n19 & ~n658 ;
  assign n660 = n22 & n262 ;
  assign n661 = n216 & n500 ;
  assign n662 = ~n660 & ~n661 ;
  assign n663 = n46 & ~n662 ;
  assign n664 = ~n29 & n296 ;
  assign n665 = n409 & ~n664 ;
  assign n666 = ~n663 & ~n665 ;
  assign n667 = ~n408 & n666 ;
  assign n668 = n41 & ~n667 ;
  assign n669 = ~n112 & ~n333 ;
  assign n670 = ~n668 & ~n669 ;
  assign n671 = n31 & n53 ;
  assign n672 = ~n296 & n671 ;
  assign n673 = ~n105 & ~n359 ;
  assign n674 = ~n102 & n307 ;
  assign n675 = n17 & n94 ;
  assign n676 = n186 & n675 ;
  assign n677 = n215 & n319 ;
  assign n678 = n187 & n276 ;
  assign n679 = ~n677 & ~n678 ;
  assign n680 = n46 & ~n679 ;
  assign n681 = ~n676 & ~n680 ;
  assign n682 = ~n674 & n681 ;
  assign n683 = ~n673 & n682 ;
  assign n684 = ~n672 & n683 ;
  assign n685 = n75 & ~n684 ;
  assign n686 = ~n359 & ~n630 ;
  assign n687 = ~n188 & n566 ;
  assign n688 = n22 & n63 ;
  assign n689 = n23 & n394 ;
  assign n690 = ~n688 & ~n689 ;
  assign n691 = n267 & ~n690 ;
  assign n692 = ~n409 & ~n660 ;
  assign n693 = n58 & ~n692 ;
  assign n694 = ~n691 & ~n693 ;
  assign n695 = ~n20 & n31 ;
  assign n696 = n29 & n695 ;
  assign n697 = ~n23 & n24 ;
  assign n698 = ~n34 & n697 ;
  assign n699 = ~n696 & ~n698 ;
  assign n700 = n38 & n393 ;
  assign n701 = ~n294 & n700 ;
  assign n702 = n699 & ~n701 ;
  assign n703 = n53 & ~n702 ;
  assign n704 = n694 & ~n703 ;
  assign n705 = ~n687 & n704 ;
  assign n706 = ~n40 & ~n662 ;
  assign n707 = n705 & ~n706 ;
  assign n708 = ~n686 & n707 ;
  assign n709 = ~n685 & n708 ;
  assign n710 = n670 & n709 ;
  assign n711 = ~n659 & n710 ;
  assign n712 = n90 & ~n711 ;
  assign n713 = ~n144 & ~n333 ;
  assign n714 = n41 & ~n158 ;
  assign n715 = n633 & ~n714 ;
  assign n716 = ~n359 & ~n715 ;
  assign n717 = n307 & ~n518 ;
  assign n718 = n606 & ~n664 ;
  assign n719 = n186 & n406 ;
  assign n720 = n187 & n500 ;
  assign n721 = ~n29 & n720 ;
  assign n722 = ~n719 & ~n721 ;
  assign n723 = ~n363 & ~n722 ;
  assign n724 = ~n718 & ~n723 ;
  assign n725 = ~n717 & n724 ;
  assign n726 = ~n716 & n725 ;
  assign n727 = n90 & ~n726 ;
  assign n728 = n22 & n283 ;
  assign n729 = n182 & n500 ;
  assign n730 = ~n728 & ~n729 ;
  assign n731 = ~n40 & ~n730 ;
  assign n732 = ~n188 & n486 ;
  assign n733 = n22 & n84 ;
  assign n734 = n25 & n67 ;
  assign n735 = ~n733 & ~n734 ;
  assign n736 = n267 & ~n735 ;
  assign n737 = ~n732 & ~n736 ;
  assign n738 = ~n485 & ~n728 ;
  assign n739 = n58 & ~n738 ;
  assign n740 = n737 & ~n739 ;
  assign n741 = ~n731 & n740 ;
  assign n742 = n740 ^ n49 ;
  assign n743 = n741 ^ n702 ;
  assign n744 = n742 & n743 ;
  assign n745 = n744 ^ n702 ;
  assign n746 = n741 & n745 ;
  assign n747 = ~n727 & n746 ;
  assign n748 = ~n24 & ~n407 ;
  assign n749 = n261 & ~n748 ;
  assign n750 = n275 & n500 ;
  assign n751 = n32 & n407 ;
  assign n752 = ~n750 & ~n751 ;
  assign n753 = ~n27 & ~n752 ;
  assign n754 = ~n26 & n267 ;
  assign n755 = n24 & ~n327 ;
  assign n756 = ~n754 & ~n755 ;
  assign n757 = ~n753 & n756 ;
  assign n758 = ~n749 & n757 ;
  assign n759 = n90 & ~n758 ;
  assign n760 = n46 & ~n730 ;
  assign n761 = n485 & ~n664 ;
  assign n762 = n20 & n285 ;
  assign n763 = ~n761 & ~n762 ;
  assign n764 = ~n760 & n763 ;
  assign n765 = ~n759 & n764 ;
  assign n766 = n41 & ~n765 ;
  assign n767 = ~n153 & ~n359 ;
  assign n768 = ~n766 & ~n767 ;
  assign n769 = n747 & n768 ;
  assign n770 = ~n713 & n769 ;
  assign n771 = n76 & ~n770 ;
  assign n772 = ~n88 & ~n662 ;
  assign n773 = ~n82 & ~n662 ;
  assign n774 = ~n183 & n566 ;
  assign n775 = n118 & n215 ;
  assign n776 = n25 & n54 ;
  assign n777 = ~n775 & ~n776 ;
  assign n778 = n267 & ~n777 ;
  assign n779 = ~n78 & n697 ;
  assign n780 = n53 & n779 ;
  assign n781 = ~n778 & ~n780 ;
  assign n782 = n29 & n297 ;
  assign n783 = ~n20 & n782 ;
  assign n784 = n781 & ~n783 ;
  assign n785 = n49 & ~n692 ;
  assign n786 = n114 & n350 ;
  assign n787 = ~n785 & ~n786 ;
  assign n788 = n38 & ~n787 ;
  assign n789 = n784 & ~n788 ;
  assign n790 = ~n774 & n789 ;
  assign n791 = ~n773 & n790 ;
  assign n792 = n791 ^ x2 ;
  assign n793 = n792 ^ x3 ;
  assign n794 = n793 ^ n791 ;
  assign n795 = n794 ^ n772 ;
  assign n796 = ~n397 & ~n777 ;
  assign n814 = n52 & ~n692 ;
  assign n797 = ~n21 & n32 ;
  assign n798 = ~n23 & n52 ;
  assign n799 = ~n797 & n798 ;
  assign n800 = ~n49 & ~n799 ;
  assign n801 = n800 ^ n53 ;
  assign n802 = x9 ^ x8 ;
  assign n803 = x4 & ~n32 ;
  assign n804 = n803 ^ x8 ;
  assign n805 = n802 & n804 ;
  assign n806 = n805 ^ x8 ;
  assign n807 = n806 ^ n800 ;
  assign n808 = ~n801 & ~n807 ;
  assign n809 = n808 ^ n805 ;
  assign n810 = n809 ^ x8 ;
  assign n811 = n810 ^ n53 ;
  assign n812 = ~n800 & n811 ;
  assign n813 = n812 ^ n800 ;
  assign n815 = n814 ^ n813 ;
  assign n816 = n815 ^ n29 ;
  assign n826 = n816 ^ n815 ;
  assign n817 = n129 & ~n260 ;
  assign n818 = ~n110 & ~n817 ;
  assign n819 = ~n53 & n818 ;
  assign n820 = n819 ^ n816 ;
  assign n821 = n820 ^ n815 ;
  assign n822 = n816 ^ n813 ;
  assign n823 = n822 ^ n819 ;
  assign n824 = n823 ^ n821 ;
  assign n825 = n821 & n824 ;
  assign n827 = n826 ^ n825 ;
  assign n828 = n827 ^ n821 ;
  assign n829 = n815 ^ n49 ;
  assign n830 = n825 ^ n821 ;
  assign n831 = ~n829 & n830 ;
  assign n832 = n831 ^ n815 ;
  assign n833 = ~n828 & ~n832 ;
  assign n834 = n833 ^ n815 ;
  assign n835 = n834 ^ n814 ;
  assign n836 = n835 ^ n815 ;
  assign n837 = ~n796 & ~n836 ;
  assign n838 = n837 ^ x3 ;
  assign n839 = ~n837 & ~n838 ;
  assign n840 = n839 ^ n791 ;
  assign n841 = n840 ^ n837 ;
  assign n842 = n795 & n841 ;
  assign n843 = n842 ^ n839 ;
  assign n844 = n843 ^ n837 ;
  assign n845 = ~n772 & ~n844 ;
  assign n846 = n845 ^ n772 ;
  assign n847 = ~n771 & ~n846 ;
  assign n848 = ~n712 & n847 ;
  assign n849 = ~n622 & n848 ;
  assign n850 = n425 & n849 ;
  assign y0 = ~n850 ;
endmodule
