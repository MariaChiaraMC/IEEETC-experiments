module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 ;
  assign n11 = ~x0 & x4 ;
  assign n12 = ~x2 & x3 ;
  assign n13 = x5 & ~x6 ;
  assign n14 = x7 & x8 ;
  assign n15 = ~x9 & n14 ;
  assign n16 = n13 & n15 ;
  assign n17 = ~x5 & x6 ;
  assign n18 = ~x8 & x9 ;
  assign n19 = ~x7 & n18 ;
  assign n20 = n17 & n19 ;
  assign n21 = ~n16 & ~n20 ;
  assign n22 = n12 & ~n21 ;
  assign n23 = x2 & ~x9 ;
  assign n24 = ~x6 & x7 ;
  assign n25 = ~x3 & ~x5 ;
  assign n26 = n24 & n25 ;
  assign n27 = n23 & n26 ;
  assign n28 = ~x8 & n27 ;
  assign n29 = ~n22 & ~n28 ;
  assign n30 = n11 & ~n29 ;
  assign n31 = x4 ^ x1 ;
  assign n32 = x2 & ~x5 ;
  assign n33 = ~x7 & ~x8 ;
  assign n34 = x6 & n33 ;
  assign n35 = n34 ^ x1 ;
  assign n36 = ~x3 & ~x9 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = n37 ^ n24 ;
  assign n40 = ~n38 & n39 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = x8 & x9 ;
  assign n43 = x3 & n42 ;
  assign n44 = ~n37 & ~n43 ;
  assign n45 = n44 ^ n35 ;
  assign n46 = ~n41 & ~n45 ;
  assign n47 = n46 ^ n44 ;
  assign n48 = ~n35 & n47 ;
  assign n49 = n48 ^ n34 ;
  assign n50 = n49 ^ n35 ;
  assign n51 = n32 & ~n50 ;
  assign n52 = n51 ^ n31 ;
  assign n53 = n52 ^ x4 ;
  assign n54 = n53 ^ n52 ;
  assign n83 = x4 ^ x2 ;
  assign n95 = n83 ^ x2 ;
  assign n55 = x5 & x6 ;
  assign n56 = x8 & ~x9 ;
  assign n57 = n55 & n56 ;
  assign n58 = ~x7 & n57 ;
  assign n59 = ~x6 & ~x7 ;
  assign n60 = ~x5 & n59 ;
  assign n61 = x9 ^ x6 ;
  assign n62 = x7 & n61 ;
  assign n63 = ~n60 & ~n62 ;
  assign n64 = ~x5 & ~n56 ;
  assign n65 = ~n63 & ~n64 ;
  assign n66 = n65 ^ x3 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = x9 ^ x5 ;
  assign n69 = x9 ^ x7 ;
  assign n70 = n69 ^ x7 ;
  assign n71 = x6 & x7 ;
  assign n72 = n71 ^ x7 ;
  assign n73 = n70 & ~n72 ;
  assign n74 = n73 ^ x7 ;
  assign n75 = ~n68 & ~n74 ;
  assign n76 = ~x8 & n75 ;
  assign n77 = n76 ^ n65 ;
  assign n78 = ~n67 & n77 ;
  assign n79 = n78 ^ n65 ;
  assign n80 = ~n58 & ~n79 ;
  assign n81 = ~x4 & ~n80 ;
  assign n82 = n81 ^ x2 ;
  assign n84 = n83 ^ n82 ;
  assign n85 = n84 ^ n83 ;
  assign n86 = n85 ^ x2 ;
  assign n87 = x6 & ~x7 ;
  assign n88 = x3 & x5 ;
  assign n89 = n42 & n88 ;
  assign n90 = n87 & n89 ;
  assign n91 = n90 ^ n84 ;
  assign n92 = n91 ^ n84 ;
  assign n93 = n92 ^ n86 ;
  assign n94 = ~n86 & n93 ;
  assign n96 = n95 ^ n94 ;
  assign n97 = n96 ^ n86 ;
  assign n98 = ~x6 & ~x9 ;
  assign n99 = ~x2 & x5 ;
  assign n100 = n33 ^ n14 ;
  assign n101 = ~x3 & n100 ;
  assign n102 = n101 ^ n33 ;
  assign n103 = n99 & n102 ;
  assign n104 = n98 & n103 ;
  assign n105 = n18 & n71 ;
  assign n106 = ~x2 & n25 ;
  assign n107 = ~n88 & ~n106 ;
  assign n108 = n105 & ~n107 ;
  assign n109 = x5 & n71 ;
  assign n110 = ~n60 & ~n109 ;
  assign n111 = n18 & ~n25 ;
  assign n112 = n111 ^ x3 ;
  assign n113 = n112 ^ n111 ;
  assign n114 = n111 ^ n42 ;
  assign n115 = n114 ^ n111 ;
  assign n116 = ~n113 & n115 ;
  assign n117 = n116 ^ n111 ;
  assign n118 = ~x2 & n117 ;
  assign n119 = n118 ^ n111 ;
  assign n120 = ~n110 & n119 ;
  assign n121 = ~n108 & ~n120 ;
  assign n122 = ~n104 & n121 ;
  assign n123 = n122 ^ x2 ;
  assign n124 = n94 ^ n86 ;
  assign n125 = ~n123 & ~n124 ;
  assign n126 = n125 ^ x2 ;
  assign n127 = n97 & ~n126 ;
  assign n128 = n127 ^ x2 ;
  assign n129 = n128 ^ x4 ;
  assign n130 = n129 ^ x2 ;
  assign n131 = n130 ^ n52 ;
  assign n132 = n131 ^ n31 ;
  assign n133 = ~n54 & ~n132 ;
  assign n134 = n133 ^ n130 ;
  assign n135 = x2 & x3 ;
  assign n136 = ~n59 & ~n71 ;
  assign n137 = x5 & x8 ;
  assign n138 = ~n136 & n137 ;
  assign n139 = ~n34 & ~n138 ;
  assign n140 = x9 & ~n139 ;
  assign n141 = ~n16 & ~n140 ;
  assign n142 = n135 & ~n141 ;
  assign n143 = ~n130 & ~n142 ;
  assign n144 = n143 ^ n31 ;
  assign n145 = ~n134 & ~n144 ;
  assign n146 = n145 ^ n143 ;
  assign n147 = ~n31 & n146 ;
  assign n148 = n147 ^ n133 ;
  assign n149 = n148 ^ x1 ;
  assign n150 = n149 ^ n130 ;
  assign n151 = x0 & n150 ;
  assign n152 = n151 ^ n30 ;
  assign n156 = x3 & x4 ;
  assign n157 = ~x2 & n156 ;
  assign n158 = x6 & x9 ;
  assign n159 = ~x7 & n158 ;
  assign n160 = n157 & n159 ;
  assign n153 = ~x3 & ~x4 ;
  assign n161 = ~x4 & ~x7 ;
  assign n162 = ~x3 & n24 ;
  assign n163 = ~n161 & ~n162 ;
  assign n164 = n23 & ~n163 ;
  assign n165 = ~n153 & n164 ;
  assign n166 = ~n160 & ~n165 ;
  assign n154 = ~x2 & n24 ;
  assign n155 = n153 & n154 ;
  assign n167 = n166 ^ n155 ;
  assign n168 = n167 ^ n166 ;
  assign n169 = n166 ^ x9 ;
  assign n170 = n169 ^ n166 ;
  assign n171 = n168 & ~n170 ;
  assign n172 = n171 ^ n166 ;
  assign n173 = x8 & ~n172 ;
  assign n174 = n173 ^ n166 ;
  assign n175 = ~x5 & ~n174 ;
  assign n176 = ~x4 & ~x9 ;
  assign n177 = ~n137 & n176 ;
  assign n178 = x6 ^ x5 ;
  assign n179 = n177 & n178 ;
  assign n180 = n179 ^ x4 ;
  assign n181 = n180 ^ x7 ;
  assign n193 = n181 ^ n180 ;
  assign n182 = n136 ^ x6 ;
  assign n183 = n178 ^ x6 ;
  assign n184 = ~n182 & n183 ;
  assign n185 = n184 ^ x6 ;
  assign n186 = n18 & ~n185 ;
  assign n187 = n186 ^ n181 ;
  assign n188 = n187 ^ n180 ;
  assign n189 = n181 ^ n179 ;
  assign n190 = n189 ^ n186 ;
  assign n191 = n190 ^ n188 ;
  assign n192 = n188 & ~n191 ;
  assign n194 = n193 ^ n192 ;
  assign n195 = n194 ^ n188 ;
  assign n196 = n180 ^ n57 ;
  assign n197 = n192 ^ n188 ;
  assign n198 = ~n196 & n197 ;
  assign n199 = n198 ^ n180 ;
  assign n200 = ~n195 & n199 ;
  assign n201 = n200 ^ n180 ;
  assign n202 = n201 ^ x4 ;
  assign n203 = n202 ^ n180 ;
  assign n204 = ~x2 & n203 ;
  assign n205 = x7 & x9 ;
  assign n206 = x4 & n205 ;
  assign n207 = ~x5 & ~x6 ;
  assign n208 = n206 & n207 ;
  assign n209 = ~n204 & ~n208 ;
  assign n210 = x2 & x4 ;
  assign n211 = x7 & ~x9 ;
  assign n212 = n55 & n211 ;
  assign n213 = n212 ^ x5 ;
  assign n214 = n213 ^ n212 ;
  assign n215 = ~n59 & ~n205 ;
  assign n216 = n215 ^ n212 ;
  assign n217 = n216 ^ n212 ;
  assign n218 = ~n214 & n217 ;
  assign n219 = n218 ^ n212 ;
  assign n220 = x8 & n219 ;
  assign n221 = n220 ^ n212 ;
  assign n222 = n210 & n221 ;
  assign n223 = ~x3 & ~n222 ;
  assign n224 = n209 & n223 ;
  assign n225 = ~x2 & ~x6 ;
  assign n226 = x4 & ~x5 ;
  assign n227 = n226 ^ x8 ;
  assign n228 = n227 ^ x7 ;
  assign n233 = n228 ^ n226 ;
  assign n229 = n228 ^ x7 ;
  assign n230 = n229 ^ n226 ;
  assign n231 = n230 ^ n70 ;
  assign n232 = ~n230 & ~n231 ;
  assign n234 = n233 ^ n232 ;
  assign n235 = n234 ^ n230 ;
  assign n236 = ~x4 & x5 ;
  assign n237 = n236 ^ n226 ;
  assign n238 = n232 ^ n230 ;
  assign n239 = n237 & ~n238 ;
  assign n240 = n239 ^ n226 ;
  assign n241 = ~n235 & n240 ;
  assign n242 = n241 ^ n226 ;
  assign n243 = n242 ^ n226 ;
  assign n244 = n225 & n243 ;
  assign n261 = n13 & n206 ;
  assign n262 = ~x7 & ~x9 ;
  assign n263 = n207 & n262 ;
  assign n264 = ~n261 & ~n263 ;
  assign n245 = n71 & n226 ;
  assign n246 = x4 & x9 ;
  assign n247 = x5 & ~x7 ;
  assign n248 = n246 & n247 ;
  assign n249 = ~n245 & ~n248 ;
  assign n250 = ~x4 & x9 ;
  assign n251 = n59 & n250 ;
  assign n252 = n251 ^ n62 ;
  assign n253 = n252 ^ n251 ;
  assign n254 = n251 ^ x4 ;
  assign n255 = n254 ^ n251 ;
  assign n256 = n253 & ~n255 ;
  assign n257 = n256 ^ n251 ;
  assign n258 = x5 & n257 ;
  assign n259 = n258 ^ n251 ;
  assign n260 = n249 & ~n259 ;
  assign n265 = n264 ^ n260 ;
  assign n266 = n264 ^ x8 ;
  assign n267 = n266 ^ n264 ;
  assign n268 = n267 ^ n135 ;
  assign n269 = n268 ^ x3 ;
  assign n270 = n265 & n269 ;
  assign n271 = n270 ^ n264 ;
  assign n272 = n135 & n271 ;
  assign n273 = n272 ^ n135 ;
  assign n274 = n273 ^ x3 ;
  assign n275 = ~n244 & n274 ;
  assign n276 = ~n224 & ~n275 ;
  assign n277 = n109 & n210 ;
  assign n278 = n42 & n277 ;
  assign n279 = ~n276 & ~n278 ;
  assign n280 = ~x0 & ~n279 ;
  assign n281 = ~n175 & ~n280 ;
  assign n282 = n281 ^ x1 ;
  assign n283 = n282 ^ n281 ;
  assign n284 = ~x5 & x8 ;
  assign n285 = ~x2 & ~x3 ;
  assign n286 = ~x4 & x6 ;
  assign n287 = n285 & n286 ;
  assign n288 = x3 & ~x6 ;
  assign n289 = ~n98 & ~n286 ;
  assign n290 = x2 & ~n153 ;
  assign n291 = ~n289 & n290 ;
  assign n292 = n291 ^ n246 ;
  assign n293 = ~n288 & n292 ;
  assign n294 = n293 ^ n246 ;
  assign n295 = ~n287 & ~n294 ;
  assign n296 = ~x7 & ~n295 ;
  assign n297 = ~x2 & x9 ;
  assign n298 = n156 ^ n153 ;
  assign n299 = n298 ^ n297 ;
  assign n300 = n156 ^ x7 ;
  assign n301 = n156 ^ x6 ;
  assign n302 = n301 ^ n300 ;
  assign n303 = n300 & n302 ;
  assign n304 = n303 ^ n156 ;
  assign n305 = n304 ^ n300 ;
  assign n306 = n299 & n305 ;
  assign n307 = n306 ^ n303 ;
  assign n308 = n307 ^ n300 ;
  assign n309 = n297 & n308 ;
  assign n310 = ~n296 & ~n309 ;
  assign n311 = ~x9 & n71 ;
  assign n312 = ~x2 & n311 ;
  assign n313 = x4 ^ x3 ;
  assign n314 = n312 & n313 ;
  assign n315 = n310 & ~n314 ;
  assign n316 = ~x0 & ~n315 ;
  assign n317 = ~n136 & ~n225 ;
  assign n318 = n250 & n317 ;
  assign n319 = x4 & ~n98 ;
  assign n320 = ~n154 & ~n262 ;
  assign n321 = n319 & ~n320 ;
  assign n322 = x0 & n321 ;
  assign n323 = ~n318 & ~n322 ;
  assign n324 = ~x3 & ~n323 ;
  assign n325 = x0 & ~x2 ;
  assign n326 = n71 & n325 ;
  assign n327 = ~x3 & x4 ;
  assign n328 = ~n176 & ~n327 ;
  assign n329 = n326 & n328 ;
  assign n330 = ~n324 & ~n329 ;
  assign n331 = ~n316 & n330 ;
  assign n332 = n284 & ~n331 ;
  assign n333 = ~x0 & x7 ;
  assign n334 = n32 & n333 ;
  assign n335 = n158 & n334 ;
  assign n336 = x0 & n247 ;
  assign n337 = x3 & n336 ;
  assign n338 = n297 ^ n23 ;
  assign n339 = ~x6 & n338 ;
  assign n340 = n339 ^ n297 ;
  assign n341 = n337 & n340 ;
  assign n342 = ~n335 & ~n341 ;
  assign n343 = ~x4 & ~n342 ;
  assign n344 = x3 & n17 ;
  assign n345 = n325 & n344 ;
  assign n346 = n206 & n345 ;
  assign n347 = ~n343 & ~n346 ;
  assign n348 = ~n60 & ~n262 ;
  assign n349 = n319 & ~n348 ;
  assign n350 = x0 & ~n55 ;
  assign n351 = n161 & ~n350 ;
  assign n352 = ~n261 & ~n351 ;
  assign n353 = ~n349 & n352 ;
  assign n354 = ~x0 & ~n251 ;
  assign n355 = ~x2 & ~n354 ;
  assign n356 = ~n353 & n355 ;
  assign n357 = ~x3 & ~n335 ;
  assign n358 = n13 & n333 ;
  assign n359 = ~n297 & n358 ;
  assign n360 = n359 ^ x4 ;
  assign n361 = n359 ^ n23 ;
  assign n362 = n361 ^ n23 ;
  assign n363 = n362 ^ n360 ;
  assign n364 = ~x6 & n23 ;
  assign n365 = n364 ^ n336 ;
  assign n366 = n364 & n365 ;
  assign n367 = n366 ^ n23 ;
  assign n368 = n367 ^ n364 ;
  assign n369 = ~n363 & ~n368 ;
  assign n370 = n369 ^ n366 ;
  assign n371 = n370 ^ n364 ;
  assign n372 = n360 & n371 ;
  assign n373 = n372 ^ n359 ;
  assign n374 = n357 & ~n373 ;
  assign n375 = ~n356 & n374 ;
  assign n376 = x4 & n99 ;
  assign n377 = n24 & n376 ;
  assign n378 = n59 & n236 ;
  assign n379 = x7 ^ x4 ;
  assign n380 = n379 ^ x7 ;
  assign n381 = ~n55 & ~n87 ;
  assign n382 = n381 ^ x7 ;
  assign n383 = n380 & ~n382 ;
  assign n384 = n383 ^ x7 ;
  assign n385 = x2 & n384 ;
  assign n386 = ~n286 & n385 ;
  assign n387 = ~n378 & ~n386 ;
  assign n388 = x0 & ~n387 ;
  assign n389 = ~n377 & ~n388 ;
  assign n390 = ~x9 & ~n389 ;
  assign n391 = n262 & n376 ;
  assign n392 = x2 & ~n348 ;
  assign n393 = n392 ^ n55 ;
  assign n394 = n393 ^ x9 ;
  assign n395 = n394 ^ n392 ;
  assign n396 = n395 ^ n394 ;
  assign n397 = n297 ^ n205 ;
  assign n398 = x4 & n397 ;
  assign n399 = n398 ^ n297 ;
  assign n400 = n399 ^ n394 ;
  assign n401 = n400 ^ n393 ;
  assign n402 = n396 & ~n401 ;
  assign n403 = n402 ^ n399 ;
  assign n404 = x4 & ~n399 ;
  assign n405 = n404 ^ n393 ;
  assign n406 = ~n403 & ~n405 ;
  assign n407 = n406 ^ n404 ;
  assign n408 = ~n393 & n407 ;
  assign n409 = n408 ^ n402 ;
  assign n410 = n409 ^ n55 ;
  assign n411 = n410 ^ n399 ;
  assign n412 = ~n391 & n411 ;
  assign n413 = ~x0 & ~n412 ;
  assign n414 = x3 & ~n413 ;
  assign n415 = ~n390 & n414 ;
  assign n416 = ~n375 & ~n415 ;
  assign n417 = n11 & n311 ;
  assign n418 = n32 & n417 ;
  assign n419 = ~n416 & ~n418 ;
  assign n420 = n419 ^ x8 ;
  assign n421 = n420 ^ n419 ;
  assign n422 = ~x2 & n262 ;
  assign n423 = x6 & ~n327 ;
  assign n424 = n422 & n423 ;
  assign n425 = x2 & x7 ;
  assign n426 = n176 & n425 ;
  assign n427 = x6 ^ x3 ;
  assign n428 = n426 & n427 ;
  assign n429 = ~n424 & ~n428 ;
  assign n430 = n157 & n205 ;
  assign n431 = ~x0 & ~n430 ;
  assign n432 = n429 & n431 ;
  assign n433 = ~n309 & n432 ;
  assign n434 = n153 & n211 ;
  assign n435 = ~n206 & ~n434 ;
  assign n436 = ~x6 & ~n435 ;
  assign n437 = x2 & n436 ;
  assign n438 = n211 & n286 ;
  assign n439 = ~n159 & ~n438 ;
  assign n440 = n135 & ~n439 ;
  assign n441 = ~x6 & n156 ;
  assign n442 = n422 & n441 ;
  assign n443 = x0 & ~n442 ;
  assign n444 = ~n440 & n443 ;
  assign n445 = ~n437 & n444 ;
  assign n446 = x5 & ~n445 ;
  assign n447 = ~n433 & n446 ;
  assign n448 = n447 ^ n419 ;
  assign n449 = n421 & ~n448 ;
  assign n450 = n449 ^ n419 ;
  assign n451 = n347 & n450 ;
  assign n452 = ~n332 & n451 ;
  assign n453 = n452 ^ n281 ;
  assign n454 = n283 & n453 ;
  assign n455 = n454 ^ n281 ;
  assign n456 = n455 ^ n30 ;
  assign n457 = n152 & ~n456 ;
  assign n458 = n457 ^ n454 ;
  assign n459 = n458 ^ n281 ;
  assign n460 = n459 ^ n151 ;
  assign n461 = ~n30 & ~n460 ;
  assign n462 = n461 ^ n30 ;
  assign y0 = n462 ;
endmodule
