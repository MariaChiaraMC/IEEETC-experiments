module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n21 = x1 & x2 ;
  assign n22 = x0 & x2 ;
  assign n23 = ~n21 & ~n22 ;
  assign n24 = x5 & n23 ;
  assign n25 = ~x3 & n24 ;
  assign n26 = x6 & ~n25 ;
  assign n8 = x6 ^ x3 ;
  assign n9 = x6 ^ x1 ;
  assign n10 = n9 ^ x5 ;
  assign n11 = x6 ^ x2 ;
  assign n12 = n11 ^ x5 ;
  assign n13 = n10 & n12 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = ~x5 & ~x6 ;
  assign n16 = n15 ^ n8 ;
  assign n17 = ~n14 & n16 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n8 & n18 ;
  assign n20 = n19 ^ n8 ;
  assign n27 = n26 ^ n20 ;
  assign n28 = ~x4 & n27 ;
  assign n29 = n28 ^ n20 ;
  assign y0 = n29 ;
endmodule
