module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 ;
  assign n21 = ~x9 & ~x10 ;
  assign n31 = x8 & n21 ;
  assign n60 = ~x4 & n31 ;
  assign n12 = x0 & x2 ;
  assign n13 = x4 & x10 ;
  assign n14 = ~n12 & n13 ;
  assign n15 = n14 ^ x8 ;
  assign n16 = n14 ^ x9 ;
  assign n17 = n16 ^ x9 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = ~x2 & ~x5 ;
  assign n20 = x1 & n19 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n20 & n22 ;
  assign n24 = n23 ^ x9 ;
  assign n25 = n24 ^ n20 ;
  assign n26 = n18 & n25 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = n27 ^ n20 ;
  assign n29 = ~n15 & n28 ;
  assign n30 = n29 ^ n14 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = n32 ^ x6 ;
  assign n43 = n33 ^ n32 ;
  assign n34 = x6 & ~x10 ;
  assign n35 = ~x8 & ~n34 ;
  assign n36 = ~x4 & ~n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ n32 ;
  assign n39 = n33 ^ n30 ;
  assign n40 = n39 ^ n36 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n38 & n41 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = n44 ^ n38 ;
  assign n46 = x8 & x9 ;
  assign n47 = x2 & x4 ;
  assign n48 = ~n46 & ~n47 ;
  assign n49 = x0 & n21 ;
  assign n50 = n49 ^ x9 ;
  assign n51 = n48 & n50 ;
  assign n52 = n51 ^ n32 ;
  assign n53 = n42 ^ n38 ;
  assign n54 = n52 & n53 ;
  assign n55 = n54 ^ n32 ;
  assign n56 = ~n45 & n55 ;
  assign n57 = n56 ^ n32 ;
  assign n58 = n57 ^ n31 ;
  assign n59 = n58 ^ n32 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = n61 ^ n59 ;
  assign n63 = ~x6 & n19 ;
  assign n64 = n63 ^ n59 ;
  assign n65 = n64 ^ n59 ;
  assign n66 = n62 & n65 ;
  assign n67 = n66 ^ n59 ;
  assign n68 = x7 & n67 ;
  assign n69 = n68 ^ n59 ;
  assign n70 = ~x3 & n69 ;
  assign y0 = n70 ;
endmodule
