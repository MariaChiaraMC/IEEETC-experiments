module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 ;
  output y0 ;
  wire n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 ;
  assign n23 = x5 ^ x3 ;
  assign n26 = ~x0 & ~x2 ;
  assign n24 = x5 ^ x0 ;
  assign n25 = x5 & n24 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = n27 ^ x5 ;
  assign n29 = n26 ^ x1 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n30 ^ n23 ;
  assign n32 = n28 & n31 ;
  assign n33 = n32 ^ n25 ;
  assign n34 = n33 ^ x5 ;
  assign n35 = ~n23 & n34 ;
  assign n36 = ~x4 & n35 ;
  assign n225 = ~x19 & ~x20 ;
  assign n37 = ~x11 & x13 ;
  assign n38 = ~x6 & ~x7 ;
  assign n39 = ~x13 & ~n38 ;
  assign n40 = x9 & ~n39 ;
  assign n41 = ~n37 & n40 ;
  assign n42 = x11 ^ x10 ;
  assign n43 = n42 ^ n38 ;
  assign n44 = x16 ^ x15 ;
  assign n45 = x11 & n44 ;
  assign n46 = n45 ^ x15 ;
  assign n47 = n43 & n46 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = n48 ^ x15 ;
  assign n50 = n49 ^ x11 ;
  assign n51 = n38 & n50 ;
  assign n52 = ~n41 & ~n51 ;
  assign n53 = ~x8 & ~x15 ;
  assign n54 = x9 & x10 ;
  assign n55 = ~n53 & n54 ;
  assign n56 = ~x12 & n55 ;
  assign n57 = ~x10 & x11 ;
  assign n58 = ~x11 & ~x12 ;
  assign n59 = ~n57 & ~n58 ;
  assign n60 = x11 & ~x16 ;
  assign n61 = n53 & ~n60 ;
  assign n62 = ~n59 & n61 ;
  assign n63 = x13 & ~n62 ;
  assign n64 = x8 & n38 ;
  assign n65 = ~x17 & ~n64 ;
  assign n66 = x8 & x10 ;
  assign n67 = x7 & x11 ;
  assign n68 = n66 & n67 ;
  assign n69 = x6 & n68 ;
  assign n70 = n65 & ~n69 ;
  assign n71 = ~n63 & n70 ;
  assign n72 = ~n56 & n71 ;
  assign n73 = n72 ^ n52 ;
  assign n74 = x12 & ~x13 ;
  assign n75 = x7 & ~x16 ;
  assign n76 = n74 & ~n75 ;
  assign n77 = n76 ^ x6 ;
  assign n78 = n77 ^ n76 ;
  assign n79 = x11 & ~x12 ;
  assign n80 = x9 & n79 ;
  assign n81 = n80 ^ x12 ;
  assign n82 = x7 & n81 ;
  assign n83 = ~x13 & ~n82 ;
  assign n84 = n83 ^ n76 ;
  assign n85 = n78 & ~n84 ;
  assign n86 = n85 ^ n76 ;
  assign n87 = n86 ^ n52 ;
  assign n88 = n73 & ~n87 ;
  assign n89 = n88 ^ n85 ;
  assign n90 = n89 ^ n76 ;
  assign n91 = n90 ^ n72 ;
  assign n92 = n52 & ~n91 ;
  assign n93 = n92 ^ n52 ;
  assign n94 = x2 & ~n93 ;
  assign n95 = ~x9 & n58 ;
  assign n96 = ~x1 & ~n95 ;
  assign n97 = x13 & ~n96 ;
  assign n98 = ~x8 & x9 ;
  assign n99 = ~x10 & n98 ;
  assign n100 = n37 & n99 ;
  assign n101 = n54 & n79 ;
  assign n102 = ~x12 & x13 ;
  assign n103 = n67 & n102 ;
  assign n104 = ~n101 & ~n103 ;
  assign n105 = ~n100 & n104 ;
  assign n106 = n79 & n98 ;
  assign n107 = ~x1 & ~n106 ;
  assign n108 = ~x0 & ~n107 ;
  assign n109 = x4 & ~n108 ;
  assign n110 = n105 & n109 ;
  assign n111 = ~n97 & n110 ;
  assign n112 = ~n94 & n111 ;
  assign n113 = ~x3 & x5 ;
  assign n114 = ~x0 & x2 ;
  assign n115 = ~x4 & ~n114 ;
  assign n116 = n113 & ~n115 ;
  assign n117 = ~n112 & n116 ;
  assign n118 = x3 & ~x5 ;
  assign n119 = x2 & x21 ;
  assign n120 = n118 & ~n119 ;
  assign n121 = ~n114 & ~n120 ;
  assign n122 = x1 & x4 ;
  assign n123 = ~n121 & n122 ;
  assign n124 = x0 & ~x1 ;
  assign n125 = x5 ^ x4 ;
  assign n126 = n125 ^ n124 ;
  assign n127 = ~x12 & ~x13 ;
  assign n128 = x9 & n127 ;
  assign n129 = n64 & n128 ;
  assign n130 = n129 ^ x3 ;
  assign n131 = n130 ^ n129 ;
  assign n132 = n129 ^ x2 ;
  assign n133 = ~n131 & n132 ;
  assign n134 = n133 ^ n129 ;
  assign n135 = ~x8 & ~x9 ;
  assign n136 = ~n129 & ~n135 ;
  assign n137 = n136 ^ n57 ;
  assign n138 = ~n134 & n137 ;
  assign n139 = n138 ^ n136 ;
  assign n140 = n57 & n139 ;
  assign n141 = n140 ^ n57 ;
  assign n142 = n141 ^ x3 ;
  assign n143 = x4 & n142 ;
  assign n144 = n143 ^ n141 ;
  assign n145 = ~n126 & n144 ;
  assign n146 = n145 ^ n143 ;
  assign n147 = n146 ^ n141 ;
  assign n148 = n147 ^ x4 ;
  assign n149 = n124 & n148 ;
  assign n150 = ~n123 & ~n149 ;
  assign n151 = n57 & n64 ;
  assign n152 = x1 & x2 ;
  assign n153 = ~x3 & n152 ;
  assign n154 = ~x5 & n26 ;
  assign n155 = ~n153 & ~n154 ;
  assign n156 = n151 & ~n155 ;
  assign n157 = ~x8 & n38 ;
  assign n158 = ~x11 & n157 ;
  assign n159 = ~x11 & n66 ;
  assign n160 = ~n158 & ~n159 ;
  assign n161 = n154 & n157 ;
  assign n162 = x3 ^ x1 ;
  assign n163 = x0 & ~x5 ;
  assign n164 = n163 ^ x3 ;
  assign n165 = x3 ^ x2 ;
  assign n166 = n165 ^ n163 ;
  assign n167 = n163 & n166 ;
  assign n168 = n167 ^ n163 ;
  assign n169 = ~n164 & n168 ;
  assign n170 = n169 ^ n167 ;
  assign n171 = n170 ^ n163 ;
  assign n172 = n171 ^ n165 ;
  assign n173 = ~n162 & n172 ;
  assign n174 = n173 ^ n165 ;
  assign n175 = ~n161 & ~n174 ;
  assign n176 = ~n160 & ~n175 ;
  assign n177 = ~n156 & ~n176 ;
  assign n178 = n128 & ~n177 ;
  assign n180 = x10 & n158 ;
  assign n181 = n127 & n180 ;
  assign n179 = ~x1 & n26 ;
  assign n182 = n181 ^ n179 ;
  assign n183 = n179 ^ n153 ;
  assign n184 = n183 ^ n153 ;
  assign n185 = n153 ^ x3 ;
  assign n186 = n184 & n185 ;
  assign n187 = n186 ^ n153 ;
  assign n188 = n182 & ~n187 ;
  assign n189 = n188 ^ n181 ;
  assign n190 = ~n178 & ~n189 ;
  assign n191 = ~x4 & ~n190 ;
  assign n192 = x3 & ~x4 ;
  assign n193 = ~n151 & n160 ;
  assign n194 = n128 & ~n193 ;
  assign n195 = n57 & n135 ;
  assign n196 = ~n39 & n195 ;
  assign n197 = ~n74 & n196 ;
  assign n198 = ~n181 & ~n197 ;
  assign n199 = ~n194 & n198 ;
  assign n200 = n192 & ~n199 ;
  assign n201 = ~x3 & ~n102 ;
  assign n202 = ~x1 & ~n201 ;
  assign n203 = n202 ^ x4 ;
  assign n204 = x3 ^ x0 ;
  assign n205 = n204 ^ x0 ;
  assign n206 = n128 ^ x0 ;
  assign n207 = n205 & n206 ;
  assign n208 = n207 ^ x0 ;
  assign n209 = n208 ^ n202 ;
  assign n210 = n203 & ~n209 ;
  assign n211 = n210 ^ n207 ;
  assign n212 = n211 ^ x0 ;
  assign n213 = n212 ^ x4 ;
  assign n214 = ~n202 & ~n213 ;
  assign n215 = n214 ^ n202 ;
  assign n216 = n215 ^ n202 ;
  assign n217 = n216 ^ x1 ;
  assign n218 = ~x2 & ~n217 ;
  assign n219 = n218 ^ x1 ;
  assign n220 = ~n200 & ~n219 ;
  assign n221 = x5 & ~n220 ;
  assign n222 = ~n191 & ~n221 ;
  assign n223 = n150 & n222 ;
  assign n224 = ~n117 & n223 ;
  assign n226 = n225 ^ n224 ;
  assign n227 = n226 ^ n224 ;
  assign n228 = n224 ^ x18 ;
  assign n229 = ~n227 & n228 ;
  assign n230 = n229 ^ n224 ;
  assign n231 = ~n36 & n230 ;
  assign n232 = x14 & ~n231 ;
  assign y0 = n232 ;
endmodule
