module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n8 = x0 & ~x6 ;
  assign n9 = x5 & ~n8 ;
  assign n10 = x4 & ~n9 ;
  assign n11 = x1 & x3 ;
  assign n12 = ~n10 & n11 ;
  assign n13 = n12 ^ x2 ;
  assign n19 = n13 ^ n12 ;
  assign n14 = n13 ^ x4 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = x4 ^ x0 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = ~n15 & n17 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = n20 ^ n15 ;
  assign n22 = n12 ^ x3 ;
  assign n23 = n18 ^ n15 ;
  assign n24 = ~n22 & ~n23 ;
  assign n25 = n24 ^ n12 ;
  assign n26 = n21 & n25 ;
  assign n27 = n26 ^ n12 ;
  assign n28 = n27 ^ n12 ;
  assign y0 = n28 ;
endmodule
