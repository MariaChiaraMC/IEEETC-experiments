// Benchmark "restrictions/spla.pla.uscita15.plaopt.pla_res_0" written by ABC on Mon Jun 28 06:10:30 2021

module \restrictions/spla.pla.uscita15.plaopt.pla_res_0  ( 
    x0, x1,
    z0  );
  input  x0, x1;
  output z0;
  assign z0 = ~x0 | x1;
endmodule


