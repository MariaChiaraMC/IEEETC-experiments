// Benchmark "./pla/f51m.pla_res_7NonExact" written by ABC on Fri Nov 20 10:22:17 2020

module \./pla/f51m.pla_res_7NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = ~x0;
endmodule


