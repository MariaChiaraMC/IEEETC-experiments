module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n13 = x6 & ~x9 ;
  assign n14 = ~x8 & ~x10 ;
  assign n15 = ~n13 & ~n14 ;
  assign n16 = ~x7 & ~n15 ;
  assign n17 = ~x0 & n16 ;
  assign n18 = x11 ^ x6 ;
  assign n19 = n18 ^ n17 ;
  assign n21 = x2 & ~x5 ;
  assign n22 = x3 & ~n21 ;
  assign n23 = ~x4 & ~x9 ;
  assign n24 = n22 & n23 ;
  assign n25 = x1 & n24 ;
  assign n20 = x8 & x10 ;
  assign n26 = n25 ^ n20 ;
  assign n27 = ~x11 & n26 ;
  assign n28 = n27 ^ n20 ;
  assign n29 = ~n19 & ~n28 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n30 ^ n20 ;
  assign n32 = n31 ^ x11 ;
  assign n33 = n17 & n32 ;
  assign y0 = n33 ;
endmodule
