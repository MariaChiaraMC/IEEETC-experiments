module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 ;
  assign n22 = ~x0 & ~x2 ;
  assign n23 = ~x3 & ~x4 ;
  assign n24 = x1 & n23 ;
  assign n25 = n22 & n24 ;
  assign n26 = ~x1 & x3 ;
  assign n27 = ~n22 & ~n26 ;
  assign n28 = ~x1 & x2 ;
  assign n29 = n27 & ~n28 ;
  assign n30 = ~x0 & ~x1 ;
  assign n31 = ~x4 & ~n30 ;
  assign n32 = x5 & n31 ;
  assign n33 = ~n29 & n32 ;
  assign n34 = n33 ^ x14 ;
  assign n228 = ~x19 & ~x20 ;
  assign n35 = x3 & x4 ;
  assign n36 = n35 ^ x2 ;
  assign n37 = n36 ^ x5 ;
  assign n76 = n37 ^ x1 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = n38 ^ n37 ;
  assign n75 = n39 ^ x1 ;
  assign n77 = n76 ^ n75 ;
  assign n41 = ~x12 & ~x13 ;
  assign n47 = ~x6 & ~x7 ;
  assign n42 = ~x8 & ~x11 ;
  assign n43 = ~x9 & ~x10 ;
  assign n44 = n42 & ~n43 ;
  assign n48 = n47 ^ n44 ;
  assign n57 = n48 ^ n44 ;
  assign n45 = x8 & x9 ;
  assign n46 = n45 ^ n44 ;
  assign n49 = n48 ^ n46 ;
  assign n50 = n49 ^ n48 ;
  assign n51 = n50 ^ n44 ;
  assign n52 = n49 ^ x11 ;
  assign n53 = n52 ^ x10 ;
  assign n54 = n53 ^ n49 ;
  assign n55 = n54 ^ n51 ;
  assign n56 = n51 & n55 ;
  assign n58 = n57 ^ n56 ;
  assign n59 = n58 ^ n51 ;
  assign n60 = n44 ^ x10 ;
  assign n61 = n56 ^ n51 ;
  assign n62 = ~n60 & n61 ;
  assign n63 = n62 ^ n44 ;
  assign n64 = n59 & ~n63 ;
  assign n65 = n64 ^ n44 ;
  assign n66 = n65 ^ n47 ;
  assign n67 = n66 ^ n44 ;
  assign n68 = n23 & n67 ;
  assign n69 = n41 & n68 ;
  assign n70 = n69 ^ n38 ;
  assign n40 = n39 ^ n36 ;
  assign n71 = n70 ^ n40 ;
  assign n72 = n40 ^ x1 ;
  assign n73 = n71 & ~n72 ;
  assign n74 = n73 ^ x1 ;
  assign n78 = n77 ^ n74 ;
  assign n79 = n78 ^ n70 ;
  assign n80 = n77 ^ n76 ;
  assign n81 = n80 ^ n40 ;
  assign n82 = ~n76 & ~n81 ;
  assign n83 = ~x0 & x4 ;
  assign n84 = n76 ^ n70 ;
  assign n85 = n83 & ~n84 ;
  assign n86 = n85 ^ n83 ;
  assign n87 = n86 ^ n70 ;
  assign n88 = n87 ^ n40 ;
  assign n89 = n82 & n88 ;
  assign n90 = n89 ^ x1 ;
  assign n91 = ~n79 & ~n90 ;
  assign n92 = n91 ^ n82 ;
  assign n93 = n92 ^ n89 ;
  assign n94 = n93 ^ x1 ;
  assign n95 = n94 ^ n76 ;
  assign n96 = n95 ^ n77 ;
  assign n97 = n96 ^ x2 ;
  assign n98 = n97 ^ n39 ;
  assign n99 = ~n30 & n98 ;
  assign n100 = ~x9 & ~n30 ;
  assign n101 = ~x2 & n26 ;
  assign n102 = ~n22 & ~n101 ;
  assign n103 = ~n100 & ~n102 ;
  assign n104 = ~x5 & ~n103 ;
  assign n105 = n43 ^ x11 ;
  assign n106 = x13 ^ x5 ;
  assign n107 = n43 ^ x5 ;
  assign n108 = n107 ^ x5 ;
  assign n109 = ~n106 & ~n108 ;
  assign n110 = n109 ^ x5 ;
  assign n111 = ~n105 & n110 ;
  assign n112 = ~x8 & n111 ;
  assign n113 = x12 & ~x13 ;
  assign n114 = ~x13 & ~n47 ;
  assign n115 = ~n113 & ~n114 ;
  assign n116 = n112 & n115 ;
  assign n117 = ~n104 & n116 ;
  assign n128 = ~x10 & x11 ;
  assign n129 = n47 & n128 ;
  assign n130 = ~n27 & n129 ;
  assign n118 = x8 ^ x5 ;
  assign n120 = n118 ^ x2 ;
  assign n119 = n118 ^ x8 ;
  assign n121 = n120 ^ n119 ;
  assign n131 = n130 ^ n121 ;
  assign n135 = n131 ^ n120 ;
  assign n136 = n135 ^ n118 ;
  assign n122 = n121 ^ n120 ;
  assign n123 = n122 ^ n118 ;
  assign n124 = n123 ^ n118 ;
  assign n125 = n120 ^ n101 ;
  assign n126 = n125 ^ n118 ;
  assign n127 = ~n124 & ~n126 ;
  assign n132 = n131 ^ n127 ;
  assign n133 = n132 ^ n118 ;
  assign n134 = ~n123 & ~n133 ;
  assign n137 = n136 ^ n134 ;
  assign n138 = n137 ^ n123 ;
  assign n139 = x10 & ~x11 ;
  assign n140 = n139 ^ n118 ;
  assign n141 = n136 ^ n133 ;
  assign n142 = n141 ^ n123 ;
  assign n143 = ~n140 & ~n142 ;
  assign n144 = n143 ^ n118 ;
  assign n145 = n138 & n144 ;
  assign n146 = n145 ^ n143 ;
  assign n147 = n146 ^ n118 ;
  assign n148 = n147 ^ x8 ;
  assign n149 = n41 & n148 ;
  assign n150 = x9 & n149 ;
  assign n151 = ~n117 & ~n150 ;
  assign n152 = ~x4 & ~n151 ;
  assign n153 = ~n99 & ~n152 ;
  assign n154 = x9 & ~x10 ;
  assign n155 = n42 & n154 ;
  assign n156 = x15 ^ x12 ;
  assign n157 = x2 & ~n156 ;
  assign n158 = n157 ^ x12 ;
  assign n159 = ~n155 & n158 ;
  assign n160 = ~x1 & n159 ;
  assign n161 = x13 & ~n160 ;
  assign n162 = x9 & ~x12 ;
  assign n163 = x11 & n162 ;
  assign n164 = x10 & n163 ;
  assign n165 = ~x2 & ~n164 ;
  assign n166 = ~x8 & ~x9 ;
  assign n167 = ~x17 & ~n113 ;
  assign n168 = n166 & n167 ;
  assign n169 = n129 & n168 ;
  assign n170 = x16 & n169 ;
  assign n171 = ~n165 & ~n170 ;
  assign n172 = ~x0 & x1 ;
  assign n173 = x4 & ~n172 ;
  assign n174 = ~n171 & n173 ;
  assign n175 = ~n161 & n174 ;
  assign n176 = x5 & ~n175 ;
  assign n177 = ~x8 & n163 ;
  assign n178 = x5 & n177 ;
  assign n179 = n178 ^ x1 ;
  assign n180 = n179 ^ n178 ;
  assign n181 = n178 ^ x4 ;
  assign n182 = n181 ^ n179 ;
  assign n183 = n182 ^ x0 ;
  assign n188 = n183 ^ n179 ;
  assign n189 = n188 ^ n178 ;
  assign n190 = n189 ^ n178 ;
  assign n184 = n183 ^ x0 ;
  assign n185 = n184 ^ n179 ;
  assign n186 = n185 ^ n178 ;
  assign n187 = n186 ^ n180 ;
  assign n191 = n190 ^ n187 ;
  assign n192 = n180 & n191 ;
  assign n193 = n192 ^ n189 ;
  assign n194 = n193 ^ n180 ;
  assign n195 = n194 ^ n190 ;
  assign n196 = n128 & n166 ;
  assign n197 = n183 ^ x2 ;
  assign n198 = n197 ^ x0 ;
  assign n199 = n198 ^ n180 ;
  assign n200 = ~n196 & ~n199 ;
  assign n201 = n200 ^ n186 ;
  assign n202 = n196 ^ n189 ;
  assign n203 = n196 ^ n186 ;
  assign n204 = ~n202 & n203 ;
  assign n205 = n204 ^ n189 ;
  assign n206 = n205 ^ n180 ;
  assign n207 = n206 ^ n198 ;
  assign n208 = n207 ^ n186 ;
  assign n209 = ~n201 & n208 ;
  assign n210 = n209 ^ n189 ;
  assign n211 = n210 ^ n180 ;
  assign n212 = ~n195 & n211 ;
  assign n213 = n212 ^ x1 ;
  assign n214 = ~n176 & n213 ;
  assign n215 = n214 ^ x3 ;
  assign n216 = n215 ^ n214 ;
  assign n217 = n216 ^ n153 ;
  assign n218 = ~x2 & x5 ;
  assign n219 = n218 ^ x1 ;
  assign n220 = n218 & ~n219 ;
  assign n221 = n220 ^ n214 ;
  assign n222 = n221 ^ n218 ;
  assign n223 = n217 & ~n222 ;
  assign n224 = n223 ^ n220 ;
  assign n225 = n224 ^ n218 ;
  assign n226 = n153 & n225 ;
  assign n227 = n226 ^ n153 ;
  assign n229 = n228 ^ n227 ;
  assign n230 = n229 ^ n227 ;
  assign n231 = n227 ^ x18 ;
  assign n232 = ~n230 & n231 ;
  assign n233 = n232 ^ n227 ;
  assign n234 = n233 ^ n33 ;
  assign n235 = ~n34 & ~n234 ;
  assign n236 = n235 ^ n232 ;
  assign n237 = n236 ^ n227 ;
  assign n238 = n237 ^ x14 ;
  assign n239 = ~n33 & n238 ;
  assign n240 = n239 ^ n33 ;
  assign n241 = ~n25 & ~n240 ;
  assign y0 = ~n241 ;
endmodule
