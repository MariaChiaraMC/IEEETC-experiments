module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 ;
  assign n25 = ~x1 & x2 ;
  assign n18 = ~x4 & ~x6 ;
  assign n26 = x14 & n18 ;
  assign n27 = n25 & ~n26 ;
  assign n28 = x7 & x10 ;
  assign n29 = n28 ^ x2 ;
  assign n30 = n28 ^ x6 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = x9 ^ x1 ;
  assign n33 = x6 & ~n32 ;
  assign n34 = n33 ^ x1 ;
  assign n35 = ~n31 & ~n34 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = n36 ^ x1 ;
  assign n38 = n37 ^ x6 ;
  assign n39 = n29 & ~n38 ;
  assign n40 = n39 ^ x2 ;
  assign n41 = ~n27 & n40 ;
  assign n16 = ~x9 & ~x10 ;
  assign n17 = ~x7 & n16 ;
  assign n19 = ~x1 & ~x2 ;
  assign n20 = n18 & n19 ;
  assign n21 = n17 & n20 ;
  assign n42 = n41 ^ n21 ;
  assign n43 = n42 ^ n21 ;
  assign n22 = x1 & ~x9 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n23 ^ n21 ;
  assign n44 = n43 ^ n24 ;
  assign n45 = x4 & ~x14 ;
  assign n46 = ~n25 & ~n45 ;
  assign n47 = n46 ^ n21 ;
  assign n48 = n47 ^ n21 ;
  assign n49 = n48 ^ n43 ;
  assign n50 = n43 & ~n49 ;
  assign n51 = n50 ^ n43 ;
  assign n52 = ~n44 & n51 ;
  assign n53 = n52 ^ n50 ;
  assign n54 = n53 ^ n21 ;
  assign n55 = n54 ^ n43 ;
  assign n56 = x3 & n55 ;
  assign n57 = n56 ^ n21 ;
  assign n58 = ~x5 & n57 ;
  assign n59 = x2 & x3 ;
  assign n60 = n45 & n59 ;
  assign n61 = x1 & ~x6 ;
  assign n62 = x1 & ~x10 ;
  assign n63 = ~n61 & ~n62 ;
  assign n64 = ~x7 & ~n63 ;
  assign n65 = n60 & n64 ;
  assign n66 = x9 & n65 ;
  assign n67 = ~n58 & ~n66 ;
  assign n68 = ~x12 & ~n67 ;
  assign n69 = n68 ^ x14 ;
  assign n70 = n68 ^ x13 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = ~n69 & ~n71 ;
  assign n73 = n72 ^ n68 ;
  assign n74 = n73 ^ n69 ;
  assign n75 = n68 ^ x10 ;
  assign n76 = n75 ^ n70 ;
  assign n77 = n76 ^ x12 ;
  assign n78 = n77 ^ x14 ;
  assign n79 = n78 ^ n76 ;
  assign n80 = ~x3 & n25 ;
  assign n81 = x5 & ~x6 ;
  assign n82 = x4 & x9 ;
  assign n83 = n81 & n82 ;
  assign n84 = n80 & n83 ;
  assign n85 = n84 ^ n76 ;
  assign n86 = n85 ^ n76 ;
  assign n87 = n76 ^ n70 ;
  assign n88 = n87 ^ n68 ;
  assign n89 = n86 & n88 ;
  assign n90 = n89 ^ n72 ;
  assign n91 = n90 ^ n68 ;
  assign n92 = n91 ^ n69 ;
  assign n93 = n79 & ~n92 ;
  assign n94 = n93 ^ n71 ;
  assign n95 = ~n74 & ~n94 ;
  assign n96 = n95 ^ n93 ;
  assign n97 = n96 ^ n68 ;
  assign n98 = n97 ^ n71 ;
  assign n99 = n98 ^ x13 ;
  assign n100 = n99 ^ n68 ;
  assign n101 = ~x0 & n100 ;
  assign n102 = ~x4 & ~x5 ;
  assign n103 = n16 & n102 ;
  assign n104 = x7 & ~x14 ;
  assign n105 = x12 & x13 ;
  assign n106 = n104 & n105 ;
  assign n107 = ~x2 & x3 ;
  assign n108 = x0 & x6 ;
  assign n109 = ~n107 & n108 ;
  assign n110 = n106 & n109 ;
  assign n111 = n103 & n110 ;
  assign n112 = ~n80 & n111 ;
  assign n113 = ~n101 & ~n112 ;
  assign n114 = ~x8 & ~n113 ;
  assign n115 = ~x11 & n114 ;
  assign y0 = n115 ;
endmodule
