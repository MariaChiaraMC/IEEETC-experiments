module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 ;
  assign n17 = ~x1 & x4 ;
  assign n18 = x5 & n17 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = n19 ^ x0 ;
  assign n107 = n20 ^ n19 ;
  assign n23 = x12 & ~x13 ;
  assign n24 = x14 & ~x15 ;
  assign n25 = ~n23 & ~n24 ;
  assign n21 = ~x0 & ~x5 ;
  assign n26 = x6 & x7 ;
  assign n27 = n21 & ~n26 ;
  assign n28 = x5 & x7 ;
  assign n29 = ~n27 & ~n28 ;
  assign n30 = ~x8 & ~x9 ;
  assign n31 = x8 & x9 ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = n21 & n32 ;
  assign n34 = n33 ^ x10 ;
  assign n35 = n34 ^ n33 ;
  assign n36 = x5 & x6 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n35 & n37 ;
  assign n39 = n38 ^ n33 ;
  assign n40 = ~x11 & n39 ;
  assign n41 = n29 & ~n40 ;
  assign n42 = ~n25 & ~n41 ;
  assign n43 = x15 ^ x13 ;
  assign n44 = n36 & n43 ;
  assign n45 = x12 & x14 ;
  assign n46 = ~x10 & x11 ;
  assign n47 = n45 & n46 ;
  assign n48 = n44 & n47 ;
  assign n49 = ~n42 & ~n48 ;
  assign n22 = x6 & n21 ;
  assign n50 = n49 ^ n22 ;
  assign n51 = n50 ^ x1 ;
  assign n89 = n51 ^ n50 ;
  assign n52 = ~x11 & ~x12 ;
  assign n53 = ~x13 & ~x15 ;
  assign n54 = n53 ^ x8 ;
  assign n55 = n54 ^ x14 ;
  assign n62 = n55 ^ n53 ;
  assign n56 = n55 ^ x1 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = x14 ^ x1 ;
  assign n59 = n58 ^ x1 ;
  assign n60 = n59 ^ n57 ;
  assign n61 = n57 & ~n60 ;
  assign n63 = n62 ^ n61 ;
  assign n64 = n63 ^ n57 ;
  assign n65 = n53 ^ n43 ;
  assign n66 = n61 ^ n57 ;
  assign n67 = n65 & n66 ;
  assign n68 = n67 ^ n53 ;
  assign n69 = n64 & n68 ;
  assign n70 = n69 ^ n53 ;
  assign n71 = n70 ^ n53 ;
  assign n72 = n52 & n71 ;
  assign n73 = x7 & x14 ;
  assign n74 = n73 ^ x9 ;
  assign n75 = n74 ^ x9 ;
  assign n76 = n31 ^ x9 ;
  assign n77 = n76 ^ x9 ;
  assign n78 = ~n75 & ~n77 ;
  assign n79 = n78 ^ x9 ;
  assign n80 = x10 & n79 ;
  assign n81 = n80 ^ x9 ;
  assign n82 = n72 & n81 ;
  assign n83 = n82 ^ n51 ;
  assign n84 = n83 ^ n50 ;
  assign n85 = n82 ^ n22 ;
  assign n86 = n85 ^ n82 ;
  assign n87 = n86 ^ n84 ;
  assign n88 = n84 & n87 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = n90 ^ n84 ;
  assign n92 = n50 ^ x7 ;
  assign n93 = n88 ^ n84 ;
  assign n94 = n92 & n93 ;
  assign n95 = n94 ^ n50 ;
  assign n96 = ~n91 & ~n95 ;
  assign n97 = n96 ^ n50 ;
  assign n98 = n97 ^ n22 ;
  assign n99 = n98 ^ n50 ;
  assign n100 = x4 & n99 ;
  assign n101 = n100 ^ n20 ;
  assign n102 = n101 ^ n19 ;
  assign n103 = n20 ^ n18 ;
  assign n104 = n103 ^ n100 ;
  assign n105 = n104 ^ n102 ;
  assign n106 = ~n102 & n105 ;
  assign n108 = n107 ^ n106 ;
  assign n109 = n108 ^ n102 ;
  assign n110 = ~x4 & ~x7 ;
  assign n111 = ~x6 & x7 ;
  assign n112 = n30 & n111 ;
  assign n113 = n46 & n112 ;
  assign n114 = ~n110 & ~n113 ;
  assign n115 = x5 & ~n114 ;
  assign n116 = ~n25 & n115 ;
  assign n120 = ~x6 & ~n32 ;
  assign n121 = n28 & ~n120 ;
  assign n117 = ~x4 & ~x5 ;
  assign n118 = x7 ^ x6 ;
  assign n119 = n117 & n118 ;
  assign n122 = n121 ^ n119 ;
  assign n123 = n122 ^ x10 ;
  assign n130 = n123 ^ n122 ;
  assign n124 = n123 ^ n25 ;
  assign n125 = n124 ^ n122 ;
  assign n126 = n119 ^ n25 ;
  assign n127 = n126 ^ n25 ;
  assign n128 = n127 ^ n125 ;
  assign n129 = n125 & ~n128 ;
  assign n131 = n130 ^ n129 ;
  assign n132 = n131 ^ n125 ;
  assign n133 = n122 ^ n112 ;
  assign n134 = n129 ^ n125 ;
  assign n135 = n133 & n134 ;
  assign n136 = n135 ^ n122 ;
  assign n137 = ~n132 & n136 ;
  assign n138 = n137 ^ n122 ;
  assign n139 = n138 ^ n119 ;
  assign n140 = n139 ^ n122 ;
  assign n141 = ~x11 & n140 ;
  assign n142 = ~n116 & ~n141 ;
  assign n143 = ~x1 & ~n142 ;
  assign n144 = n143 ^ n19 ;
  assign n145 = n106 ^ n102 ;
  assign n146 = n144 & ~n145 ;
  assign n147 = n146 ^ n19 ;
  assign n148 = ~n109 & ~n147 ;
  assign n149 = n148 ^ n19 ;
  assign n150 = n149 ^ x2 ;
  assign n151 = n150 ^ n19 ;
  assign n152 = ~x3 & ~n151 ;
  assign y0 = n152 ;
endmodule
