module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 ;
  assign n13 = x1 ^ x0 ;
  assign n15 = x5 & ~x6 ;
  assign n16 = ~x8 & n15 ;
  assign n26 = ~x7 & x9 ;
  assign n27 = n16 & n26 ;
  assign n14 = x4 & x7 ;
  assign n17 = x3 & ~x9 ;
  assign n18 = n16 & n17 ;
  assign n19 = x8 & ~x10 ;
  assign n20 = x9 & n19 ;
  assign n21 = ~x3 & ~x5 ;
  assign n22 = n20 & n21 ;
  assign n23 = x6 & n22 ;
  assign n24 = ~n18 & ~n23 ;
  assign n25 = n14 & ~n24 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = x2 & n28 ;
  assign n30 = n28 ^ n25 ;
  assign n31 = ~x4 & ~x10 ;
  assign n32 = x3 & ~n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = ~n30 & n33 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = n29 & n35 ;
  assign n37 = n36 ^ n27 ;
  assign n38 = n37 ^ x11 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = n14 & n15 ;
  assign n41 = ~x2 & n20 ;
  assign n42 = n40 & n41 ;
  assign n43 = n42 ^ n37 ;
  assign n44 = n39 & n43 ;
  assign n45 = n44 ^ n37 ;
  assign n46 = n45 ^ x1 ;
  assign n47 = n13 & n46 ;
  assign n48 = n47 ^ n44 ;
  assign n49 = n48 ^ n37 ;
  assign n50 = n49 ^ x0 ;
  assign n51 = x1 & n50 ;
  assign n52 = n51 ^ x1 ;
  assign y0 = n52 ;
endmodule
