module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n17 = ~x0 & ~x3 ;
  assign n18 = ~x6 & n17 ;
  assign n19 = ~x4 & n18 ;
  assign n20 = x10 ^ x9 ;
  assign n21 = n20 ^ x11 ;
  assign n22 = n21 ^ x8 ;
  assign n23 = ~x1 & ~x2 ;
  assign n24 = x5 & x7 ;
  assign n25 = n23 & n24 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = x11 ^ x10 ;
  assign n28 = x10 ^ x8 ;
  assign n29 = n27 & n28 ;
  assign n30 = n29 ^ x10 ;
  assign n31 = n30 ^ n22 ;
  assign n32 = n26 & ~n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ x10 ;
  assign n35 = n34 ^ n25 ;
  assign n36 = n22 & ~n35 ;
  assign n37 = n36 ^ n22 ;
  assign n38 = n19 & n37 ;
  assign y0 = n38 ;
endmodule
