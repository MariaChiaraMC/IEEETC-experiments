module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n8 = x5 ^ x4 ;
  assign n9 = n8 ^ x5 ;
  assign n10 = n9 ^ x6 ;
  assign n12 = ~x1 & ~x3 ;
  assign n15 = ~x2 & n12 ;
  assign n11 = ~x2 & ~x3 ;
  assign n13 = ~x0 & n12 ;
  assign n14 = ~n11 & ~n13 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n16 ^ n9 ;
  assign n18 = x5 & ~n17 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n19 ^ x5 ;
  assign n21 = n20 ^ n9 ;
  assign n22 = n21 ^ x6 ;
  assign n23 = n10 & ~n22 ;
  assign n24 = n23 ^ n18 ;
  assign n25 = n24 ^ n15 ;
  assign n26 = n25 ^ n9 ;
  assign n27 = x6 & ~n26 ;
  assign n28 = n27 ^ x6 ;
  assign n29 = n28 ^ x6 ;
  assign n30 = n29 ^ x6 ;
  assign y0 = ~n30 ;
endmodule
