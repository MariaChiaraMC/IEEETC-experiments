// Benchmark "./m4.pla" written by ABC on Thu Apr 23 10:59:56 2020

module \./m4.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z8  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z8;
  assign z8 = 1'b1;
endmodule


