module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n15 = ~x5 & ~x9 ;
  assign n16 = ~x12 & ~x13 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = ~x6 & x10 ;
  assign n19 = n18 ^ x11 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = x3 & ~x10 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = ~n20 & n22 ;
  assign n24 = n23 ^ n18 ;
  assign n25 = n24 ^ n15 ;
  assign n26 = n17 & n25 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = n27 ^ n18 ;
  assign n29 = n28 ^ n16 ;
  assign n30 = n15 & n29 ;
  assign n31 = n30 ^ n15 ;
  assign y0 = n31 ;
endmodule
