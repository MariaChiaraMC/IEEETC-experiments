module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n9 = ~x2 & x7 ;
  assign n10 = n9 ^ x6 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = x4 & x5 ;
  assign n13 = x2 & ~n12 ;
  assign n14 = n13 ^ n9 ;
  assign n15 = n14 ^ n9 ;
  assign n16 = ~n11 & ~n15 ;
  assign n17 = n16 ^ n9 ;
  assign n18 = x1 & n17 ;
  assign n19 = n18 ^ n9 ;
  assign n20 = x0 & n19 ;
  assign n21 = ~x1 & x5 ;
  assign n22 = ~x2 & ~n21 ;
  assign n23 = x3 & ~n22 ;
  assign n24 = x1 ^ x0 ;
  assign n25 = n23 & ~n24 ;
  assign n26 = ~x2 & ~x3 ;
  assign n27 = n26 ^ x4 ;
  assign n29 = ~x0 & ~x1 ;
  assign n28 = x0 & x1 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = n29 ^ n26 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = n30 & n32 ;
  assign n34 = n33 ^ n29 ;
  assign n35 = n27 & ~n34 ;
  assign n36 = n35 ^ x4 ;
  assign n37 = ~n25 & ~n36 ;
  assign n38 = ~n20 & n37 ;
  assign y0 = ~n38 ;
endmodule
