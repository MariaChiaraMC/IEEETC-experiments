module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 ;
  assign n12 = x8 & x9 ;
  assign n13 = ~x2 & x10 ;
  assign n14 = n12 & n13 ;
  assign n15 = n14 ^ x6 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = x3 & x4 ;
  assign n18 = x1 & ~n17 ;
  assign n19 = ~x5 & ~n18 ;
  assign n20 = n14 & ~n19 ;
  assign n21 = ~x7 & n20 ;
  assign n22 = n21 ^ n14 ;
  assign n23 = ~n16 & ~n22 ;
  assign n24 = n23 ^ n14 ;
  assign n25 = ~x0 & ~n24 ;
  assign y0 = n25 ;
endmodule
