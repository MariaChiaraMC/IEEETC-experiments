module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
  assign n11 = x4 & x5 ;
  assign n12 = ~x3 & ~n11 ;
  assign n13 = ~x4 & ~x5 ;
  assign n14 = ~x1 & n13 ;
  assign n15 = n14 ^ x2 ;
  assign n16 = n14 ^ x0 ;
  assign n17 = ~n15 & ~n16 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = ~x7 & ~x8 ;
  assign n20 = ~n14 & ~n19 ;
  assign n21 = n20 ^ x6 ;
  assign n22 = ~n18 & ~n21 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = ~x6 & n23 ;
  assign n25 = n24 ^ x6 ;
  assign n26 = n12 & ~n25 ;
  assign n27 = n13 ^ x1 ;
  assign n28 = ~x0 & ~x2 ;
  assign n29 = ~x8 & x9 ;
  assign n30 = ~n19 & ~n29 ;
  assign n31 = ~n28 & n30 ;
  assign n32 = n13 & n31 ;
  assign n33 = n27 & n32 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = n26 & ~n34 ;
  assign y0 = n35 ;
endmodule
