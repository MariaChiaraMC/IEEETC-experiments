module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n7 = x5 ^ x4 ;
  assign n11 = n7 ^ x5 ;
  assign n9 = x5 ^ x1 ;
  assign n8 = n7 ^ x3 ;
  assign n10 = n9 ^ n8 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = n11 ^ x5 ;
  assign n14 = ~n12 & ~n13 ;
  assign n15 = n14 ^ n9 ;
  assign n16 = n15 ^ x5 ;
  assign n18 = n10 ^ n9 ;
  assign n19 = n18 ^ x5 ;
  assign n20 = ~n18 & ~n19 ;
  assign n17 = ~x0 & ~x2 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n21 ^ n9 ;
  assign n23 = n22 ^ n10 ;
  assign n24 = ~n11 & ~n23 ;
  assign n25 = n24 ^ n17 ;
  assign n26 = n25 ^ x5 ;
  assign n27 = ~n16 & n26 ;
  assign n28 = n27 ^ n17 ;
  assign n29 = n28 ^ n20 ;
  assign n30 = n29 ^ n24 ;
  assign n31 = n30 ^ n9 ;
  assign n32 = n31 ^ n10 ;
  assign n33 = n32 ^ x4 ;
  assign n34 = n33 ^ x5 ;
  assign y0 = ~n34 ;
endmodule
