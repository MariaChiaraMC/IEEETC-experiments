module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 ;
  assign n18 = x15 ^ x14 ;
  assign n19 = n18 ^ x6 ;
  assign n20 = n19 ^ x5 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n21 ^ x15 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = x4 & n23 ;
  assign n25 = n24 ^ n18 ;
  assign n26 = x5 ^ x4 ;
  assign n27 = n26 ^ n18 ;
  assign n28 = ~n22 & ~n27 ;
  assign n29 = n28 ^ n21 ;
  assign n30 = n29 ^ n22 ;
  assign n31 = n25 & n30 ;
  assign n32 = ~n21 & n31 ;
  assign n33 = n32 ^ n24 ;
  assign n34 = n33 ^ x14 ;
  assign n35 = x12 & n34 ;
  assign n36 = ~x8 & x14 ;
  assign n37 = ~x1 & x2 ;
  assign n38 = n36 & n37 ;
  assign n39 = ~x9 & ~x10 ;
  assign n40 = x0 & ~n39 ;
  assign n41 = x5 & x6 ;
  assign n42 = ~x7 & n41 ;
  assign n43 = ~n40 & n42 ;
  assign n44 = n38 & n43 ;
  assign n45 = x4 & n44 ;
  assign n46 = ~n35 & ~n45 ;
  assign n47 = ~x13 & ~x16 ;
  assign n48 = ~n46 & n47 ;
  assign n49 = x11 ^ x2 ;
  assign n50 = n49 ^ x11 ;
  assign n51 = n50 ^ x13 ;
  assign n52 = ~x5 & x15 ;
  assign n53 = ~x4 & ~x14 ;
  assign n54 = x6 & n53 ;
  assign n55 = n52 & n54 ;
  assign n56 = ~x4 & n41 ;
  assign n57 = ~x5 & ~x6 ;
  assign n58 = ~x7 & n57 ;
  assign n59 = x4 & n58 ;
  assign n60 = ~n56 & ~n59 ;
  assign n61 = ~x15 & ~n60 ;
  assign n62 = x14 & n61 ;
  assign n63 = ~n55 & ~n62 ;
  assign n64 = ~x6 & x15 ;
  assign n65 = ~x7 & n53 ;
  assign n66 = n64 & n65 ;
  assign n67 = x5 & n66 ;
  assign n68 = x11 & ~n67 ;
  assign n69 = n63 & n68 ;
  assign n70 = ~x6 & ~x7 ;
  assign n71 = x5 & ~n70 ;
  assign n72 = ~n57 & ~n71 ;
  assign n73 = n53 & n72 ;
  assign n74 = ~x14 & ~x15 ;
  assign n75 = x5 & ~x6 ;
  assign n76 = ~x1 & ~n75 ;
  assign n77 = n74 & ~n76 ;
  assign n78 = ~n73 & ~n77 ;
  assign n79 = ~x11 & ~n61 ;
  assign n80 = n78 & n79 ;
  assign n81 = x3 & ~n80 ;
  assign n82 = ~n69 & n81 ;
  assign n83 = ~x3 & ~x11 ;
  assign n84 = n74 & n83 ;
  assign n85 = x1 & n84 ;
  assign n86 = n85 ^ n82 ;
  assign n87 = ~n82 & n86 ;
  assign n88 = n87 ^ x11 ;
  assign n89 = n88 ^ n82 ;
  assign n90 = n51 & ~n89 ;
  assign n91 = n90 ^ n87 ;
  assign n92 = n91 ^ n82 ;
  assign n93 = ~x13 & ~n92 ;
  assign n94 = n93 ^ x13 ;
  assign n95 = ~x11 & ~x13 ;
  assign n96 = x2 & ~n95 ;
  assign n97 = ~n74 & n96 ;
  assign n98 = n97 ^ x1 ;
  assign n99 = n98 ^ n97 ;
  assign n100 = x3 & n70 ;
  assign n101 = n74 & n95 ;
  assign n102 = ~x2 & n101 ;
  assign n103 = ~n100 & n102 ;
  assign n104 = x13 & n64 ;
  assign n105 = n18 ^ x15 ;
  assign n106 = ~x8 & x13 ;
  assign n107 = n106 ^ x15 ;
  assign n108 = n105 & ~n107 ;
  assign n109 = n108 ^ x15 ;
  assign n110 = ~n104 & ~n109 ;
  assign n111 = n96 & ~n110 ;
  assign n112 = ~n103 & ~n111 ;
  assign n113 = ~x5 & ~n112 ;
  assign n114 = x7 & n97 ;
  assign n115 = ~n102 & ~n114 ;
  assign n116 = n41 & ~n115 ;
  assign n117 = ~n113 & ~n116 ;
  assign n118 = x4 & ~n117 ;
  assign n119 = ~x2 & x3 ;
  assign n120 = ~x14 & n106 ;
  assign n121 = ~n119 & ~n120 ;
  assign n122 = ~n57 & ~n121 ;
  assign n123 = ~x8 & n41 ;
  assign n124 = x13 & n123 ;
  assign n125 = x2 & ~n124 ;
  assign n126 = ~n101 & ~n125 ;
  assign n127 = x4 ^ x2 ;
  assign n128 = ~n74 & ~n95 ;
  assign n129 = n128 ^ x4 ;
  assign n130 = n129 ^ n128 ;
  assign n131 = n128 ^ n75 ;
  assign n132 = n130 & ~n131 ;
  assign n133 = n132 ^ n128 ;
  assign n134 = n127 & n133 ;
  assign n135 = n134 ^ x2 ;
  assign n136 = ~n126 & ~n135 ;
  assign n137 = ~n122 & n136 ;
  assign n138 = ~n118 & ~n137 ;
  assign n139 = n138 ^ n97 ;
  assign n140 = ~n99 & ~n139 ;
  assign n141 = n140 ^ n97 ;
  assign n142 = n94 & ~n141 ;
  assign n143 = n40 & ~n142 ;
  assign n144 = ~x14 & x15 ;
  assign n145 = x3 & x5 ;
  assign n146 = ~x2 & n145 ;
  assign n147 = n144 & n146 ;
  assign n148 = x13 & n147 ;
  assign n149 = x1 & n148 ;
  assign n150 = x0 & n149 ;
  assign n151 = x2 & ~n74 ;
  assign n152 = ~x4 & n70 ;
  assign n153 = ~x13 & ~n152 ;
  assign n154 = n147 & ~n153 ;
  assign n155 = ~n151 & ~n154 ;
  assign n156 = x1 & ~n155 ;
  assign n157 = ~x2 & ~x13 ;
  assign n158 = ~n63 & n157 ;
  assign n159 = x3 & n158 ;
  assign n160 = ~n156 & ~n159 ;
  assign n161 = ~n40 & ~n160 ;
  assign n162 = x1 & x13 ;
  assign n163 = ~n145 & n162 ;
  assign n164 = ~x14 & n163 ;
  assign n165 = x4 & x14 ;
  assign n166 = x3 & ~x13 ;
  assign n167 = n165 & n166 ;
  assign n168 = n72 & n167 ;
  assign n169 = ~n164 & ~n168 ;
  assign n170 = ~x2 & x15 ;
  assign n171 = ~n169 & n170 ;
  assign n172 = ~n161 & ~n171 ;
  assign n173 = x6 & x13 ;
  assign n174 = n165 & n173 ;
  assign n178 = x13 ^ x5 ;
  assign n179 = n178 ^ x14 ;
  assign n183 = n179 ^ n178 ;
  assign n175 = x4 & ~x15 ;
  assign n176 = n175 ^ x13 ;
  assign n177 = n176 ^ n175 ;
  assign n180 = n179 ^ n175 ;
  assign n181 = n180 ^ n178 ;
  assign n182 = n177 & ~n181 ;
  assign n184 = n183 ^ n182 ;
  assign n185 = ~x4 & x6 ;
  assign n186 = n185 ^ n179 ;
  assign n187 = n183 & n186 ;
  assign n188 = n187 ^ n185 ;
  assign n189 = n184 & n188 ;
  assign n190 = n189 ^ n182 ;
  assign n191 = n190 ^ n179 ;
  assign n192 = n191 ^ x13 ;
  assign n193 = n192 ^ n178 ;
  assign n194 = ~n174 & ~n193 ;
  assign n195 = ~x8 & ~n194 ;
  assign n196 = n151 & ~n195 ;
  assign n197 = n56 ^ x5 ;
  assign n198 = n196 & ~n197 ;
  assign n199 = n65 & n166 ;
  assign n200 = ~x2 & ~n199 ;
  assign n201 = ~x13 & n36 ;
  assign n202 = x5 & n201 ;
  assign n203 = ~n74 & n197 ;
  assign n204 = ~n202 & ~n203 ;
  assign n205 = ~n200 & ~n204 ;
  assign n206 = x6 & x7 ;
  assign n207 = n165 & ~n206 ;
  assign n208 = n207 ^ x13 ;
  assign n209 = n208 ^ x8 ;
  assign n210 = n53 ^ x6 ;
  assign n211 = n210 ^ n208 ;
  assign n212 = ~n207 & ~n211 ;
  assign n213 = n212 ^ x6 ;
  assign n214 = n213 ^ n207 ;
  assign n215 = n214 ^ n208 ;
  assign n216 = n215 ^ x8 ;
  assign n217 = ~n209 & ~n216 ;
  assign n218 = n217 ^ n212 ;
  assign n219 = n218 ^ x6 ;
  assign n220 = n219 ^ n208 ;
  assign n221 = ~x8 & ~n220 ;
  assign n222 = n221 ^ x8 ;
  assign n223 = n222 ^ x8 ;
  assign n224 = n205 & ~n223 ;
  assign n225 = ~n198 & ~n224 ;
  assign n226 = ~n40 & ~n225 ;
  assign n227 = ~x5 & n64 ;
  assign n228 = x8 & ~n74 ;
  assign n229 = n228 ^ n41 ;
  assign n230 = n228 ^ x6 ;
  assign n231 = n228 ^ x14 ;
  assign n232 = n228 & n231 ;
  assign n233 = n232 ^ n228 ;
  assign n234 = n230 & n233 ;
  assign n235 = n234 ^ n232 ;
  assign n236 = n235 ^ n228 ;
  assign n237 = n236 ^ x14 ;
  assign n238 = ~n229 & n237 ;
  assign n239 = n238 ^ n228 ;
  assign n240 = ~n227 & ~n239 ;
  assign n241 = ~x2 & ~n240 ;
  assign n242 = x15 & n123 ;
  assign n243 = ~x4 & ~n242 ;
  assign n244 = ~n65 & ~n243 ;
  assign n245 = ~n241 & ~n244 ;
  assign n246 = x5 & ~n206 ;
  assign n247 = ~x5 & n36 ;
  assign n248 = n247 ^ x14 ;
  assign n249 = ~n227 & ~n248 ;
  assign n250 = ~n246 & ~n249 ;
  assign n251 = ~n144 & ~n250 ;
  assign n252 = ~x2 & ~n251 ;
  assign n253 = ~x5 & ~x15 ;
  assign n254 = n36 & n253 ;
  assign n255 = n206 & n254 ;
  assign n256 = x4 & ~n255 ;
  assign n257 = ~n252 & n256 ;
  assign n258 = x13 & ~n257 ;
  assign n259 = ~n245 & n258 ;
  assign n260 = ~n226 & ~n259 ;
  assign n261 = n260 ^ x1 ;
  assign n262 = n261 ^ n260 ;
  assign n263 = n262 ^ n172 ;
  assign n264 = x13 & x14 ;
  assign n265 = n264 ^ x2 ;
  assign n266 = n264 & ~n265 ;
  assign n267 = n266 ^ n260 ;
  assign n268 = n267 ^ n264 ;
  assign n269 = n263 & ~n268 ;
  assign n270 = n269 ^ n266 ;
  assign n271 = n270 ^ n264 ;
  assign n272 = n172 & n271 ;
  assign n273 = n272 ^ n172 ;
  assign n274 = ~n150 & n273 ;
  assign n275 = ~n143 & n274 ;
  assign n276 = ~x16 & ~n275 ;
  assign n277 = x16 & n53 ;
  assign n278 = n253 & n277 ;
  assign n279 = ~x1 & ~n206 ;
  assign n280 = n106 & n279 ;
  assign n281 = n278 & n280 ;
  assign n282 = x2 & n40 ;
  assign n283 = ~n264 & ~n282 ;
  assign n284 = x8 & ~n40 ;
  assign n285 = x2 & n284 ;
  assign n286 = ~x16 & ~n285 ;
  assign n287 = x15 & n106 ;
  assign n288 = x14 & n287 ;
  assign n289 = x4 & n128 ;
  assign n290 = ~n288 & n289 ;
  assign n291 = ~x1 & n246 ;
  assign n292 = n290 & n291 ;
  assign n293 = n286 & n292 ;
  assign n294 = ~n283 & n293 ;
  assign n295 = ~n281 & ~n294 ;
  assign n296 = ~n276 & n295 ;
  assign n297 = ~x12 & ~n296 ;
  assign n306 = ~x6 & ~x13 ;
  assign n307 = x12 & n306 ;
  assign n298 = ~x4 & x14 ;
  assign n299 = x14 & ~x15 ;
  assign n300 = ~x5 & ~n299 ;
  assign n301 = ~n298 & ~n300 ;
  assign n302 = x4 & ~x14 ;
  assign n303 = x5 & ~x15 ;
  assign n304 = ~n302 & ~n303 ;
  assign n305 = n301 & n304 ;
  assign n308 = n307 ^ n305 ;
  assign n309 = n305 ^ n278 ;
  assign n310 = n309 ^ n278 ;
  assign n311 = ~x16 & n70 ;
  assign n312 = n280 & ~n311 ;
  assign n313 = ~x12 & n312 ;
  assign n314 = n313 ^ n278 ;
  assign n315 = n310 & ~n314 ;
  assign n316 = n315 ^ n278 ;
  assign n317 = n308 & ~n316 ;
  assign n318 = n317 ^ n307 ;
  assign n319 = ~n297 & ~n318 ;
  assign n320 = ~n48 & n319 ;
  assign y0 = ~n320 ;
endmodule
