module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 ;
  assign n15 = x12 ^ x10 ;
  assign n16 = x12 ^ x6 ;
  assign n17 = x12 ^ x11 ;
  assign n18 = ~x12 & ~n17 ;
  assign n19 = n18 ^ x12 ;
  assign n20 = ~n16 & ~n19 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n21 ^ x12 ;
  assign n23 = n22 ^ x11 ;
  assign n24 = n15 & ~n23 ;
  assign n25 = n24 ^ x10 ;
  assign n26 = ~x5 & ~n25 ;
  assign n27 = ~x6 & x13 ;
  assign n28 = x13 ^ x4 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = x3 & ~x11 ;
  assign n31 = ~x10 & ~n30 ;
  assign n32 = ~x8 & ~x12 ;
  assign n33 = ~n31 & n32 ;
  assign n34 = n33 ^ x0 ;
  assign n35 = ~x4 & n34 ;
  assign n36 = n35 ^ x0 ;
  assign n37 = n29 & ~n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = n38 ^ x0 ;
  assign n40 = n39 ^ x4 ;
  assign n41 = ~n27 & n40 ;
  assign n42 = n41 ^ x9 ;
  assign n43 = n42 ^ n41 ;
  assign n45 = ~x6 & ~n28 ;
  assign n46 = n45 ^ x4 ;
  assign n44 = x13 ^ x11 ;
  assign n47 = n46 ^ n44 ;
  assign n48 = n47 ^ x12 ;
  assign n49 = n48 ^ n44 ;
  assign n50 = n49 ^ n17 ;
  assign n51 = n44 ^ x10 ;
  assign n52 = ~n50 & n51 ;
  assign n53 = n52 ^ n44 ;
  assign n54 = n53 ^ n48 ;
  assign n55 = n54 ^ x10 ;
  assign n56 = n17 ^ x11 ;
  assign n57 = x10 & n56 ;
  assign n58 = n57 ^ n44 ;
  assign n59 = n58 ^ n48 ;
  assign n60 = n59 ^ x11 ;
  assign n61 = n60 ^ x10 ;
  assign n62 = n44 ^ x0 ;
  assign n63 = n62 ^ n17 ;
  assign n64 = n63 ^ x10 ;
  assign n65 = ~n62 & ~n64 ;
  assign n66 = n65 ^ n48 ;
  assign n67 = n66 ^ x10 ;
  assign n68 = ~n61 & ~n67 ;
  assign n69 = n68 ^ n48 ;
  assign n70 = ~n55 & ~n69 ;
  assign n71 = n70 ^ n57 ;
  assign n72 = n71 ^ n52 ;
  assign n73 = n72 ^ n44 ;
  assign n74 = n73 ^ n48 ;
  assign n75 = n74 ^ x11 ;
  assign n76 = n75 ^ n17 ;
  assign n77 = n76 ^ x10 ;
  assign n78 = n77 ^ n41 ;
  assign n79 = n43 & ~n78 ;
  assign n80 = n79 ^ n41 ;
  assign n81 = n26 & n80 ;
  assign y0 = n81 ;
endmodule
