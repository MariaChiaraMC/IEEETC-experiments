module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 ;
  assign n13 = x6 & ~x8 ;
  assign n14 = x3 & x5 ;
  assign n15 = n13 & n14 ;
  assign n10 = ~x6 & ~x7 ;
  assign n11 = x5 & n10 ;
  assign n12 = ~x8 & n11 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = n16 ^ x1 ;
  assign n24 = n17 ^ n16 ;
  assign n18 = n17 ^ x6 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n17 ^ n12 ;
  assign n21 = n20 ^ x6 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n19 & n22 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ n19 ;
  assign n27 = ~x5 & ~x7 ;
  assign n28 = n27 ^ n16 ;
  assign n29 = n23 ^ n19 ;
  assign n30 = n28 & n29 ;
  assign n31 = n30 ^ n16 ;
  assign n32 = ~n26 & n31 ;
  assign n33 = n32 ^ n16 ;
  assign n34 = n33 ^ n15 ;
  assign n35 = n34 ^ n16 ;
  assign n36 = ~x4 & n35 ;
  assign n37 = ~x4 & ~x5 ;
  assign n38 = x8 & n37 ;
  assign n39 = x6 & x7 ;
  assign n40 = n39 ^ x7 ;
  assign n41 = ~x3 & ~n40 ;
  assign n42 = n41 ^ x7 ;
  assign n43 = n38 & ~n42 ;
  assign n44 = x4 & ~x8 ;
  assign n45 = x5 & n44 ;
  assign n47 = x6 & ~x7 ;
  assign n46 = ~x6 & x7 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = n47 ^ x1 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = n49 & ~n51 ;
  assign n53 = n52 ^ n47 ;
  assign n54 = x3 & n53 ;
  assign n55 = n54 ^ n47 ;
  assign n56 = n45 & n55 ;
  assign n57 = ~n43 & ~n56 ;
  assign n58 = ~x3 & ~x6 ;
  assign n59 = ~x7 & ~x8 ;
  assign n60 = x7 & x8 ;
  assign n61 = x5 & n60 ;
  assign n62 = ~n59 & ~n61 ;
  assign n63 = n58 & ~n62 ;
  assign n64 = ~x5 & x6 ;
  assign n65 = x7 & ~x8 ;
  assign n66 = n64 & n65 ;
  assign n69 = n66 ^ n47 ;
  assign n70 = n69 ^ n66 ;
  assign n67 = n66 ^ x5 ;
  assign n68 = n67 ^ n66 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = n66 ^ x1 ;
  assign n73 = n72 ^ n66 ;
  assign n74 = n73 ^ n70 ;
  assign n75 = n70 & n74 ;
  assign n76 = n75 ^ n70 ;
  assign n77 = n71 & n76 ;
  assign n78 = n77 ^ n75 ;
  assign n79 = n78 ^ n66 ;
  assign n80 = n79 ^ n70 ;
  assign n81 = ~x3 & n80 ;
  assign n82 = n81 ^ n66 ;
  assign n83 = ~n63 & ~n82 ;
  assign n84 = ~x4 & ~n83 ;
  assign n85 = x7 ^ x6 ;
  assign n86 = x4 & ~x5 ;
  assign n87 = ~x6 & n86 ;
  assign n88 = n87 ^ n85 ;
  assign n89 = x8 ^ x6 ;
  assign n90 = n89 ^ x8 ;
  assign n91 = x4 & x5 ;
  assign n92 = n91 ^ x8 ;
  assign n93 = n90 & n92 ;
  assign n94 = n93 ^ x8 ;
  assign n95 = n94 ^ n85 ;
  assign n96 = n88 & ~n95 ;
  assign n97 = n96 ^ n93 ;
  assign n98 = n97 ^ x8 ;
  assign n99 = n98 ^ n87 ;
  assign n100 = ~n85 & ~n99 ;
  assign n101 = n100 ^ n85 ;
  assign n102 = n101 ^ n87 ;
  assign n103 = x3 & ~n102 ;
  assign n104 = ~n13 & ~n58 ;
  assign n105 = n27 & ~n104 ;
  assign n106 = x5 & n47 ;
  assign n107 = ~x4 & x8 ;
  assign n108 = n106 & n107 ;
  assign n109 = ~n105 & ~n108 ;
  assign n110 = x7 & ~n107 ;
  assign n111 = ~x3 & x5 ;
  assign n112 = ~x6 & ~x8 ;
  assign n113 = ~n111 & ~n112 ;
  assign n114 = ~n44 & ~n113 ;
  assign n115 = n110 & n114 ;
  assign n116 = ~x1 & ~n115 ;
  assign n117 = n109 & n116 ;
  assign n118 = ~n103 & n117 ;
  assign n119 = x4 & ~x6 ;
  assign n120 = ~n65 & ~n119 ;
  assign n121 = n14 & ~n120 ;
  assign n122 = n121 ^ x1 ;
  assign n123 = ~x7 & n64 ;
  assign n124 = ~n37 & ~n123 ;
  assign n125 = ~x3 & n39 ;
  assign n126 = ~x4 & n39 ;
  assign n127 = ~n125 & ~n126 ;
  assign n128 = n124 & n127 ;
  assign n129 = n128 ^ x8 ;
  assign n130 = n129 ^ n128 ;
  assign n131 = n128 ^ n87 ;
  assign n132 = ~n130 & ~n131 ;
  assign n133 = n132 ^ n128 ;
  assign n134 = n133 ^ n121 ;
  assign n135 = ~n122 & ~n134 ;
  assign n136 = n135 ^ n132 ;
  assign n137 = n136 ^ n128 ;
  assign n138 = n137 ^ x1 ;
  assign n139 = ~n121 & n138 ;
  assign n140 = n139 ^ n121 ;
  assign n141 = ~n118 & n140 ;
  assign n142 = ~n84 & ~n141 ;
  assign n143 = n142 ^ x2 ;
  assign n144 = n143 ^ n142 ;
  assign n145 = n45 & n58 ;
  assign n146 = n60 & n119 ;
  assign n147 = ~x3 & n126 ;
  assign n148 = ~n146 & ~n147 ;
  assign n149 = x6 & n91 ;
  assign n150 = n149 ^ x8 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = n151 ^ x3 ;
  assign n153 = ~n47 & ~n119 ;
  assign n154 = n153 ^ n86 ;
  assign n155 = ~n86 & n154 ;
  assign n156 = n155 ^ n149 ;
  assign n157 = n156 ^ n86 ;
  assign n158 = ~n152 & n157 ;
  assign n159 = n158 ^ n155 ;
  assign n160 = n159 ^ n86 ;
  assign n161 = x3 & ~n160 ;
  assign n162 = n161 ^ x3 ;
  assign n163 = n148 & ~n162 ;
  assign n164 = ~n145 & n163 ;
  assign n165 = x1 & ~n164 ;
  assign n166 = x8 ^ x3 ;
  assign n167 = ~x4 & ~n166 ;
  assign n168 = n167 ^ x3 ;
  assign n169 = n64 & ~n168 ;
  assign n170 = ~n110 & n169 ;
  assign n171 = ~x3 & ~n91 ;
  assign n172 = x7 & ~n37 ;
  assign n173 = n112 & ~n172 ;
  assign n174 = ~n171 & n173 ;
  assign n175 = ~n170 & ~n174 ;
  assign n176 = ~n165 & n175 ;
  assign n177 = n176 ^ n142 ;
  assign n178 = ~n144 & n177 ;
  assign n179 = n178 ^ n142 ;
  assign n180 = n57 & n179 ;
  assign n181 = ~n36 & n180 ;
  assign n182 = ~x0 & ~n181 ;
  assign n183 = x5 ^ x4 ;
  assign n184 = x4 ^ x3 ;
  assign n185 = ~n183 & ~n184 ;
  assign n186 = n185 ^ x3 ;
  assign n187 = ~x0 & n186 ;
  assign n188 = x3 & ~n172 ;
  assign n189 = x8 & ~n188 ;
  assign n190 = n187 & n189 ;
  assign n191 = x8 ^ x0 ;
  assign n201 = n191 ^ x8 ;
  assign n202 = n201 ^ x3 ;
  assign n192 = x8 ^ x7 ;
  assign n193 = n192 ^ n191 ;
  assign n194 = n193 ^ n191 ;
  assign n195 = n194 ^ x8 ;
  assign n196 = n195 ^ x3 ;
  assign n197 = n193 ^ x4 ;
  assign n198 = n197 ^ n193 ;
  assign n199 = n198 ^ n196 ;
  assign n200 = n196 & ~n199 ;
  assign n203 = n202 ^ n200 ;
  assign n204 = n203 ^ n196 ;
  assign n205 = n202 ^ x3 ;
  assign n206 = n205 ^ n202 ;
  assign n207 = x8 ^ x5 ;
  assign n210 = n207 ^ x8 ;
  assign n211 = n210 ^ n207 ;
  assign n212 = n211 ^ n202 ;
  assign n213 = n212 ^ n205 ;
  assign n214 = n212 & ~n213 ;
  assign n208 = n207 ^ n198 ;
  assign n209 = ~n205 & ~n208 ;
  assign n215 = n214 ^ n209 ;
  assign n216 = n215 ^ n207 ;
  assign n217 = n206 & n216 ;
  assign n218 = n217 ^ n209 ;
  assign n219 = n218 ^ n210 ;
  assign n220 = n219 ^ n202 ;
  assign n221 = ~n204 & n220 ;
  assign n222 = n221 ^ n209 ;
  assign n223 = n222 ^ n214 ;
  assign n224 = n223 ^ n217 ;
  assign n225 = n224 ^ n207 ;
  assign n226 = n225 ^ n202 ;
  assign n227 = n226 ^ n205 ;
  assign n228 = x6 & ~n227 ;
  assign n229 = ~n46 & ~n106 ;
  assign n230 = n107 & n229 ;
  assign n231 = ~x4 & n10 ;
  assign n232 = ~n45 & ~n231 ;
  assign n233 = x0 & ~n232 ;
  assign n234 = x4 & n47 ;
  assign n235 = x0 & n87 ;
  assign n236 = ~n234 & ~n235 ;
  assign n237 = n236 ^ x8 ;
  assign n238 = n237 ^ n236 ;
  assign n239 = n238 ^ n233 ;
  assign n240 = x7 & n37 ;
  assign n241 = n240 ^ x6 ;
  assign n242 = n240 & ~n241 ;
  assign n243 = n242 ^ n236 ;
  assign n244 = n243 ^ n240 ;
  assign n245 = n239 & ~n244 ;
  assign n246 = n245 ^ n242 ;
  assign n247 = n246 ^ n240 ;
  assign n248 = ~n233 & n247 ;
  assign n249 = n248 ^ n233 ;
  assign n250 = ~n230 & ~n249 ;
  assign n251 = ~x3 & ~n250 ;
  assign n252 = ~n228 & ~n251 ;
  assign n253 = ~n190 & n252 ;
  assign n254 = ~x2 & ~n253 ;
  assign n255 = ~x1 & n254 ;
  assign n256 = ~n182 & ~n255 ;
  assign y0 = ~n256 ;
endmodule
