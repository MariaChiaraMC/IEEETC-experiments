module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 ;
  assign n9 = ~x3 & x4 ;
  assign n10 = x6 & x7 ;
  assign n11 = n9 & n10 ;
  assign n12 = x5 ^ x0 ;
  assign n13 = n11 & n12 ;
  assign n16 = x5 ^ x3 ;
  assign n17 = n16 ^ x6 ;
  assign n20 = n17 ^ x4 ;
  assign n21 = n20 ^ x5 ;
  assign n22 = n21 ^ x6 ;
  assign n29 = n22 ^ x5 ;
  assign n30 = n29 ^ x7 ;
  assign n14 = x3 ^ x0 ;
  assign n31 = n30 ^ n14 ;
  assign n15 = n14 ^ x6 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n18 ^ x7 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n17 ^ n14 ;
  assign n26 = n24 ^ n14 ;
  assign n25 = n24 ^ n23 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = n23 & ~n27 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = n32 ^ n24 ;
  assign n34 = n31 ^ n22 ;
  assign n35 = n34 ^ n17 ;
  assign n43 = n35 ^ n23 ;
  assign n44 = n31 ^ n23 ;
  assign n45 = n44 ^ n26 ;
  assign n46 = ~n43 & ~n45 ;
  assign n36 = n14 ^ x7 ;
  assign n37 = n36 ^ n19 ;
  assign n38 = n37 ^ n19 ;
  assign n39 = n38 ^ n30 ;
  assign n40 = n39 ^ n31 ;
  assign n41 = n40 ^ n26 ;
  assign n42 = ~n35 & n41 ;
  assign n47 = n46 ^ n42 ;
  assign n48 = n47 ^ n39 ;
  assign n49 = n48 ^ n23 ;
  assign n50 = n49 ^ n24 ;
  assign n51 = n26 & n50 ;
  assign n52 = n51 ^ n42 ;
  assign n53 = n52 ^ n31 ;
  assign n54 = n53 ^ n39 ;
  assign n55 = n54 ^ n23 ;
  assign n56 = n55 ^ n24 ;
  assign n57 = n56 ^ n26 ;
  assign n58 = n57 ^ n35 ;
  assign n59 = n33 & n58 ;
  assign n60 = n59 ^ n42 ;
  assign n61 = n60 ^ n46 ;
  assign n62 = n61 ^ n28 ;
  assign n63 = n62 ^ n51 ;
  assign n64 = n63 ^ n31 ;
  assign n65 = n64 ^ n39 ;
  assign n66 = n65 ^ n23 ;
  assign n67 = n66 ^ x1 ;
  assign n68 = n67 ^ n66 ;
  assign n69 = x5 & ~x6 ;
  assign n70 = x7 & n69 ;
  assign n71 = x6 & ~x7 ;
  assign n72 = ~n70 & ~n71 ;
  assign n73 = ~x0 & x5 ;
  assign n74 = n9 & ~n73 ;
  assign n75 = ~n72 & n74 ;
  assign n82 = x3 & x5 ;
  assign n83 = n10 & n82 ;
  assign n76 = n10 ^ x3 ;
  assign n77 = ~x5 & ~x7 ;
  assign n78 = ~n10 & n77 ;
  assign n79 = n76 & n78 ;
  assign n80 = n79 ^ n76 ;
  assign n81 = ~n69 & n80 ;
  assign n84 = n83 ^ n81 ;
  assign n85 = n84 ^ n81 ;
  assign n86 = ~x3 & ~x5 ;
  assign n87 = ~x6 & n86 ;
  assign n88 = n87 ^ n81 ;
  assign n89 = n88 ^ n81 ;
  assign n90 = ~n85 & ~n89 ;
  assign n91 = n90 ^ n81 ;
  assign n92 = ~x0 & ~n91 ;
  assign n93 = n92 ^ n81 ;
  assign n94 = ~x4 & n93 ;
  assign n95 = ~n75 & ~n94 ;
  assign n96 = n95 ^ n66 ;
  assign n97 = n68 & ~n96 ;
  assign n98 = n97 ^ n66 ;
  assign n99 = ~n13 & ~n98 ;
  assign n100 = ~x2 & ~n99 ;
  assign n101 = ~x0 & ~x5 ;
  assign n102 = ~x1 & ~x3 ;
  assign n103 = x2 & x7 ;
  assign n104 = ~n102 & n103 ;
  assign n105 = n101 & n104 ;
  assign n106 = x1 & x3 ;
  assign n107 = x4 & x6 ;
  assign n108 = n107 ^ x4 ;
  assign n109 = ~n106 & ~n108 ;
  assign n110 = n109 ^ x4 ;
  assign n111 = n105 & ~n110 ;
  assign n112 = x2 & x3 ;
  assign n113 = n71 & n112 ;
  assign n114 = ~x4 & ~x5 ;
  assign n115 = n113 & n114 ;
  assign n116 = x1 & n115 ;
  assign n117 = ~n111 & ~n116 ;
  assign n118 = x4 & x7 ;
  assign n119 = x2 & ~x3 ;
  assign n120 = ~n118 & ~n119 ;
  assign n121 = x1 & ~n9 ;
  assign n122 = ~x6 & n121 ;
  assign n123 = ~n120 & n122 ;
  assign n124 = x7 ^ x3 ;
  assign n131 = x2 ^ x1 ;
  assign n125 = x7 ^ x2 ;
  assign n126 = n125 ^ x1 ;
  assign n127 = n126 ^ x2 ;
  assign n137 = n127 ^ x2 ;
  assign n128 = n127 ^ x6 ;
  assign n138 = n137 ^ n128 ;
  assign n139 = n131 & ~n138 ;
  assign n129 = x6 ^ x4 ;
  assign n130 = n129 ^ x6 ;
  assign n132 = n131 ^ n130 ;
  assign n133 = ~n128 & n132 ;
  assign n145 = n139 ^ n133 ;
  assign n134 = n133 ^ n127 ;
  assign n135 = n134 ^ n131 ;
  assign n136 = n135 ^ n128 ;
  assign n140 = n139 ^ n127 ;
  assign n141 = n140 ^ n131 ;
  assign n142 = n141 ^ n128 ;
  assign n143 = n142 ^ n124 ;
  assign n144 = n136 & n143 ;
  assign n146 = n145 ^ n144 ;
  assign n147 = n124 & n146 ;
  assign n148 = ~n123 & ~n147 ;
  assign n149 = n73 & ~n148 ;
  assign n150 = ~x4 & n69 ;
  assign n151 = ~n107 & ~n150 ;
  assign n152 = n121 & ~n151 ;
  assign n153 = ~x5 & ~x6 ;
  assign n154 = ~x1 & ~x4 ;
  assign n155 = ~n153 & n154 ;
  assign n156 = n16 & n155 ;
  assign n157 = ~n152 & ~n156 ;
  assign n158 = x2 & ~n157 ;
  assign n159 = ~x5 & n107 ;
  assign n160 = n102 & n159 ;
  assign n161 = ~n158 & ~n160 ;
  assign n162 = x0 & x7 ;
  assign n163 = ~n161 & n162 ;
  assign n164 = ~n149 & ~n163 ;
  assign n165 = n117 & n164 ;
  assign n166 = ~n100 & n165 ;
  assign y0 = ~n166 ;
endmodule
