module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 ;
  assign n11 = x7 ^ x6 ;
  assign n19 = n11 ^ x9 ;
  assign n20 = n19 ^ x6 ;
  assign n17 = n11 ^ x8 ;
  assign n18 = n17 ^ x3 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n21 ^ x3 ;
  assign n23 = n18 ^ n11 ;
  assign n24 = n23 ^ x3 ;
  assign n25 = n24 ^ x6 ;
  assign n26 = ~n22 & ~n25 ;
  assign n13 = x4 & x5 ;
  assign n14 = ~x2 & ~n13 ;
  assign n12 = x6 ^ x3 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = ~n11 & n15 ;
  assign n27 = n26 ^ n16 ;
  assign n28 = n27 ^ n20 ;
  assign n29 = n28 ^ x3 ;
  assign n30 = n29 ^ x6 ;
  assign n31 = n30 ^ n14 ;
  assign n32 = n21 ^ x6 ;
  assign n33 = n24 ^ n14 ;
  assign n34 = ~n32 & n33 ;
  assign n35 = n34 ^ n26 ;
  assign n36 = n35 ^ x3 ;
  assign n37 = n36 ^ n14 ;
  assign n38 = n14 & ~n37 ;
  assign n39 = n38 ^ n14 ;
  assign n40 = n31 & n39 ;
  assign n41 = ~x6 & ~x7 ;
  assign n42 = ~x4 & ~x5 ;
  assign n43 = n42 ^ x8 ;
  assign n44 = n43 ^ x8 ;
  assign n45 = x8 ^ x3 ;
  assign n46 = n44 & ~n45 ;
  assign n47 = n46 ^ x8 ;
  assign n48 = n41 & n47 ;
  assign n49 = n48 ^ n42 ;
  assign n50 = n40 & n49 ;
  assign n51 = ~x3 & x9 ;
  assign n52 = n41 & n42 ;
  assign n53 = n51 & n52 ;
  assign n54 = x2 & n53 ;
  assign n55 = ~n50 & ~n54 ;
  assign n56 = ~x0 & ~x1 ;
  assign n57 = ~n55 & n56 ;
  assign y0 = n57 ;
endmodule
