module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
  assign n9 = ~x0 & ~x1 ;
  assign n10 = ~x3 & n9 ;
  assign n11 = ~x4 & ~x7 ;
  assign n12 = n11 ^ x5 ;
  assign n13 = n11 ^ x2 ;
  assign n14 = n13 ^ n11 ;
  assign n15 = ~n12 & ~n14 ;
  assign n16 = n15 ^ n11 ;
  assign n17 = ~x6 & ~n11 ;
  assign n18 = n17 ^ n10 ;
  assign n19 = ~n16 & n18 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n10 & n20 ;
  assign n22 = n21 ^ n10 ;
  assign n23 = n22 ^ n10 ;
  assign n24 = x7 ^ x5 ;
  assign n25 = n24 ^ x7 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = x6 ^ x2 ;
  assign n28 = x7 & ~n27 ;
  assign n29 = n28 ^ x6 ;
  assign n30 = n26 & ~n29 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n31 ^ x6 ;
  assign n33 = n32 ^ x7 ;
  assign n34 = x4 & ~n33 ;
  assign n35 = n23 & ~n34 ;
  assign y0 = n35 ;
endmodule
