module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 ;
  assign n8 = x3 & ~x4 ;
  assign n9 = n8 ^ x0 ;
  assign n10 = n9 ^ x1 ;
  assign n11 = n9 ^ n8 ;
  assign n12 = ~x3 & x4 ;
  assign n13 = n12 ^ n8 ;
  assign n14 = n8 & n13 ;
  assign n15 = n14 ^ n8 ;
  assign n16 = ~n11 & n15 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = n17 ^ n8 ;
  assign n19 = n18 ^ n12 ;
  assign n20 = n10 & n19 ;
  assign n21 = n20 ^ n9 ;
  assign n22 = x2 & n21 ;
  assign n7 = x0 & x3 ;
  assign n23 = n22 ^ n7 ;
  assign n24 = n23 ^ x5 ;
  assign n31 = n24 ^ n23 ;
  assign n25 = n24 ^ x2 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n7 ^ x2 ;
  assign n28 = n27 ^ x2 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = n26 & n29 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = n32 ^ n26 ;
  assign n34 = n23 ^ x1 ;
  assign n35 = n30 ^ n26 ;
  assign n36 = ~n34 & n35 ;
  assign n37 = n36 ^ n23 ;
  assign n38 = n33 & ~n37 ;
  assign n39 = n38 ^ n23 ;
  assign n40 = n39 ^ n7 ;
  assign n41 = n40 ^ n23 ;
  assign n57 = ~x2 & x4 ;
  assign n58 = ~x4 & ~x5 ;
  assign n59 = ~n57 & ~n58 ;
  assign n60 = ~x2 & n8 ;
  assign n61 = ~n59 & ~n60 ;
  assign n45 = x5 ^ x3 ;
  assign n42 = x2 ^ x0 ;
  assign n43 = n42 ^ x5 ;
  assign n44 = n43 ^ x5 ;
  assign n46 = n45 ^ n44 ;
  assign n47 = n46 ^ x4 ;
  assign n48 = ~x4 & ~n47 ;
  assign n49 = n48 ^ n43 ;
  assign n50 = n49 ^ x4 ;
  assign n51 = n43 ^ x2 ;
  assign n52 = n45 & ~n51 ;
  assign n53 = n52 ^ n43 ;
  assign n54 = ~n50 & n53 ;
  assign n55 = n54 ^ n43 ;
  assign n56 = n55 ^ n45 ;
  assign n62 = n61 ^ n56 ;
  assign n63 = ~x1 & ~n62 ;
  assign n64 = n63 ^ n56 ;
  assign n65 = ~n41 & n64 ;
  assign y0 = ~n65 ;
endmodule
