module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 ;
  assign n17 = ~x0 & ~x3 ;
  assign n18 = ~x1 & n17 ;
  assign n19 = x11 & n18 ;
  assign n20 = ~x2 & n19 ;
  assign n21 = x6 ^ x5 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = ~x8 & ~x9 ;
  assign n24 = ~x10 & n23 ;
  assign n25 = x7 & ~n24 ;
  assign n26 = n25 ^ x6 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = x9 ^ x8 ;
  assign n29 = x7 & ~n28 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = ~n27 & n30 ;
  assign n32 = n31 ^ n25 ;
  assign n33 = n32 ^ n21 ;
  assign n34 = ~n22 & ~n33 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = n35 ^ n25 ;
  assign n37 = n36 ^ x4 ;
  assign n38 = n21 & n37 ;
  assign n39 = n38 ^ n21 ;
  assign n40 = n39 ^ x4 ;
  assign n41 = n20 & n40 ;
  assign n42 = ~x5 & x6 ;
  assign n43 = x6 & ~x10 ;
  assign n45 = x12 & x13 ;
  assign n44 = x14 & x15 ;
  assign n46 = n45 ^ n44 ;
  assign n47 = x8 & x9 ;
  assign n48 = ~n23 & ~n47 ;
  assign n49 = n48 ^ n45 ;
  assign n50 = n46 & n49 ;
  assign n51 = n50 ^ n45 ;
  assign n52 = n43 & n51 ;
  assign n53 = x5 & ~n52 ;
  assign n54 = ~x7 & n53 ;
  assign n55 = ~n42 & ~n54 ;
  assign n56 = n28 ^ x13 ;
  assign n57 = ~x6 & x14 ;
  assign n58 = ~x15 & n57 ;
  assign n59 = n58 ^ x12 ;
  assign n60 = n59 ^ n58 ;
  assign n61 = x7 & n44 ;
  assign n62 = n61 ^ n58 ;
  assign n63 = n60 & n62 ;
  assign n64 = n63 ^ n58 ;
  assign n65 = n64 ^ n28 ;
  assign n66 = ~n56 & n65 ;
  assign n67 = n66 ^ n63 ;
  assign n68 = n67 ^ n58 ;
  assign n69 = n68 ^ x13 ;
  assign n70 = n28 & ~n69 ;
  assign n71 = n70 ^ n28 ;
  assign n72 = x4 & ~n71 ;
  assign n73 = ~n55 & n72 ;
  assign n74 = n41 & ~n73 ;
  assign y0 = n74 ;
endmodule
