module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;
  assign n18 = ~x13 & ~x14 ;
  assign n17 = ~x8 & ~x15 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = x13 & x14 ;
  assign n21 = ~x11 & ~x12 ;
  assign n22 = ~n20 & n21 ;
  assign n23 = x8 & x15 ;
  assign n24 = x9 ^ x8 ;
  assign n25 = x10 ^ x8 ;
  assign n26 = ~n24 & ~n25 ;
  assign n27 = n26 ^ n22 ;
  assign n28 = n23 & n27 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = n22 & n29 ;
  assign n31 = n30 ^ n22 ;
  assign n32 = n19 & n31 ;
  assign n33 = ~x7 & ~n32 ;
  assign n34 = ~x0 & x1 ;
  assign n35 = ~x5 & x6 ;
  assign n36 = n34 & n35 ;
  assign n37 = ~x2 & n36 ;
  assign n38 = ~n33 & n37 ;
  assign n39 = ~x1 & x5 ;
  assign n40 = x0 & n39 ;
  assign n41 = ~n38 & ~n40 ;
  assign n42 = ~x3 & ~n41 ;
  assign n43 = ~x4 & n42 ;
  assign y0 = n43 ;
endmodule
