module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 ;
  assign n11 = x8 & x9 ;
  assign n12 = ~x3 & ~n11 ;
  assign n13 = ~x8 & ~x9 ;
  assign n14 = x7 & n13 ;
  assign n15 = n12 & ~n14 ;
  assign n16 = x2 & ~x6 ;
  assign n17 = ~x5 & n16 ;
  assign n18 = ~n15 & n17 ;
  assign n19 = x3 & x5 ;
  assign n20 = ~n13 & ~n19 ;
  assign n21 = ~x7 & n20 ;
  assign n22 = ~x2 & x3 ;
  assign n23 = n22 ^ x5 ;
  assign n24 = x6 & n23 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = n21 & n25 ;
  assign n27 = ~x2 & ~x6 ;
  assign n28 = ~x3 & ~x5 ;
  assign n29 = ~x8 & x9 ;
  assign n30 = n28 & n29 ;
  assign n31 = x3 & n11 ;
  assign n32 = x5 & ~x7 ;
  assign n33 = n31 & n32 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = n30 & n34 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = n27 & n36 ;
  assign n38 = ~n26 & ~n37 ;
  assign n39 = ~n18 & n38 ;
  assign n40 = ~x0 & ~n39 ;
  assign n41 = ~x7 & x9 ;
  assign n42 = x8 & n41 ;
  assign n43 = x6 & ~x7 ;
  assign n44 = ~x2 & ~x5 ;
  assign n45 = ~n43 & n44 ;
  assign n46 = ~n42 & n45 ;
  assign n47 = x3 & n46 ;
  assign n48 = ~n40 & ~n47 ;
  assign n49 = ~x1 & ~n48 ;
  assign n50 = x2 & x3 ;
  assign n51 = x6 & ~n50 ;
  assign n52 = x5 & n50 ;
  assign n53 = ~n51 & ~n52 ;
  assign n54 = ~x5 & ~x6 ;
  assign n55 = ~x0 & ~n54 ;
  assign n56 = x7 & n55 ;
  assign n57 = n53 & n56 ;
  assign n58 = n19 & ~n27 ;
  assign n59 = ~x0 & ~x3 ;
  assign n60 = x8 & n44 ;
  assign n61 = ~x6 & ~n60 ;
  assign n62 = n59 & ~n61 ;
  assign n63 = ~x4 & ~n62 ;
  assign n64 = ~n58 & n63 ;
  assign n65 = ~n57 & n64 ;
  assign n66 = ~n49 & n65 ;
  assign n67 = ~x2 & ~x7 ;
  assign n68 = n28 & n67 ;
  assign n69 = x4 & n68 ;
  assign n70 = ~n66 & ~n69 ;
  assign n71 = ~x3 & n32 ;
  assign n72 = n11 & n71 ;
  assign n73 = ~x0 & ~x5 ;
  assign n74 = n11 ^ x3 ;
  assign n75 = n74 ^ n11 ;
  assign n76 = n13 ^ n11 ;
  assign n77 = ~n75 & n76 ;
  assign n78 = n77 ^ n11 ;
  assign n79 = ~x7 & ~n78 ;
  assign n80 = n73 & ~n79 ;
  assign n81 = ~n72 & ~n80 ;
  assign n82 = n16 & ~n81 ;
  assign n83 = ~x7 & ~n11 ;
  assign n84 = ~x6 & n83 ;
  assign n85 = x5 & ~n84 ;
  assign n86 = ~x0 & n11 ;
  assign n87 = n43 & ~n86 ;
  assign n88 = n22 & ~n87 ;
  assign n89 = ~n85 & n88 ;
  assign n90 = ~x4 & ~n89 ;
  assign n91 = x7 ^ x5 ;
  assign n92 = n13 ^ x7 ;
  assign n93 = n92 ^ n13 ;
  assign n94 = n29 ^ n13 ;
  assign n95 = ~n93 & ~n94 ;
  assign n96 = n95 ^ n13 ;
  assign n97 = n91 & n96 ;
  assign n98 = n27 & n97 ;
  assign n99 = n59 & n98 ;
  assign n100 = n90 & ~n99 ;
  assign n101 = ~n82 & n100 ;
  assign n102 = x1 & ~n101 ;
  assign n103 = ~x5 & x7 ;
  assign n104 = n50 & n103 ;
  assign n105 = ~x4 & ~n104 ;
  assign n106 = x1 & x5 ;
  assign n107 = ~x3 & ~n106 ;
  assign n108 = x5 & x9 ;
  assign n109 = ~x1 & ~n108 ;
  assign n110 = ~n107 & ~n109 ;
  assign n111 = x9 ^ x1 ;
  assign n112 = n111 ^ x8 ;
  assign n113 = x9 ^ x8 ;
  assign n114 = n28 ^ x9 ;
  assign n115 = n113 & ~n114 ;
  assign n116 = n112 & n115 ;
  assign n117 = n116 ^ n111 ;
  assign n118 = x2 & ~n117 ;
  assign n119 = ~n110 & ~n118 ;
  assign n120 = ~x7 & ~n119 ;
  assign n121 = ~n19 & ~n107 ;
  assign n122 = ~x1 & ~x5 ;
  assign n123 = x7 & ~n122 ;
  assign n124 = ~x1 & ~x8 ;
  assign n125 = ~n123 & ~n124 ;
  assign n126 = ~x9 & n125 ;
  assign n127 = ~n121 & ~n126 ;
  assign n128 = ~x2 & ~n127 ;
  assign n129 = x3 & n103 ;
  assign n130 = ~x6 & ~n52 ;
  assign n131 = ~n129 & n130 ;
  assign n132 = ~n128 & n131 ;
  assign n133 = ~n120 & n132 ;
  assign n134 = n51 ^ x3 ;
  assign n135 = n41 & n122 ;
  assign n136 = n135 ^ n51 ;
  assign n137 = n136 ^ n135 ;
  assign n138 = n137 ^ n134 ;
  assign n139 = n106 ^ x2 ;
  assign n140 = ~x2 & ~n139 ;
  assign n141 = n140 ^ n135 ;
  assign n142 = n141 ^ x2 ;
  assign n143 = n138 & n142 ;
  assign n144 = n143 ^ n140 ;
  assign n145 = n144 ^ x2 ;
  assign n146 = ~n134 & ~n145 ;
  assign n147 = n146 ^ n51 ;
  assign n148 = ~n133 & ~n147 ;
  assign n149 = n105 & n148 ;
  assign n150 = x0 & ~n149 ;
  assign n151 = ~n102 & ~n150 ;
  assign n152 = ~n70 & n151 ;
  assign y0 = ~n152 ;
endmodule
