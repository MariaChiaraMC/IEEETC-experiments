module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 ;
  assign n10 = ~x1 & ~x5 ;
  assign n11 = x6 & n10 ;
  assign n12 = x7 & ~n11 ;
  assign n13 = x1 & ~x5 ;
  assign n14 = ~x0 & ~x7 ;
  assign n15 = ~x1 & ~n14 ;
  assign n16 = x6 & n15 ;
  assign n17 = ~n13 & ~n16 ;
  assign n18 = ~x2 & x8 ;
  assign n19 = ~x3 & ~x4 ;
  assign n20 = ~x0 & ~x6 ;
  assign n21 = n19 & ~n20 ;
  assign n22 = n18 & n21 ;
  assign n23 = ~n17 & n22 ;
  assign n24 = ~n12 & n23 ;
  assign n25 = x2 & ~x5 ;
  assign n26 = x3 & x4 ;
  assign n27 = ~x5 & n26 ;
  assign n28 = x2 & n19 ;
  assign n29 = ~n27 & ~n28 ;
  assign n30 = ~n25 & ~n29 ;
  assign n31 = x1 & ~x7 ;
  assign n32 = ~n15 & ~n31 ;
  assign n33 = ~x6 & ~n32 ;
  assign n34 = n30 & n33 ;
  assign n35 = ~x6 & ~x7 ;
  assign n36 = x0 & ~n35 ;
  assign n37 = n19 & n36 ;
  assign n38 = x1 & ~x2 ;
  assign n39 = n37 & n38 ;
  assign n40 = ~x5 & n39 ;
  assign n41 = ~n34 & ~n40 ;
  assign n42 = ~x8 & ~n41 ;
  assign n43 = ~x6 & ~x8 ;
  assign n44 = x6 & x8 ;
  assign n45 = ~n43 & ~n44 ;
  assign n46 = ~x7 & n45 ;
  assign n47 = ~x1 & ~x2 ;
  assign n48 = n27 & n47 ;
  assign n49 = n46 & n48 ;
  assign n50 = ~n42 & ~n49 ;
  assign n51 = ~n24 & n50 ;
  assign n52 = ~x2 & x5 ;
  assign n53 = ~n25 & ~n52 ;
  assign n54 = ~x1 & ~x8 ;
  assign n55 = n35 & n54 ;
  assign n56 = n26 & n55 ;
  assign n57 = ~n19 & ~n26 ;
  assign n58 = ~n14 & n43 ;
  assign n59 = ~n46 & ~n58 ;
  assign n60 = ~x1 & ~n59 ;
  assign n61 = n31 & n43 ;
  assign n62 = ~n60 & ~n61 ;
  assign n63 = n57 & ~n62 ;
  assign n64 = x1 & ~n58 ;
  assign n65 = n19 & ~n64 ;
  assign n66 = ~x7 & ~n20 ;
  assign n67 = n66 ^ x1 ;
  assign n68 = n67 ^ n66 ;
  assign n69 = n66 ^ n36 ;
  assign n70 = n69 ^ n66 ;
  assign n71 = ~n68 & ~n70 ;
  assign n72 = n71 ^ n66 ;
  assign n73 = ~x8 & ~n72 ;
  assign n74 = n73 ^ n66 ;
  assign n75 = n65 & n74 ;
  assign n76 = ~n63 & ~n75 ;
  assign n77 = ~n56 & n76 ;
  assign n78 = ~n53 & ~n77 ;
  assign n79 = x5 ^ x2 ;
  assign n80 = x2 ^ x1 ;
  assign n81 = n80 ^ x5 ;
  assign n82 = n81 ^ x7 ;
  assign n83 = n82 ^ x5 ;
  assign n84 = n83 ^ x7 ;
  assign n85 = ~n79 & ~n84 ;
  assign n86 = x7 ^ x5 ;
  assign n87 = n86 ^ n84 ;
  assign n88 = x0 & x7 ;
  assign n89 = n88 ^ n85 ;
  assign n90 = ~n87 & n89 ;
  assign n91 = n90 ^ n88 ;
  assign n92 = n85 & n91 ;
  assign n93 = n92 ^ n82 ;
  assign n94 = n45 & ~n93 ;
  assign n95 = n94 ^ n26 ;
  assign n96 = n95 ^ n94 ;
  assign n97 = n13 & ~n59 ;
  assign n98 = n44 ^ x7 ;
  assign n100 = n98 ^ n43 ;
  assign n99 = n98 ^ x0 ;
  assign n101 = n100 ^ n99 ;
  assign n102 = n98 ^ n44 ;
  assign n103 = n102 ^ n98 ;
  assign n104 = n103 ^ n100 ;
  assign n105 = ~n100 & n104 ;
  assign n106 = n105 ^ n100 ;
  assign n107 = ~n101 & ~n106 ;
  assign n108 = n107 ^ n105 ;
  assign n109 = n108 ^ n98 ;
  assign n110 = n109 ^ n100 ;
  assign n111 = n10 & ~n110 ;
  assign n112 = ~n97 & ~n111 ;
  assign n113 = ~x2 & ~n112 ;
  assign n114 = ~x1 & x2 ;
  assign n115 = x5 & ~x7 ;
  assign n116 = n43 & n115 ;
  assign n117 = n114 & n116 ;
  assign n118 = ~n113 & ~n117 ;
  assign n119 = n118 ^ n94 ;
  assign n120 = n119 ^ n94 ;
  assign n121 = ~n96 & ~n120 ;
  assign n122 = n121 ^ n94 ;
  assign n123 = ~n19 & n122 ;
  assign n124 = n123 ^ n94 ;
  assign n125 = ~n78 & ~n124 ;
  assign n126 = n51 & n125 ;
  assign y0 = ~n126 ;
endmodule
