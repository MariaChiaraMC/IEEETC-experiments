module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 ;
  assign n17 = x14 & ~x15 ;
  assign n18 = ~x14 & x15 ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = x12 & ~x13 ;
  assign n21 = ~x12 & x13 ;
  assign n22 = ~n20 & ~n21 ;
  assign n23 = n19 & n22 ;
  assign n42 = ~x4 & ~x5 ;
  assign n24 = x8 & ~x9 ;
  assign n25 = x5 & ~x10 ;
  assign n26 = n24 & n25 ;
  assign n27 = ~x11 & n26 ;
  assign n28 = x6 ^ x4 ;
  assign n29 = x6 ^ x5 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = x10 & ~x11 ;
  assign n32 = x11 & n25 ;
  assign n33 = ~n31 & ~n32 ;
  assign n34 = ~x8 & ~x9 ;
  assign n35 = ~n33 & n34 ;
  assign n36 = n35 ^ x5 ;
  assign n37 = ~n30 & ~n36 ;
  assign n38 = n37 ^ x5 ;
  assign n39 = ~n28 & ~n38 ;
  assign n40 = n39 ^ x4 ;
  assign n41 = ~n27 & ~n40 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = n43 ^ x7 ;
  assign n55 = n44 ^ n43 ;
  assign n45 = x7 & ~x10 ;
  assign n46 = ~x8 & ~x11 ;
  assign n47 = n45 & n46 ;
  assign n48 = x9 & n47 ;
  assign n49 = n48 ^ n44 ;
  assign n50 = n49 ^ n43 ;
  assign n51 = n44 ^ n41 ;
  assign n52 = n51 ^ n48 ;
  assign n53 = n52 ^ n50 ;
  assign n54 = ~n50 & n53 ;
  assign n56 = n55 ^ n54 ;
  assign n57 = n56 ^ n50 ;
  assign n58 = x4 & x5 ;
  assign n59 = n58 ^ n43 ;
  assign n60 = n54 ^ n50 ;
  assign n61 = n59 & ~n60 ;
  assign n62 = n61 ^ n43 ;
  assign n63 = ~n57 & n62 ;
  assign n64 = n63 ^ n43 ;
  assign n65 = n64 ^ n42 ;
  assign n66 = n65 ^ n43 ;
  assign n67 = ~n23 & ~n66 ;
  assign n70 = x10 ^ x7 ;
  assign n71 = ~n17 & ~n20 ;
  assign n72 = n71 ^ x10 ;
  assign n73 = n72 ^ n71 ;
  assign n74 = n73 ^ n70 ;
  assign n75 = ~x5 & ~n24 ;
  assign n76 = n75 ^ n23 ;
  assign n77 = ~n75 & n76 ;
  assign n78 = n77 ^ n71 ;
  assign n79 = n78 ^ n75 ;
  assign n80 = ~n74 & n79 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n81 ^ n75 ;
  assign n83 = n70 & ~n82 ;
  assign n84 = ~x11 & n83 ;
  assign n87 = x13 ^ x12 ;
  assign n88 = n87 ^ x14 ;
  assign n89 = n88 ^ x15 ;
  assign n90 = x15 ^ x13 ;
  assign n91 = x14 ^ x13 ;
  assign n92 = n90 & n91 ;
  assign n93 = n92 ^ x13 ;
  assign n94 = n89 & n93 ;
  assign n95 = n32 & n94 ;
  assign n85 = n42 ^ x7 ;
  assign n86 = n85 ^ n42 ;
  assign n96 = n95 ^ n86 ;
  assign n97 = n96 ^ n95 ;
  assign n98 = n97 ^ n85 ;
  assign n99 = n98 ^ n97 ;
  assign n100 = n24 & ~n99 ;
  assign n101 = n100 ^ n95 ;
  assign n102 = n95 ^ n31 ;
  assign n103 = n98 & ~n102 ;
  assign n104 = n103 ^ n97 ;
  assign n105 = n104 ^ n98 ;
  assign n106 = ~n101 & ~n105 ;
  assign n107 = ~n97 & n106 ;
  assign n108 = n107 ^ n100 ;
  assign n109 = n108 ^ x7 ;
  assign n110 = ~n84 & n109 ;
  assign n68 = x7 & n31 ;
  assign n69 = n42 & n68 ;
  assign n111 = n110 ^ n69 ;
  assign n112 = ~x6 & ~n111 ;
  assign n113 = n112 ^ n110 ;
  assign n114 = ~n67 & n113 ;
  assign n115 = ~x0 & ~x3 ;
  assign n116 = ~x1 & n115 ;
  assign n117 = ~x2 & n116 ;
  assign n118 = ~n114 & n117 ;
  assign y0 = n118 ;
endmodule
