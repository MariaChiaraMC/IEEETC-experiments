module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 ;
  assign n17 = ~x2 & ~x3 ;
  assign n18 = ~x0 & ~x1 ;
  assign n19 = n17 & n18 ;
  assign n20 = x12 & x13 ;
  assign n21 = x14 & x15 ;
  assign n22 = ~n20 & ~n21 ;
  assign n31 = x7 ^ x4 ;
  assign n25 = ~x5 & x6 ;
  assign n26 = ~x8 & ~x9 ;
  assign n27 = n25 & n26 ;
  assign n28 = x11 ^ x10 ;
  assign n29 = n27 & n28 ;
  assign n32 = n31 ^ n29 ;
  assign n23 = x6 ^ x4 ;
  assign n24 = n23 ^ x5 ;
  assign n30 = n29 ^ n24 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n32 ^ x5 ;
  assign n35 = n33 ^ x4 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = n34 & n36 ;
  assign n38 = n37 ^ n32 ;
  assign n39 = n32 ^ n29 ;
  assign n40 = n35 & ~n39 ;
  assign n41 = n40 ^ n33 ;
  assign n42 = n41 ^ n35 ;
  assign n43 = ~n38 & n42 ;
  assign n44 = n33 & n43 ;
  assign n45 = n44 ^ n37 ;
  assign n46 = n45 ^ n29 ;
  assign n47 = ~n22 & n46 ;
  assign n48 = x12 & x14 ;
  assign n49 = x4 & x5 ;
  assign n50 = n48 & n49 ;
  assign n51 = x13 & x15 ;
  assign n52 = x6 & ~x10 ;
  assign n53 = n51 & n52 ;
  assign n54 = n50 & n53 ;
  assign n55 = x11 & n54 ;
  assign n56 = x10 & x11 ;
  assign n57 = n48 & ~n51 ;
  assign n58 = x10 & ~n57 ;
  assign n59 = ~n56 & ~n58 ;
  assign n60 = x6 & ~n22 ;
  assign n61 = x5 ^ x4 ;
  assign n62 = ~x10 & ~x11 ;
  assign n63 = n62 ^ x5 ;
  assign n64 = ~n61 & n63 ;
  assign n65 = n60 & n64 ;
  assign n66 = n59 & n65 ;
  assign n67 = x5 & ~x6 ;
  assign n68 = ~x12 & n67 ;
  assign n69 = ~x15 & n68 ;
  assign n70 = ~x7 & ~n69 ;
  assign n71 = x11 & ~n70 ;
  assign n73 = x12 & x15 ;
  assign n74 = x7 & ~n73 ;
  assign n72 = x7 & n67 ;
  assign n75 = n74 ^ n72 ;
  assign n76 = n75 ^ n72 ;
  assign n77 = ~x13 & x14 ;
  assign n78 = n77 ^ n72 ;
  assign n79 = n78 ^ n72 ;
  assign n80 = ~n76 & n79 ;
  assign n81 = n80 ^ n72 ;
  assign n82 = x4 & n81 ;
  assign n83 = n82 ^ n72 ;
  assign n84 = n71 & n83 ;
  assign n85 = ~n66 & ~n84 ;
  assign n86 = x9 ^ x8 ;
  assign n87 = ~n85 & n86 ;
  assign n88 = ~n55 & ~n87 ;
  assign n89 = ~n47 & n88 ;
  assign n90 = n19 & ~n89 ;
  assign y0 = n90 ;
endmodule
