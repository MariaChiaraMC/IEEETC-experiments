module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 ;
  assign n16 = x12 ^ x11 ;
  assign n17 = ~x0 & ~x2 ;
  assign n18 = x1 & n17 ;
  assign n21 = n18 ^ x3 ;
  assign n19 = ~x2 & x4 ;
  assign n20 = n19 ^ n18 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n20 ^ n18 ;
  assign n24 = n23 ^ x13 ;
  assign n25 = n22 & ~n24 ;
  assign n26 = n25 ^ n18 ;
  assign n27 = x0 & ~x1 ;
  assign n28 = ~n18 & n27 ;
  assign n29 = n28 ^ x13 ;
  assign n30 = ~n26 & ~n29 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = ~x13 & n31 ;
  assign n33 = n32 ^ n25 ;
  assign n34 = n33 ^ n18 ;
  assign n35 = n34 ^ n18 ;
  assign n36 = ~x10 & ~n35 ;
  assign n37 = ~x9 & n36 ;
  assign n38 = x10 & ~x13 ;
  assign n39 = ~x2 & ~x3 ;
  assign n40 = n27 & ~n39 ;
  assign n41 = n40 ^ x9 ;
  assign n42 = x14 ^ x9 ;
  assign n43 = n42 ^ x9 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = ~n41 & n44 ;
  assign n46 = n45 ^ n40 ;
  assign n47 = n38 & n46 ;
  assign n48 = n47 ^ x10 ;
  assign n49 = ~n37 & ~n48 ;
  assign n50 = n49 ^ x12 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = n51 ^ n16 ;
  assign n53 = n38 ^ x9 ;
  assign n54 = n38 & n53 ;
  assign n55 = n54 ^ n49 ;
  assign n56 = n55 ^ n38 ;
  assign n57 = ~n52 & ~n56 ;
  assign n58 = n57 ^ n54 ;
  assign n59 = n58 ^ n38 ;
  assign n60 = ~n16 & n59 ;
  assign y0 = n60 ;
endmodule
