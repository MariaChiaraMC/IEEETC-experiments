module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 ;
  assign n9 = ~x5 & x7 ;
  assign n10 = x4 ^ x3 ;
  assign n11 = x3 ^ x2 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = x4 ^ x0 ;
  assign n14 = n13 ^ x0 ;
  assign n15 = x1 ^ x0 ;
  assign n16 = n14 & n15 ;
  assign n17 = n16 ^ x0 ;
  assign n18 = n17 ^ n10 ;
  assign n19 = n12 & ~n18 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = n20 ^ x0 ;
  assign n22 = n21 ^ n11 ;
  assign n23 = n10 & ~n22 ;
  assign n24 = n23 ^ n10 ;
  assign n25 = n9 & n24 ;
  assign n26 = ~x2 & ~x4 ;
  assign n27 = x5 & x7 ;
  assign n28 = ~x0 & n27 ;
  assign n29 = n26 & n28 ;
  assign n30 = x5 & ~x7 ;
  assign n31 = x2 & ~n30 ;
  assign n32 = n31 ^ x4 ;
  assign n33 = x3 & ~x5 ;
  assign n34 = ~x5 & ~x7 ;
  assign n35 = ~n33 & ~n34 ;
  assign n36 = ~x3 & n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ n31 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = n39 ^ n32 ;
  assign n41 = n33 ^ x3 ;
  assign n42 = x7 & ~n41 ;
  assign n43 = n42 ^ x3 ;
  assign n44 = ~x3 & x5 ;
  assign n45 = n44 ^ n43 ;
  assign n46 = n43 & ~n45 ;
  assign n47 = n46 ^ n37 ;
  assign n48 = n47 ^ n43 ;
  assign n49 = n40 & ~n48 ;
  assign n50 = n49 ^ n46 ;
  assign n51 = n50 ^ n43 ;
  assign n52 = n32 & n51 ;
  assign n53 = n52 ^ x0 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = x4 & ~x7 ;
  assign n56 = x2 & x3 ;
  assign n57 = n56 ^ x2 ;
  assign n58 = n55 & ~n57 ;
  assign n59 = n58 ^ x2 ;
  assign n60 = ~n35 & ~n59 ;
  assign n61 = n60 ^ n52 ;
  assign n62 = ~n54 & n61 ;
  assign n63 = n62 ^ n52 ;
  assign n64 = ~n29 & ~n63 ;
  assign n65 = x1 & ~n64 ;
  assign n66 = ~x6 & ~n65 ;
  assign n67 = ~n25 & n66 ;
  assign n68 = ~x3 & ~x5 ;
  assign n69 = ~x1 & ~x2 ;
  assign n70 = n55 & n69 ;
  assign n71 = n68 & n70 ;
  assign n72 = x6 & ~n71 ;
  assign n73 = ~x3 & x4 ;
  assign n74 = n69 & n73 ;
  assign n75 = n27 & n74 ;
  assign n76 = x2 ^ x1 ;
  assign n77 = n68 ^ x5 ;
  assign n78 = n77 ^ x5 ;
  assign n79 = x5 ^ x2 ;
  assign n80 = n79 ^ x5 ;
  assign n81 = n78 & n80 ;
  assign n82 = n81 ^ x5 ;
  assign n83 = ~n76 & n82 ;
  assign n84 = n83 ^ x5 ;
  assign n85 = n55 & n84 ;
  assign n86 = ~x4 & ~n44 ;
  assign n87 = n31 & n86 ;
  assign n88 = ~n9 & ~n33 ;
  assign n89 = n88 ^ x1 ;
  assign n90 = n87 & n89 ;
  assign n91 = ~n85 & ~n90 ;
  assign n92 = ~n75 & n91 ;
  assign n93 = n92 ^ x0 ;
  assign n94 = n93 ^ n92 ;
  assign n95 = x1 & ~x2 ;
  assign n96 = n33 & n95 ;
  assign n97 = n56 ^ x1 ;
  assign n98 = n30 ^ n9 ;
  assign n99 = n9 ^ x4 ;
  assign n100 = n99 ^ n9 ;
  assign n101 = n98 & ~n100 ;
  assign n102 = n101 ^ n9 ;
  assign n103 = n102 ^ n56 ;
  assign n104 = ~n97 & n103 ;
  assign n105 = n104 ^ n101 ;
  assign n106 = n105 ^ n9 ;
  assign n107 = n106 ^ x1 ;
  assign n108 = n56 & ~n107 ;
  assign n109 = n108 ^ n56 ;
  assign n110 = ~n96 & ~n109 ;
  assign n111 = ~x3 & ~x4 ;
  assign n112 = n9 ^ x1 ;
  assign n113 = n112 ^ n9 ;
  assign n114 = n98 & n113 ;
  assign n115 = n114 ^ n9 ;
  assign n116 = n111 & n115 ;
  assign n117 = n110 & ~n116 ;
  assign n118 = n117 ^ n92 ;
  assign n119 = n94 & n118 ;
  assign n120 = n119 ^ n92 ;
  assign n121 = n72 & n120 ;
  assign n122 = ~n67 & ~n121 ;
  assign n123 = n28 & n111 ;
  assign n124 = n95 & n123 ;
  assign n125 = ~n122 & ~n124 ;
  assign y0 = ~n125 ;
endmodule
