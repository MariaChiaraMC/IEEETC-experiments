module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 ;
  assign n10 = ~x5 & x7 ;
  assign n11 = ~x3 & x4 ;
  assign n12 = x2 & n11 ;
  assign n13 = n10 & n12 ;
  assign n14 = x4 & x7 ;
  assign n15 = ~x2 & n14 ;
  assign n16 = ~x0 & n15 ;
  assign n17 = x5 & n16 ;
  assign n18 = ~x3 & ~x7 ;
  assign n19 = ~x4 & ~x5 ;
  assign n20 = ~x0 & n19 ;
  assign n21 = n18 & n20 ;
  assign n22 = ~n17 & ~n21 ;
  assign n23 = x0 & ~x3 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n24 ^ x2 ;
  assign n26 = x7 ^ x5 ;
  assign n27 = n26 ^ x8 ;
  assign n28 = x8 & ~n27 ;
  assign n29 = n28 ^ x5 ;
  assign n30 = n29 ^ x8 ;
  assign n31 = n25 & ~n30 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = n32 ^ x8 ;
  assign n34 = ~x2 & n33 ;
  assign n35 = n34 ^ x4 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = x2 & ~x5 ;
  assign n38 = ~x0 & x7 ;
  assign n39 = x8 & n38 ;
  assign n40 = x3 & ~n39 ;
  assign n41 = n37 & ~n40 ;
  assign n42 = x7 ^ x2 ;
  assign n43 = n42 ^ x2 ;
  assign n44 = x0 & x2 ;
  assign n45 = n44 ^ x2 ;
  assign n46 = n43 & ~n45 ;
  assign n47 = n46 ^ x2 ;
  assign n48 = x5 & ~n47 ;
  assign n49 = ~n41 & ~n48 ;
  assign n50 = n49 ^ n34 ;
  assign n51 = n36 & ~n50 ;
  assign n52 = n51 ^ n34 ;
  assign n53 = x6 & n52 ;
  assign n54 = n22 & ~n53 ;
  assign n55 = ~n13 & n54 ;
  assign n56 = ~x1 & ~n55 ;
  assign n57 = x1 & n44 ;
  assign n58 = ~n19 & n57 ;
  assign n59 = ~x1 & x5 ;
  assign n60 = x8 & n59 ;
  assign n61 = ~x0 & x4 ;
  assign n62 = ~n14 & ~n61 ;
  assign n63 = n60 & ~n62 ;
  assign n64 = ~x1 & ~x2 ;
  assign n65 = n20 & n64 ;
  assign n66 = x4 & x5 ;
  assign n67 = x2 & x8 ;
  assign n68 = n66 & n67 ;
  assign n69 = ~x7 & n68 ;
  assign n70 = ~n65 & ~n69 ;
  assign n71 = ~n63 & n70 ;
  assign n72 = ~n58 & n71 ;
  assign n73 = x3 & ~n72 ;
  assign n74 = ~n56 & ~n73 ;
  assign n75 = x0 & x4 ;
  assign n76 = x7 & x8 ;
  assign n77 = ~n14 & ~n76 ;
  assign n78 = ~n75 & ~n77 ;
  assign n79 = x1 & ~x3 ;
  assign n80 = x5 & n79 ;
  assign n81 = ~n78 & n80 ;
  assign n82 = ~x2 & n81 ;
  assign n83 = n82 ^ n74 ;
  assign n91 = ~x0 & ~x3 ;
  assign n92 = ~x1 & ~x5 ;
  assign n93 = n91 & n92 ;
  assign n94 = n76 & n79 ;
  assign n95 = ~x0 & ~n94 ;
  assign n87 = x1 & x7 ;
  assign n96 = ~x7 & ~x8 ;
  assign n97 = n64 & n96 ;
  assign n98 = ~n87 & ~n97 ;
  assign n99 = ~n95 & ~n98 ;
  assign n100 = ~x0 & ~x8 ;
  assign n101 = ~x7 & x8 ;
  assign n102 = ~n100 & ~n101 ;
  assign n103 = x3 & ~n102 ;
  assign n104 = ~x2 & n103 ;
  assign n105 = ~n99 & ~n104 ;
  assign n106 = x5 & ~n105 ;
  assign n107 = ~n93 & ~n106 ;
  assign n84 = x3 & ~x7 ;
  assign n85 = ~n64 & ~n84 ;
  assign n86 = x0 & ~n85 ;
  assign n88 = x3 & n87 ;
  assign n89 = ~n67 & n88 ;
  assign n90 = ~n86 & ~n89 ;
  assign n108 = n107 ^ n90 ;
  assign n109 = n108 ^ n107 ;
  assign n110 = n107 ^ x5 ;
  assign n111 = n110 ^ n107 ;
  assign n112 = ~n109 & ~n111 ;
  assign n113 = n112 ^ n107 ;
  assign n114 = x4 & ~n113 ;
  assign n115 = n114 ^ n107 ;
  assign n116 = x0 & ~x4 ;
  assign n117 = ~x1 & x3 ;
  assign n118 = n117 ^ x3 ;
  assign n119 = ~x5 & ~n118 ;
  assign n120 = n119 ^ x3 ;
  assign n121 = n116 & ~n120 ;
  assign n122 = x3 & x7 ;
  assign n123 = n116 & n122 ;
  assign n124 = ~n93 & ~n123 ;
  assign n125 = x8 & ~n124 ;
  assign n126 = ~x0 & x1 ;
  assign n127 = ~n96 & ~n126 ;
  assign n128 = ~n79 & n127 ;
  assign n129 = n19 & ~n84 ;
  assign n130 = ~n128 & n129 ;
  assign n131 = ~n125 & ~n130 ;
  assign n151 = n91 & n96 ;
  assign n152 = x4 & n84 ;
  assign n153 = ~n151 & ~n152 ;
  assign n132 = n14 ^ x0 ;
  assign n133 = n132 ^ x3 ;
  assign n140 = n133 ^ n132 ;
  assign n134 = n133 ^ n117 ;
  assign n135 = n134 ^ n132 ;
  assign n136 = n133 ^ n14 ;
  assign n137 = n136 ^ n117 ;
  assign n138 = n137 ^ n135 ;
  assign n139 = ~n135 & n138 ;
  assign n141 = n140 ^ n139 ;
  assign n142 = n141 ^ n135 ;
  assign n143 = n132 ^ x4 ;
  assign n144 = n139 ^ n135 ;
  assign n145 = n143 & ~n144 ;
  assign n146 = n145 ^ n132 ;
  assign n147 = ~n142 & ~n146 ;
  assign n148 = n147 ^ n132 ;
  assign n149 = n148 ^ x0 ;
  assign n150 = n149 ^ n132 ;
  assign n154 = n153 ^ n150 ;
  assign n155 = n154 ^ n150 ;
  assign n156 = n150 ^ x1 ;
  assign n157 = n156 ^ n150 ;
  assign n158 = ~n155 & n157 ;
  assign n159 = n158 ^ n150 ;
  assign n160 = ~x5 & ~n159 ;
  assign n161 = n160 ^ n150 ;
  assign n162 = n131 & n161 ;
  assign n163 = ~n121 & n162 ;
  assign n164 = n163 ^ x2 ;
  assign n165 = n164 ^ n163 ;
  assign n166 = n165 ^ n115 ;
  assign n167 = ~x3 & x5 ;
  assign n168 = n167 ^ n14 ;
  assign n169 = n14 & n168 ;
  assign n170 = n169 ^ n163 ;
  assign n171 = n170 ^ n14 ;
  assign n172 = ~n166 & ~n171 ;
  assign n173 = n172 ^ n169 ;
  assign n174 = n173 ^ n14 ;
  assign n175 = n115 & n174 ;
  assign n176 = n175 ^ n115 ;
  assign n177 = n176 ^ x6 ;
  assign n178 = n177 ^ n176 ;
  assign n179 = n75 & n97 ;
  assign n180 = x0 & ~n64 ;
  assign n181 = n10 & ~n180 ;
  assign n182 = x2 & ~x7 ;
  assign n183 = x8 ^ x0 ;
  assign n184 = n182 & n183 ;
  assign n185 = ~n181 & ~n184 ;
  assign n186 = ~x4 & ~n185 ;
  assign n187 = x1 & x5 ;
  assign n188 = n116 & n187 ;
  assign n189 = ~n186 & ~n188 ;
  assign n190 = x4 & n182 ;
  assign n191 = ~x1 & x2 ;
  assign n192 = ~x8 & n191 ;
  assign n193 = ~n190 & ~n192 ;
  assign n194 = ~n16 & n193 ;
  assign n195 = ~n44 & n194 ;
  assign n196 = n195 ^ n126 ;
  assign n197 = n196 ^ n195 ;
  assign n198 = n195 ^ x2 ;
  assign n199 = n198 ^ n195 ;
  assign n200 = n197 & ~n199 ;
  assign n201 = n200 ^ n195 ;
  assign n202 = ~x5 & ~n201 ;
  assign n203 = n202 ^ n195 ;
  assign n204 = n189 & n203 ;
  assign n205 = ~n179 & n204 ;
  assign n206 = x3 & ~n205 ;
  assign n207 = n37 & n116 ;
  assign n208 = ~x1 & ~x7 ;
  assign n209 = ~n117 & ~n208 ;
  assign n210 = n207 & n209 ;
  assign n211 = n15 & n126 ;
  assign n212 = n94 ^ x2 ;
  assign n213 = n212 ^ n94 ;
  assign n214 = n213 ^ n211 ;
  assign n215 = n39 ^ n11 ;
  assign n216 = n11 & n215 ;
  assign n217 = n216 ^ n94 ;
  assign n218 = n217 ^ n11 ;
  assign n219 = ~n214 & n218 ;
  assign n220 = n219 ^ n216 ;
  assign n221 = n220 ^ n11 ;
  assign n222 = ~n211 & n221 ;
  assign n223 = n222 ^ n211 ;
  assign n224 = ~x5 & n223 ;
  assign n225 = n19 & n182 ;
  assign n226 = n225 ^ x2 ;
  assign n227 = n226 ^ n225 ;
  assign n228 = n225 ^ n66 ;
  assign n229 = n228 ^ n225 ;
  assign n230 = ~n227 & n229 ;
  assign n231 = n230 ^ n225 ;
  assign n232 = ~x1 & n231 ;
  assign n233 = n232 ^ n225 ;
  assign n234 = ~x8 & n233 ;
  assign n235 = x2 & n38 ;
  assign n236 = ~n18 & ~n235 ;
  assign n237 = ~x4 & n187 ;
  assign n238 = ~n236 & n237 ;
  assign n239 = ~n234 & ~n238 ;
  assign n240 = ~n224 & n239 ;
  assign n241 = ~n210 & n240 ;
  assign n242 = ~n206 & n241 ;
  assign n243 = n242 ^ n176 ;
  assign n244 = n178 & n243 ;
  assign n245 = n244 ^ n176 ;
  assign n246 = n245 ^ n74 ;
  assign n247 = ~n83 & n246 ;
  assign n248 = n247 ^ n244 ;
  assign n249 = n248 ^ n176 ;
  assign n250 = n249 ^ n82 ;
  assign n251 = n74 & ~n250 ;
  assign n252 = n251 ^ n74 ;
  assign y0 = ~n252 ;
endmodule
