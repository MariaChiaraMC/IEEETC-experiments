module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 ;
  assign n11 = ~x0 & ~x6 ;
  assign n12 = x2 & x3 ;
  assign n13 = ~n11 & n12 ;
  assign n14 = ~x7 & ~n13 ;
  assign n15 = ~x8 & n14 ;
  assign n16 = x3 & x6 ;
  assign n17 = n15 & ~n16 ;
  assign n18 = x5 & ~x9 ;
  assign n19 = ~x1 & ~n18 ;
  assign n20 = ~x4 & ~x8 ;
  assign n21 = n19 & ~n20 ;
  assign n22 = ~n17 & n21 ;
  assign n23 = ~x8 & ~n18 ;
  assign n24 = ~x4 & ~n23 ;
  assign n25 = ~x2 & x6 ;
  assign n26 = ~n24 & ~n25 ;
  assign n27 = ~n22 & n26 ;
  assign n28 = x9 ^ x5 ;
  assign n29 = ~x1 & ~n15 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = ~x3 & x7 ;
  assign n32 = n31 ^ x5 ;
  assign n33 = x5 & ~n32 ;
  assign n34 = n33 ^ x5 ;
  assign n35 = n30 & n34 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = n36 ^ x5 ;
  assign n38 = n37 ^ n31 ;
  assign n39 = n28 & ~n38 ;
  assign n40 = n39 ^ n31 ;
  assign n41 = n27 & ~n40 ;
  assign y0 = n41 ;
endmodule
