module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 ;
  assign n9 = x6 & x7 ;
  assign n10 = x1 & ~x4 ;
  assign n11 = n10 ^ x2 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = n10 ^ x1 ;
  assign n14 = n13 ^ n10 ;
  assign n15 = ~n12 & ~n14 ;
  assign n16 = n15 ^ n10 ;
  assign n17 = x5 & n16 ;
  assign n18 = n17 ^ n10 ;
  assign n19 = ~n9 & n18 ;
  assign n20 = ~x1 & x5 ;
  assign n21 = ~x4 & x6 ;
  assign n22 = x2 & n21 ;
  assign n23 = n20 & n22 ;
  assign n24 = x2 & x4 ;
  assign n25 = x4 ^ x0 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n20 ^ n9 ;
  assign n28 = x4 & ~n27 ;
  assign n29 = n28 ^ n9 ;
  assign n30 = ~n26 & n29 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n31 ^ n9 ;
  assign n33 = n32 ^ x4 ;
  assign n34 = ~n24 & n33 ;
  assign n35 = ~n23 & ~n34 ;
  assign n36 = ~n19 & n35 ;
  assign n37 = x3 & ~n36 ;
  assign n38 = x3 ^ x1 ;
  assign n39 = x3 ^ x0 ;
  assign n40 = n39 ^ x3 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = ~x6 & ~x7 ;
  assign n43 = n42 ^ x2 ;
  assign n44 = x3 & n43 ;
  assign n45 = n44 ^ n42 ;
  assign n46 = n41 & n45 ;
  assign n47 = n46 ^ n44 ;
  assign n48 = n47 ^ n42 ;
  assign n49 = n48 ^ x3 ;
  assign n50 = ~n38 & n49 ;
  assign n51 = n50 ^ x1 ;
  assign n52 = x4 & n51 ;
  assign n53 = x4 ^ x3 ;
  assign n54 = n53 ^ x3 ;
  assign n56 = x1 & x2 ;
  assign n55 = n54 ^ n53 ;
  assign n57 = n56 ^ n55 ;
  assign n58 = ~n54 & ~n57 ;
  assign n59 = n58 ^ n53 ;
  assign n60 = n59 ^ n54 ;
  assign n64 = n54 ^ x6 ;
  assign n65 = ~n54 & n64 ;
  assign n61 = n53 ^ x5 ;
  assign n62 = n61 ^ n54 ;
  assign n63 = n42 & ~n62 ;
  assign n66 = n65 ^ n63 ;
  assign n67 = n66 ^ n53 ;
  assign n68 = n67 ^ x5 ;
  assign n69 = n68 ^ n54 ;
  assign n70 = n69 ^ n56 ;
  assign n71 = ~x5 & n70 ;
  assign n72 = n71 ^ n63 ;
  assign n73 = n72 ^ n53 ;
  assign n74 = n73 ^ n54 ;
  assign n75 = n74 ^ n56 ;
  assign n76 = n60 & ~n75 ;
  assign n77 = n76 ^ n63 ;
  assign n78 = n77 ^ n58 ;
  assign n79 = n78 ^ n71 ;
  assign n80 = n79 ^ n56 ;
  assign n81 = ~n52 & ~n80 ;
  assign n82 = ~n37 & n81 ;
  assign n83 = x4 ^ x2 ;
  assign n84 = x1 & ~n83 ;
  assign n85 = n84 ^ x2 ;
  assign n86 = x0 & n85 ;
  assign n87 = x5 ^ x2 ;
  assign n88 = x5 ^ x0 ;
  assign n89 = n88 ^ x0 ;
  assign n90 = n89 ^ n87 ;
  assign n91 = x6 ^ x4 ;
  assign n92 = x4 & ~n91 ;
  assign n93 = n92 ^ x0 ;
  assign n94 = n93 ^ x4 ;
  assign n95 = ~n90 & n94 ;
  assign n96 = n95 ^ n92 ;
  assign n97 = n96 ^ x4 ;
  assign n98 = ~n87 & n97 ;
  assign n99 = n98 ^ x5 ;
  assign n100 = n99 ^ x1 ;
  assign n101 = x3 & ~n24 ;
  assign n102 = n101 ^ n21 ;
  assign n103 = n102 ^ n101 ;
  assign n104 = n101 ^ x2 ;
  assign n105 = n103 & n104 ;
  assign n106 = n105 ^ n101 ;
  assign n107 = n106 ^ n99 ;
  assign n108 = n100 & n107 ;
  assign n109 = n108 ^ n105 ;
  assign n110 = n109 ^ n101 ;
  assign n111 = n110 ^ x1 ;
  assign n112 = ~n99 & n111 ;
  assign n113 = n112 ^ n99 ;
  assign n114 = ~n86 & n113 ;
  assign n115 = n82 & n114 ;
  assign y0 = ~n115 ;
endmodule
