module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 ;
  assign n9 = x3 & ~x4 ;
  assign n10 = ~x1 & ~x2 ;
  assign n11 = ~x5 & x7 ;
  assign n12 = n10 & n11 ;
  assign n13 = n9 & n12 ;
  assign n28 = x4 & ~x5 ;
  assign n14 = x2 & x3 ;
  assign n15 = ~x2 & ~x3 ;
  assign n16 = x7 & n15 ;
  assign n17 = ~n14 & ~n16 ;
  assign n18 = x1 & x5 ;
  assign n19 = ~n17 & n18 ;
  assign n20 = ~x4 & ~n12 ;
  assign n21 = ~n19 & n20 ;
  assign n22 = ~x5 & n16 ;
  assign n23 = x5 & n14 ;
  assign n24 = ~x1 & n23 ;
  assign n25 = x4 & ~n24 ;
  assign n26 = ~n22 & n25 ;
  assign n27 = ~n21 & ~n26 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = x1 & n15 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = n32 ^ n27 ;
  assign n34 = n30 & n33 ;
  assign n35 = n34 ^ n27 ;
  assign n36 = x6 & n35 ;
  assign n37 = n36 ^ n27 ;
  assign n38 = ~n13 & ~n37 ;
  assign n39 = x0 & ~n38 ;
  assign n40 = ~x4 & ~x5 ;
  assign n41 = ~x6 & n40 ;
  assign n84 = n41 ^ x0 ;
  assign n87 = x4 & x6 ;
  assign n88 = x5 & ~n87 ;
  assign n85 = n84 ^ x3 ;
  assign n86 = n85 ^ n41 ;
  assign n89 = n88 ^ n86 ;
  assign n90 = n89 ^ n86 ;
  assign n91 = n86 ^ n41 ;
  assign n92 = n91 ^ n84 ;
  assign n93 = ~n90 & n92 ;
  assign n94 = n93 ^ n41 ;
  assign n95 = x6 & n28 ;
  assign n96 = ~n41 & n95 ;
  assign n97 = n96 ^ n84 ;
  assign n98 = ~n94 & n97 ;
  assign n99 = n98 ^ n96 ;
  assign n100 = n84 & n99 ;
  assign n101 = n100 ^ n93 ;
  assign n102 = n101 ^ x0 ;
  assign n103 = n102 ^ n41 ;
  assign n104 = ~x2 & n103 ;
  assign n105 = ~x0 & ~x6 ;
  assign n106 = n28 & n105 ;
  assign n107 = x3 & n106 ;
  assign n108 = ~n104 & ~n107 ;
  assign n42 = n14 & n41 ;
  assign n43 = x3 ^ x2 ;
  assign n44 = n43 ^ x4 ;
  assign n45 = n44 ^ x0 ;
  assign n46 = n45 ^ x6 ;
  assign n47 = n46 ^ x4 ;
  assign n48 = n47 ^ x2 ;
  assign n49 = n48 ^ x5 ;
  assign n50 = n49 ^ x2 ;
  assign n51 = n50 ^ x5 ;
  assign n60 = n51 ^ n49 ;
  assign n54 = x4 ^ x0 ;
  assign n55 = n54 ^ x6 ;
  assign n62 = n55 ^ x6 ;
  assign n63 = n62 ^ x4 ;
  assign n56 = n55 ^ x2 ;
  assign n61 = n56 ^ x5 ;
  assign n64 = n63 ^ n61 ;
  assign n65 = n60 & ~n64 ;
  assign n52 = n51 ^ x5 ;
  assign n53 = n49 ^ x4 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n57 ^ n51 ;
  assign n59 = ~n52 & n58 ;
  assign n66 = n65 ^ n59 ;
  assign n67 = n66 ^ x5 ;
  assign n68 = n67 ^ n53 ;
  assign n69 = n68 ^ n51 ;
  assign n70 = n53 ^ n51 ;
  assign n71 = n70 ^ n49 ;
  assign n72 = ~n51 & ~n71 ;
  assign n73 = n72 ^ x5 ;
  assign n74 = n73 ^ n51 ;
  assign n75 = n59 ^ n56 ;
  assign n76 = n75 ^ n53 ;
  assign n77 = n76 ^ n49 ;
  assign n78 = ~n74 & n77 ;
  assign n79 = n78 ^ x5 ;
  assign n80 = n69 & n79 ;
  assign n81 = n80 ^ n78 ;
  assign n82 = n81 ^ x5 ;
  assign n83 = ~n42 & ~n82 ;
  assign n109 = n108 ^ n83 ;
  assign n110 = n109 ^ n83 ;
  assign n111 = x5 & n87 ;
  assign n112 = ~n41 & ~n111 ;
  assign n113 = x0 & x2 ;
  assign n114 = ~x3 & n113 ;
  assign n115 = ~n112 & n114 ;
  assign n116 = n115 ^ n83 ;
  assign n117 = n116 ^ n83 ;
  assign n118 = n110 & ~n117 ;
  assign n119 = n118 ^ n83 ;
  assign n120 = x1 & n119 ;
  assign n121 = n120 ^ n83 ;
  assign n122 = n121 ^ x7 ;
  assign n123 = n122 ^ n121 ;
  assign n138 = x6 & n40 ;
  assign n139 = x5 & ~x6 ;
  assign n140 = x2 & x4 ;
  assign n141 = ~x0 & n140 ;
  assign n142 = n139 & n141 ;
  assign n143 = ~n138 & ~n142 ;
  assign n124 = ~x2 & ~x6 ;
  assign n125 = n124 ^ x4 ;
  assign n126 = n124 ^ x5 ;
  assign n127 = n126 ^ x5 ;
  assign n128 = n127 ^ n125 ;
  assign n129 = x6 ^ x5 ;
  assign n130 = n129 ^ n113 ;
  assign n131 = ~n113 & n130 ;
  assign n132 = n131 ^ x5 ;
  assign n133 = n132 ^ n113 ;
  assign n134 = n128 & n133 ;
  assign n135 = n134 ^ n131 ;
  assign n136 = n135 ^ n113 ;
  assign n137 = ~n125 & ~n136 ;
  assign n144 = n143 ^ n137 ;
  assign n145 = n144 ^ n137 ;
  assign n146 = x0 & ~x2 ;
  assign n147 = n146 ^ n137 ;
  assign n148 = n147 ^ n137 ;
  assign n149 = ~n145 & ~n148 ;
  assign n150 = n149 ^ n137 ;
  assign n151 = x1 & n150 ;
  assign n152 = n151 ^ n137 ;
  assign n153 = ~x3 & n152 ;
  assign n154 = x0 & x6 ;
  assign n155 = ~x4 & n154 ;
  assign n156 = n24 & n155 ;
  assign n157 = ~x5 & x6 ;
  assign n158 = ~x1 & n141 ;
  assign n159 = n157 & n158 ;
  assign n160 = ~n156 & ~n159 ;
  assign n161 = ~n153 & n160 ;
  assign n162 = n161 ^ n121 ;
  assign n163 = n123 & n162 ;
  assign n164 = n163 ^ n121 ;
  assign n165 = ~n39 & n164 ;
  assign y0 = ~n165 ;
endmodule
