module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n10 = x3 & x4 ;
  assign n16 = ~x0 & x1 ;
  assign n17 = n10 & n16 ;
  assign n9 = x0 & ~x1 ;
  assign n11 = ~x5 & ~x6 ;
  assign n12 = n10 & ~n11 ;
  assign n13 = n9 & ~n12 ;
  assign n14 = n13 ^ x2 ;
  assign n15 = n14 ^ n11 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n15 ^ n14 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = n19 & n21 ;
  assign n23 = n22 ^ n14 ;
  assign n24 = ~x7 & ~n14 ;
  assign n25 = n24 ^ x2 ;
  assign n26 = ~n23 & ~n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = ~x2 & n27 ;
  assign n29 = n28 ^ n22 ;
  assign n30 = n29 ^ n13 ;
  assign n31 = n30 ^ n14 ;
  assign y0 = ~n31 ;
endmodule
