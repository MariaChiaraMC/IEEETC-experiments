module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n7 = x2 & x3 ;
  assign n8 = x1 & n7 ;
  assign n9 = n8 ^ x0 ;
  assign n19 = n9 ^ n8 ;
  assign n10 = x4 & x5 ;
  assign n11 = ~x3 & n10 ;
  assign n12 = n11 ^ n9 ;
  assign n13 = n12 ^ n8 ;
  assign n14 = ~x1 & ~x2 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = n15 ^ n11 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = ~n13 & ~n17 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = n20 ^ n13 ;
  assign n22 = x3 & ~x4 ;
  assign n23 = ~x5 & n22 ;
  assign n24 = n23 ^ n8 ;
  assign n25 = n18 ^ n13 ;
  assign n26 = n24 & ~n25 ;
  assign n27 = n26 ^ n8 ;
  assign n28 = ~n21 & ~n27 ;
  assign n29 = n28 ^ n8 ;
  assign n30 = n29 ^ x0 ;
  assign n31 = n30 ^ n8 ;
  assign y0 = n31 ;
endmodule
