// Benchmark "./pla/exep.pla_dbb_orig_62NonExact" written by ABC on Fri Nov 20 10:21:22 2020

module \./pla/exep.pla_dbb_orig_62NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = 1'b1;
endmodule


