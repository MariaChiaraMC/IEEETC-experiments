// Benchmark "./sqr6.pla" written by ABC on Thu Apr 23 11:00:04 2020

module \./sqr6.pla  ( 
    x0, x1, x2, x3, x4, x5,
    z9  );
  input  x0, x1, x2, x3, x4, x5;
  output z9;
  assign z9 = 1'b1;
endmodule


