// Benchmark "./pla/pope.rom.pla_dbb_orig_36NonExact" written by ABC on Fri Nov 20 10:28:00 2020

module \./pla/pope.rom.pla_dbb_orig_36NonExact  ( 
    x0, x1, x2, x3,
    z0  );
  input  x0, x1, x2, x3;
  output z0;
  wire new_n6_, new_n7_, new_n8_, new_n9_, new_n10_;
  assign new_n6_ = ~x0 & x1;
  assign new_n7_ = ~x1 & ~x2;
  assign new_n8_ = x3 & new_n7_;
  assign new_n9_ = ~x3 & ~new_n7_;
  assign new_n10_ = ~new_n8_ & ~new_n9_;
  assign z0 = ~new_n6_ & ~new_n10_;
endmodule


