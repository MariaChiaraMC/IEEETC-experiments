module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n11 = ~x2 & ~x4 ;
  assign n12 = ~x0 & ~x1 ;
  assign n13 = ~x3 & n12 ;
  assign n14 = n11 & n13 ;
  assign n15 = x7 ^ x6 ;
  assign n16 = n15 ^ x5 ;
  assign n17 = n14 & ~n16 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = x9 ^ x8 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n15 & n20 ;
  assign n22 = n21 ^ n15 ;
  assign n23 = n22 ^ x5 ;
  assign n24 = n18 & ~n23 ;
  assign y0 = n24 ;
endmodule
