module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 ;
  assign n16 = ~x8 & ~x11 ;
  assign n17 = ~x0 & n16 ;
  assign n18 = ~x13 & n17 ;
  assign n26 = x9 & x10 ;
  assign n27 = ~x6 & n26 ;
  assign n23 = x4 & x5 ;
  assign n28 = x2 & n23 ;
  assign n29 = ~x3 & x12 ;
  assign n30 = n28 & n29 ;
  assign n31 = n27 & n30 ;
  assign n32 = x14 & n31 ;
  assign n33 = ~x2 & ~x14 ;
  assign n34 = x9 ^ x4 ;
  assign n35 = n34 ^ x10 ;
  assign n36 = x3 & ~x6 ;
  assign n37 = n36 ^ x10 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = ~x3 & x6 ;
  assign n41 = n40 ^ x9 ;
  assign n42 = ~x9 & ~n41 ;
  assign n43 = n42 ^ n36 ;
  assign n44 = n43 ^ x9 ;
  assign n45 = n39 & ~n44 ;
  assign n46 = n45 ^ n42 ;
  assign n47 = n46 ^ x9 ;
  assign n48 = n35 & ~n47 ;
  assign n49 = x7 & n48 ;
  assign n50 = n33 & n49 ;
  assign n51 = n50 ^ x5 ;
  assign n52 = n51 ^ n50 ;
  assign n53 = n52 ^ x12 ;
  assign n54 = x7 & ~x9 ;
  assign n19 = ~x2 & ~x6 ;
  assign n55 = x10 & n19 ;
  assign n56 = n54 & n55 ;
  assign n57 = x2 & ~x14 ;
  assign n58 = x10 ^ x6 ;
  assign n59 = x10 ^ x9 ;
  assign n60 = n59 ^ x9 ;
  assign n61 = ~x7 & ~x9 ;
  assign n62 = n61 ^ x9 ;
  assign n63 = ~n60 & n62 ;
  assign n64 = n63 ^ x9 ;
  assign n65 = n58 & n64 ;
  assign n66 = n57 & n65 ;
  assign n67 = ~n56 & ~n66 ;
  assign n68 = ~x3 & x4 ;
  assign n69 = ~n67 & n68 ;
  assign n20 = ~x10 & x14 ;
  assign n21 = n19 & n20 ;
  assign n22 = x3 & n21 ;
  assign n70 = x9 ^ x7 ;
  assign n71 = ~x4 & n70 ;
  assign n72 = n22 & n71 ;
  assign n73 = n72 ^ n69 ;
  assign n74 = ~n69 & n73 ;
  assign n75 = n74 ^ n50 ;
  assign n76 = n75 ^ n69 ;
  assign n77 = ~n53 & n76 ;
  assign n78 = n77 ^ n74 ;
  assign n79 = n78 ^ n69 ;
  assign n80 = ~x12 & ~n79 ;
  assign n81 = n80 ^ x12 ;
  assign n82 = ~n32 & n81 ;
  assign n24 = ~x12 & n23 ;
  assign n25 = n22 & n24 ;
  assign n83 = n82 ^ n25 ;
  assign n84 = n83 ^ n82 ;
  assign n85 = n82 ^ n61 ;
  assign n86 = n85 ^ n82 ;
  assign n87 = n84 & n86 ;
  assign n88 = n87 ^ n82 ;
  assign n89 = x1 & ~n88 ;
  assign n90 = n89 ^ n82 ;
  assign n91 = n18 & ~n90 ;
  assign y0 = n91 ;
endmodule
