// Benchmark "./pla/x2dn.pla_res_19NonExact" written by ABC on Fri Nov 20 10:31:34 2020

module \./pla/x2dn.pla_res_19NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = x0;
endmodule


