module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 ;
  assign n15 = x2 & x13 ;
  assign n16 = ~x8 & n15 ;
  assign n17 = x4 & n16 ;
  assign n18 = x10 & ~n17 ;
  assign n19 = x13 ^ x0 ;
  assign n20 = x13 ^ x1 ;
  assign n21 = x13 ^ x8 ;
  assign n22 = x13 & n21 ;
  assign n23 = n22 ^ x13 ;
  assign n24 = ~n20 & n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n25 ^ x13 ;
  assign n27 = n26 ^ x8 ;
  assign n28 = ~n19 & n27 ;
  assign n29 = n18 & ~n28 ;
  assign n30 = x12 ^ x10 ;
  assign n31 = n30 ^ x10 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = ~x2 & ~x8 ;
  assign n34 = n33 ^ x3 ;
  assign n35 = n33 & ~n34 ;
  assign n36 = n35 ^ x10 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n32 & n37 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n39 ^ n33 ;
  assign n41 = ~n29 & n40 ;
  assign n42 = n41 ^ n29 ;
  assign n43 = ~x11 & n42 ;
  assign n44 = x10 & x12 ;
  assign n45 = ~x6 & x12 ;
  assign n46 = x11 & ~n45 ;
  assign n47 = ~x13 & n46 ;
  assign n48 = ~n44 & ~n47 ;
  assign n49 = n48 ^ x10 ;
  assign n50 = n49 ^ x8 ;
  assign n66 = n50 ^ n49 ;
  assign n52 = n15 ^ x8 ;
  assign n53 = n52 ^ n15 ;
  assign n54 = x5 & ~x6 ;
  assign n55 = x7 & n54 ;
  assign n56 = n55 ^ n15 ;
  assign n57 = n53 & ~n56 ;
  assign n58 = n57 ^ n15 ;
  assign n59 = x12 & n58 ;
  assign n60 = n59 ^ x8 ;
  assign n61 = x11 & n60 ;
  assign n51 = n50 ^ n48 ;
  assign n62 = n61 ^ n51 ;
  assign n63 = n61 ^ n50 ;
  assign n64 = n63 ^ n49 ;
  assign n65 = ~n62 & ~n64 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = ~x2 & ~x13 ;
  assign n69 = n68 ^ n50 ;
  assign n70 = n66 & n69 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = n67 & n71 ;
  assign n73 = n72 ^ n65 ;
  assign n74 = n73 ^ n50 ;
  assign n75 = n74 ^ x10 ;
  assign n76 = n75 ^ n49 ;
  assign n77 = ~n43 & n76 ;
  assign n78 = ~x9 & ~n77 ;
  assign n79 = x7 ^ x5 ;
  assign n80 = n79 ^ x7 ;
  assign n81 = x12 ^ x7 ;
  assign n82 = n80 & n81 ;
  assign n83 = n82 ^ x7 ;
  assign n84 = ~x6 & ~n83 ;
  assign n85 = n84 ^ x5 ;
  assign n86 = ~x4 & ~n85 ;
  assign n87 = ~x3 & ~n86 ;
  assign n88 = x4 & x5 ;
  assign n89 = x0 & ~n88 ;
  assign n90 = ~x10 & ~x11 ;
  assign n91 = x9 & n90 ;
  assign n92 = ~n89 & n91 ;
  assign n93 = x12 ^ x4 ;
  assign n94 = x6 ^ x4 ;
  assign n95 = n93 & ~n94 ;
  assign n96 = n95 ^ x4 ;
  assign n97 = x3 & ~n96 ;
  assign n98 = x13 & ~n97 ;
  assign n99 = n92 & ~n98 ;
  assign n100 = x8 & n99 ;
  assign n101 = ~n87 & n100 ;
  assign n102 = ~n78 & ~n101 ;
  assign y0 = ~n102 ;
endmodule
