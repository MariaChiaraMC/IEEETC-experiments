module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 ;
  output y0 ;
  wire n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 ;
  assign n25 = x3 & x5 ;
  assign n23 = ~x0 & x1 ;
  assign n24 = ~x2 & n23 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n26 ^ x4 ;
  assign n29 = x0 & ~x1 ;
  assign n28 = ~x3 & ~x5 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = n25 & ~n30 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = ~n27 & n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n34 ^ n28 ;
  assign n36 = n35 ^ n25 ;
  assign n37 = ~x4 & n36 ;
  assign n203 = ~x19 & ~x20 ;
  assign n38 = ~x12 & ~x13 ;
  assign n39 = ~x6 & ~x7 ;
  assign n40 = n39 ^ x9 ;
  assign n41 = ~x8 & n40 ;
  assign n42 = n41 ^ x9 ;
  assign n43 = ~x4 & n42 ;
  assign n44 = ~x8 & x9 ;
  assign n45 = x1 & ~x2 ;
  assign n46 = x10 & ~n45 ;
  assign n47 = ~n44 & ~n46 ;
  assign n48 = ~x11 & ~n47 ;
  assign n49 = x0 & x2 ;
  assign n50 = ~x5 & n49 ;
  assign n51 = n48 & n50 ;
  assign n52 = x1 & x2 ;
  assign n53 = ~x3 & ~n52 ;
  assign n54 = ~n51 & n53 ;
  assign n55 = n43 & ~n54 ;
  assign n61 = ~x0 & ~x2 ;
  assign n56 = ~x10 & x11 ;
  assign n57 = x8 & x9 ;
  assign n58 = n56 & n57 ;
  assign n59 = n39 & n58 ;
  assign n60 = n59 ^ n48 ;
  assign n62 = n61 ^ n60 ;
  assign n63 = n62 ^ n59 ;
  assign n71 = n63 ^ n60 ;
  assign n72 = n71 ^ n59 ;
  assign n73 = n72 ^ n59 ;
  assign n74 = x1 & x3 ;
  assign n75 = n74 ^ n60 ;
  assign n76 = n75 ^ n60 ;
  assign n77 = n76 ^ n59 ;
  assign n78 = n73 & ~n77 ;
  assign n64 = ~x1 & x9 ;
  assign n65 = ~x2 & n64 ;
  assign n66 = x3 & ~n65 ;
  assign n67 = n66 ^ n60 ;
  assign n68 = n67 ^ n63 ;
  assign n69 = n68 ^ n59 ;
  assign n70 = n63 & ~n69 ;
  assign n79 = n78 ^ n70 ;
  assign n80 = n79 ^ n63 ;
  assign n81 = n70 ^ n59 ;
  assign n82 = n81 ^ n72 ;
  assign n83 = ~n59 & n82 ;
  assign n84 = n83 ^ n70 ;
  assign n85 = n80 & n84 ;
  assign n86 = n85 ^ n78 ;
  assign n87 = n86 ^ n83 ;
  assign n88 = n87 ^ n63 ;
  assign n89 = n88 ^ n59 ;
  assign n90 = n89 ^ n72 ;
  assign n91 = n90 ^ n48 ;
  assign n92 = n55 & n91 ;
  assign n93 = n50 & n59 ;
  assign n94 = ~x1 & n93 ;
  assign n95 = ~n92 & ~n94 ;
  assign n96 = n38 & ~n95 ;
  assign n97 = x1 ^ x0 ;
  assign n98 = x2 & x4 ;
  assign n99 = n98 ^ x1 ;
  assign n100 = n99 ^ n98 ;
  assign n101 = x4 & ~n25 ;
  assign n102 = ~x8 & ~x10 ;
  assign n103 = x2 & ~x9 ;
  assign n104 = n28 & n103 ;
  assign n105 = n102 & n104 ;
  assign n106 = x11 & n105 ;
  assign n107 = ~n101 & ~n106 ;
  assign n108 = n107 ^ n98 ;
  assign n109 = ~n100 & ~n108 ;
  assign n110 = n109 ^ n98 ;
  assign n111 = n97 & n110 ;
  assign n112 = ~n96 & ~n111 ;
  assign n113 = ~x7 & n98 ;
  assign n114 = ~x3 & n113 ;
  assign n115 = x3 & ~x4 ;
  assign n116 = x9 & n115 ;
  assign n117 = n38 & n116 ;
  assign n118 = x10 & ~x11 ;
  assign n119 = n117 & n118 ;
  assign n120 = ~n114 & ~n119 ;
  assign n121 = x8 & ~n120 ;
  assign n122 = ~x12 & x13 ;
  assign n123 = ~x3 & ~n122 ;
  assign n124 = ~x1 & ~n123 ;
  assign n125 = ~n117 & ~n124 ;
  assign n126 = n125 ^ x1 ;
  assign n127 = ~x2 & ~n126 ;
  assign n128 = n127 ^ x1 ;
  assign n129 = ~x9 & ~x10 ;
  assign n130 = n129 ^ x11 ;
  assign n131 = ~x8 & n115 ;
  assign n132 = n131 ^ n130 ;
  assign n133 = ~x12 & n39 ;
  assign n134 = n133 ^ x13 ;
  assign n135 = n134 ^ n133 ;
  assign n136 = n133 ^ n129 ;
  assign n137 = n135 & n136 ;
  assign n138 = n137 ^ n133 ;
  assign n139 = n138 ^ n130 ;
  assign n140 = ~n132 & ~n139 ;
  assign n141 = n140 ^ n137 ;
  assign n142 = n141 ^ n133 ;
  assign n143 = n142 ^ n131 ;
  assign n144 = ~n130 & n143 ;
  assign n145 = n144 ^ n130 ;
  assign n146 = ~n128 & n145 ;
  assign n147 = ~n23 & ~n49 ;
  assign n148 = ~x4 & ~n147 ;
  assign n149 = ~x3 & ~n148 ;
  assign n150 = x13 ^ x1 ;
  assign n151 = n150 ^ x13 ;
  assign n152 = x11 & ~x12 ;
  assign n153 = n44 & n152 ;
  assign n154 = n153 ^ x13 ;
  assign n155 = ~n151 & ~n154 ;
  assign n156 = n155 ^ x13 ;
  assign n157 = ~n97 & n156 ;
  assign n158 = n157 ^ x0 ;
  assign n159 = x4 & n158 ;
  assign n160 = n56 ^ x2 ;
  assign n161 = n160 ^ n159 ;
  assign n175 = x13 & n102 ;
  assign n176 = ~n152 & ~n175 ;
  assign n177 = x9 & ~n176 ;
  assign n162 = ~x7 & x16 ;
  assign n163 = ~x9 & ~n162 ;
  assign n164 = ~x6 & ~x17 ;
  assign n165 = ~n163 & n164 ;
  assign n166 = x15 ^ x12 ;
  assign n167 = n166 ^ x12 ;
  assign n168 = x12 ^ x9 ;
  assign n169 = n168 ^ x12 ;
  assign n170 = ~n167 & ~n169 ;
  assign n171 = n170 ^ x12 ;
  assign n172 = x13 & ~n171 ;
  assign n173 = n172 ^ x12 ;
  assign n174 = n165 & ~n173 ;
  assign n178 = n177 ^ n174 ;
  assign n179 = n56 & n178 ;
  assign n180 = n179 ^ n177 ;
  assign n181 = ~n161 & ~n180 ;
  assign n182 = n181 ^ n179 ;
  assign n183 = n182 ^ n177 ;
  assign n184 = n183 ^ n56 ;
  assign n185 = n159 & ~n184 ;
  assign n186 = n149 & ~n185 ;
  assign n187 = n146 & ~n186 ;
  assign n188 = ~n121 & n187 ;
  assign n189 = n188 ^ x5 ;
  assign n190 = n189 ^ n188 ;
  assign n191 = n190 ^ n112 ;
  assign n192 = x2 & x21 ;
  assign n193 = x4 & ~n192 ;
  assign n194 = n193 ^ n74 ;
  assign n195 = n74 & n194 ;
  assign n196 = n195 ^ n188 ;
  assign n197 = n196 ^ n74 ;
  assign n198 = ~n191 & ~n197 ;
  assign n199 = n198 ^ n195 ;
  assign n200 = n199 ^ n74 ;
  assign n201 = n112 & n200 ;
  assign n202 = n201 ^ n112 ;
  assign n204 = n203 ^ n202 ;
  assign n205 = n204 ^ n202 ;
  assign n206 = n202 ^ x18 ;
  assign n207 = ~n205 & n206 ;
  assign n208 = n207 ^ n202 ;
  assign n209 = ~n37 & n208 ;
  assign n210 = x14 & ~n209 ;
  assign y0 = n210 ;
endmodule
