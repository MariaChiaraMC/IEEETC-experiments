module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 ;
  output y0 ;
  wire n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 ;
  assign n23 = ~x0 & x1 ;
  assign n24 = n23 ^ x2 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ x4 ;
  assign n28 = x0 & ~x1 ;
  assign n29 = n28 ^ x5 ;
  assign n27 = n23 ^ x5 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n30 ^ n25 ;
  assign n32 = n26 & n31 ;
  assign n33 = n32 ^ n27 ;
  assign n34 = n33 ^ n25 ;
  assign n37 = x4 & x5 ;
  assign n35 = x5 ^ x3 ;
  assign n36 = n35 ^ x5 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = n38 ^ x5 ;
  assign n40 = n39 ^ x4 ;
  assign n41 = n29 ^ n25 ;
  assign n42 = n36 ^ n28 ;
  assign n43 = n42 ^ x5 ;
  assign n44 = n41 & ~n43 ;
  assign n45 = n44 ^ n25 ;
  assign n46 = ~n40 & n45 ;
  assign n47 = n46 ^ n36 ;
  assign n48 = n47 ^ x4 ;
  assign n49 = n34 & ~n48 ;
  assign n50 = n49 ^ n37 ;
  assign n51 = n50 ^ x5 ;
  assign n52 = ~x19 & ~x20 ;
  assign n53 = n52 ^ x18 ;
  assign n54 = n53 ^ x18 ;
  assign n55 = ~x12 & ~x13 ;
  assign n56 = x5 & x9 ;
  assign n57 = ~x2 & n56 ;
  assign n58 = ~x10 & x11 ;
  assign n59 = x8 & n58 ;
  assign n60 = ~x6 & ~x7 ;
  assign n61 = ~x1 & n60 ;
  assign n62 = n59 & n61 ;
  assign n63 = ~x1 & ~x2 ;
  assign n64 = ~x5 & ~n63 ;
  assign n65 = n60 ^ x10 ;
  assign n66 = ~x8 & n65 ;
  assign n67 = n66 ^ x10 ;
  assign n68 = ~n64 & n67 ;
  assign n69 = ~x11 & n68 ;
  assign n70 = ~n62 & ~n69 ;
  assign n71 = x9 & ~n70 ;
  assign n72 = x3 & n71 ;
  assign n73 = ~x8 & ~x11 ;
  assign n74 = ~n59 & ~n73 ;
  assign n75 = n60 & ~n74 ;
  assign n78 = ~x0 & ~x2 ;
  assign n76 = ~x1 & x10 ;
  assign n77 = n73 & n76 ;
  assign n79 = n78 ^ n77 ;
  assign n80 = n79 ^ n75 ;
  assign n81 = x9 ^ x5 ;
  assign n82 = n78 & ~n81 ;
  assign n83 = n82 ^ x5 ;
  assign n84 = n80 & n83 ;
  assign n85 = n84 ^ n82 ;
  assign n86 = n85 ^ x5 ;
  assign n87 = n86 ^ n78 ;
  assign n88 = n75 & n87 ;
  assign n89 = ~n72 & ~n88 ;
  assign n90 = ~n57 & n89 ;
  assign n91 = n55 & ~n90 ;
  assign n92 = x3 & x5 ;
  assign n93 = ~x8 & ~x9 ;
  assign n94 = n58 & n93 ;
  assign n95 = x13 & n94 ;
  assign n96 = ~x8 & n60 ;
  assign n97 = ~x9 & n96 ;
  assign n98 = n58 & n97 ;
  assign n99 = ~x12 & n98 ;
  assign n100 = n99 ^ n92 ;
  assign n101 = n95 & n100 ;
  assign n102 = n101 ^ n99 ;
  assign n103 = n92 & n102 ;
  assign n104 = ~n91 & ~n103 ;
  assign n105 = ~x4 & ~n104 ;
  assign n106 = ~x0 & ~x1 ;
  assign n107 = ~x5 & ~n106 ;
  assign n108 = n107 ^ x4 ;
  assign n109 = x2 & n55 ;
  assign n110 = x9 & ~x10 ;
  assign n111 = x8 & n110 ;
  assign n112 = n109 & n111 ;
  assign n113 = x11 & n28 ;
  assign n114 = n112 & n113 ;
  assign n115 = n60 & n114 ;
  assign n116 = n115 ^ n108 ;
  assign n117 = n116 ^ n107 ;
  assign n118 = n117 ^ n116 ;
  assign n119 = x1 & x2 ;
  assign n120 = x0 & ~x5 ;
  assign n121 = n119 & ~n120 ;
  assign n122 = n121 ^ n116 ;
  assign n123 = n122 ^ n108 ;
  assign n124 = n118 & ~n123 ;
  assign n125 = n124 ^ n121 ;
  assign n126 = ~x3 & ~n121 ;
  assign n127 = n126 ^ n108 ;
  assign n128 = ~n125 & ~n127 ;
  assign n129 = n128 ^ n126 ;
  assign n130 = ~n108 & n129 ;
  assign n131 = n130 ^ n124 ;
  assign n132 = n131 ^ x4 ;
  assign n133 = n132 ^ n121 ;
  assign n134 = x13 & n37 ;
  assign n135 = ~x4 & n96 ;
  assign n136 = ~x11 & n55 ;
  assign n137 = n110 & n136 ;
  assign n138 = n135 & n137 ;
  assign n141 = n138 ^ x0 ;
  assign n158 = n141 ^ n138 ;
  assign n159 = n158 ^ n138 ;
  assign n160 = ~n158 & ~n159 ;
  assign n143 = x10 & ~x11 ;
  assign n144 = n96 ^ x8 ;
  assign n145 = ~x9 & n144 ;
  assign n146 = n145 ^ x8 ;
  assign n147 = n143 & n146 ;
  assign n148 = ~x0 & ~n59 ;
  assign n149 = x9 & n75 ;
  assign n150 = ~n148 & n149 ;
  assign n151 = ~n147 & ~n150 ;
  assign n139 = ~x4 & n109 ;
  assign n140 = n139 ^ n138 ;
  assign n142 = n141 ^ n140 ;
  assign n152 = n151 ^ n142 ;
  assign n153 = n152 ^ n142 ;
  assign n154 = n142 ^ n141 ;
  assign n155 = n154 ^ n138 ;
  assign n156 = ~n153 & n155 ;
  assign n163 = n160 ^ n156 ;
  assign n157 = n156 ^ x5 ;
  assign n161 = n160 ^ n158 ;
  assign n162 = n157 & ~n161 ;
  assign n164 = n163 ^ n162 ;
  assign n165 = x5 & n164 ;
  assign n166 = n165 ^ n156 ;
  assign n167 = n166 ^ n160 ;
  assign n168 = n167 ^ n162 ;
  assign n169 = n168 ^ x0 ;
  assign n170 = ~n134 & n169 ;
  assign n171 = x1 & ~n170 ;
  assign n172 = x9 & n96 ;
  assign n173 = n172 ^ n146 ;
  assign n174 = ~x10 & n173 ;
  assign n175 = n174 ^ n146 ;
  assign n176 = n136 & n175 ;
  assign n177 = ~n94 & ~n176 ;
  assign n178 = n28 & ~n177 ;
  assign n179 = x12 & ~x13 ;
  assign n180 = ~x17 & ~n179 ;
  assign n181 = n98 & n180 ;
  assign n182 = x16 & n181 ;
  assign n183 = n37 & ~n182 ;
  assign n184 = ~n178 & ~n183 ;
  assign n185 = x2 & ~n184 ;
  assign n186 = n73 & n110 ;
  assign n187 = x12 & ~n186 ;
  assign n188 = ~x2 & x13 ;
  assign n189 = ~n187 & n188 ;
  assign n190 = ~x1 & x9 ;
  assign n191 = x11 & ~x12 ;
  assign n192 = ~x8 & n191 ;
  assign n193 = n190 & n192 ;
  assign n194 = x4 & ~n193 ;
  assign n195 = ~n189 & n194 ;
  assign n196 = ~x21 & n119 ;
  assign n197 = x5 & ~n196 ;
  assign n198 = ~n195 & n197 ;
  assign n199 = x2 & n134 ;
  assign n200 = x17 & n143 ;
  assign n201 = n23 & n55 ;
  assign n202 = n135 & n201 ;
  assign n203 = n200 & n202 ;
  assign n204 = ~n199 & ~n203 ;
  assign n205 = x15 & ~n204 ;
  assign n206 = n56 & n191 ;
  assign n207 = x10 & n206 ;
  assign n208 = n207 ^ n78 ;
  assign n209 = n208 ^ n78 ;
  assign n210 = n78 ^ n28 ;
  assign n211 = n210 ^ n78 ;
  assign n212 = ~n209 & ~n211 ;
  assign n213 = n212 ^ n78 ;
  assign n214 = x4 & ~n213 ;
  assign n215 = n214 ^ n78 ;
  assign n216 = ~n205 & ~n215 ;
  assign n217 = ~n198 & n216 ;
  assign n218 = ~n185 & n217 ;
  assign n219 = ~n171 & n218 ;
  assign n220 = n219 ^ x3 ;
  assign n221 = n220 ^ n219 ;
  assign n222 = n221 ^ n133 ;
  assign n223 = ~n63 & ~n119 ;
  assign n224 = n223 ^ x5 ;
  assign n225 = ~n223 & ~n224 ;
  assign n226 = n225 ^ n219 ;
  assign n227 = n226 ^ n223 ;
  assign n228 = n222 & n227 ;
  assign n229 = n228 ^ n225 ;
  assign n230 = n229 ^ n223 ;
  assign n231 = n133 & ~n230 ;
  assign n232 = n231 ^ n133 ;
  assign n233 = ~n105 & n232 ;
  assign n234 = n233 ^ x18 ;
  assign n235 = n54 & n234 ;
  assign n236 = n235 ^ x18 ;
  assign n237 = x14 & n236 ;
  assign n238 = ~n51 & n237 ;
  assign y0 = ~n238 ;
endmodule
