module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n12 = x9 ^ x5 ;
  assign n13 = n12 ^ x10 ;
  assign n14 = n13 ^ x1 ;
  assign n15 = x6 & ~x7 ;
  assign n16 = n15 ^ x5 ;
  assign n17 = ~x10 & ~n16 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n14 & n18 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n20 ^ n15 ;
  assign n22 = n21 ^ x10 ;
  assign n23 = ~x1 & ~n22 ;
  assign n24 = ~x3 & n23 ;
  assign n25 = ~x0 & ~n24 ;
  assign n26 = ~x2 & x4 ;
  assign n27 = x8 ^ x0 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = x7 ^ x6 ;
  assign n30 = ~x8 & n29 ;
  assign n31 = n30 ^ x6 ;
  assign n32 = n28 & ~n31 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ x6 ;
  assign n35 = n34 ^ x8 ;
  assign n36 = n26 & n35 ;
  assign n37 = ~n25 & n36 ;
  assign y0 = n37 ;
endmodule
