module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n8 = ~x4 & ~x5 ;
  assign n9 = x2 & ~n8 ;
  assign n10 = ~x0 & x3 ;
  assign n11 = ~n9 & n10 ;
  assign n12 = x2 ^ x1 ;
  assign n13 = n12 ^ x1 ;
  assign n14 = n13 ^ n11 ;
  assign n15 = x4 & x5 ;
  assign n16 = x6 ^ x1 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n15 & n17 ;
  assign n19 = n18 ^ x1 ;
  assign n20 = n19 ^ n15 ;
  assign n21 = ~n14 & n20 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = n22 ^ n15 ;
  assign n24 = n11 & n23 ;
  assign y0 = n24 ;
endmodule
