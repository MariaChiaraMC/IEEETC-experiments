module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 ;
  assign n15 = x8 ^ x5 ;
  assign n11 = x8 ^ x7 ;
  assign n12 = n11 ^ x3 ;
  assign n13 = n12 ^ n11 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = n16 ^ n11 ;
  assign n14 = n13 ^ n11 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = x4 & ~n18 ;
  assign n20 = n19 ^ n13 ;
  assign n21 = n20 ^ n14 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = n11 ^ x8 ;
  assign n24 = n23 ^ x4 ;
  assign n25 = n24 ^ n13 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = n13 & n26 ;
  assign n28 = n27 ^ n14 ;
  assign n29 = x6 & ~n14 ;
  assign n30 = n29 ^ x6 ;
  assign n31 = n30 ^ n24 ;
  assign n32 = n31 ^ x4 ;
  assign n33 = ~n28 & n32 ;
  assign n34 = n33 ^ n13 ;
  assign n35 = n34 ^ n24 ;
  assign n36 = n35 ^ n14 ;
  assign n37 = n36 ^ x4 ;
  assign n38 = ~n22 & ~n37 ;
  assign n39 = n38 ^ n19 ;
  assign n40 = n39 ^ n33 ;
  assign n41 = n40 ^ n13 ;
  assign n42 = n41 ^ n24 ;
  assign n43 = n42 ^ n14 ;
  assign n44 = n43 ^ x8 ;
  assign n45 = ~x9 & n44 ;
  assign y0 = n45 ;
endmodule
