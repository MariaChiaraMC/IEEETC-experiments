module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 ;
  assign n19 = x8 & x9 ;
  assign n20 = ~x6 & n19 ;
  assign n21 = x6 ^ x1 ;
  assign n22 = n21 ^ x5 ;
  assign n28 = n22 ^ n21 ;
  assign n23 = n22 ^ x6 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = x9 ^ x6 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n24 & ~n26 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ n24 ;
  assign n31 = n21 ^ x8 ;
  assign n32 = n27 ^ n24 ;
  assign n33 = ~n31 & n32 ;
  assign n34 = n33 ^ n21 ;
  assign n35 = ~n30 & n34 ;
  assign n36 = n35 ^ n21 ;
  assign n37 = n36 ^ x1 ;
  assign n38 = n37 ^ n21 ;
  assign n39 = ~n20 & n38 ;
  assign n11 = ~x5 & x6 ;
  assign n12 = x1 & ~x8 ;
  assign n13 = ~x1 & x8 ;
  assign n14 = ~n12 & ~n13 ;
  assign n15 = ~x9 & n14 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = n11 & n16 ;
  assign n18 = ~x4 & ~n17 ;
  assign n40 = n39 ^ n18 ;
  assign n41 = ~x0 & ~n40 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = ~x2 & ~n42 ;
  assign n44 = x4 ^ x2 ;
  assign n45 = n44 ^ x3 ;
  assign n48 = ~x0 & ~x1 ;
  assign n51 = x5 & ~n48 ;
  assign n52 = x6 & ~n51 ;
  assign n53 = x1 & ~x6 ;
  assign n54 = ~x0 & x5 ;
  assign n55 = n54 ^ n19 ;
  assign n56 = n55 ^ n19 ;
  assign n57 = ~x8 & ~x9 ;
  assign n58 = ~x5 & ~x9 ;
  assign n59 = x0 & n58 ;
  assign n60 = ~n57 & ~n59 ;
  assign n61 = n60 ^ n19 ;
  assign n62 = ~n56 & ~n61 ;
  assign n63 = n62 ^ n19 ;
  assign n64 = n53 & n63 ;
  assign n65 = ~n52 & ~n64 ;
  assign n46 = ~x5 & ~n20 ;
  assign n47 = x5 & ~x6 ;
  assign n49 = ~n47 & n48 ;
  assign n50 = ~n46 & n49 ;
  assign n66 = n65 ^ n50 ;
  assign n67 = ~x2 & n66 ;
  assign n68 = n67 ^ n65 ;
  assign n69 = ~n45 & ~n68 ;
  assign n70 = n69 ^ n67 ;
  assign n71 = n70 ^ n65 ;
  assign n72 = n71 ^ x2 ;
  assign n73 = ~x3 & n72 ;
  assign n74 = ~n43 & n73 ;
  assign n75 = x1 ^ x0 ;
  assign n77 = n75 ^ x6 ;
  assign n84 = n77 ^ n75 ;
  assign n76 = n75 ^ x2 ;
  assign n78 = n77 ^ n76 ;
  assign n79 = n78 ^ x1 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = n78 ^ n77 ;
  assign n82 = n81 ^ n75 ;
  assign n83 = n80 & n82 ;
  assign n85 = n84 ^ n83 ;
  assign n86 = n19 ^ x8 ;
  assign n87 = n86 ^ n83 ;
  assign n88 = ~n75 & n87 ;
  assign n89 = n88 ^ x8 ;
  assign n90 = n89 ^ n75 ;
  assign n91 = ~n84 & n90 ;
  assign n92 = n91 ^ n75 ;
  assign n93 = ~n85 & ~n92 ;
  assign n94 = n93 ^ n91 ;
  assign n95 = n94 ^ x6 ;
  assign n96 = n95 ^ n75 ;
  assign n97 = x5 & ~n96 ;
  assign n98 = ~x1 & ~x2 ;
  assign n99 = n20 & n98 ;
  assign n100 = x3 & ~n99 ;
  assign n101 = x0 & x2 ;
  assign n102 = n58 & n101 ;
  assign n103 = x8 ^ x1 ;
  assign n104 = n102 & n103 ;
  assign n105 = n100 & ~n104 ;
  assign n106 = ~n97 & n105 ;
  assign n107 = n106 ^ x6 ;
  assign n108 = n107 ^ n106 ;
  assign n109 = x1 & n101 ;
  assign n110 = n109 ^ n106 ;
  assign n111 = n110 ^ n106 ;
  assign n112 = n111 ^ x4 ;
  assign n113 = n108 & ~n112 ;
  assign n114 = n113 ^ n108 ;
  assign n115 = n114 ^ x4 ;
  assign n116 = n106 ^ x5 ;
  assign n117 = n116 ^ n111 ;
  assign n118 = n106 ^ x9 ;
  assign n119 = n117 & ~n118 ;
  assign n120 = n119 ^ x9 ;
  assign n121 = n120 ^ n106 ;
  assign n122 = n121 ^ n111 ;
  assign n123 = n122 ^ n116 ;
  assign n124 = n123 ^ x4 ;
  assign n125 = n111 ^ n106 ;
  assign n126 = ~x4 & n125 ;
  assign n127 = n126 ^ n111 ;
  assign n128 = n127 ^ n116 ;
  assign n129 = n128 ^ x4 ;
  assign n130 = n124 & ~n129 ;
  assign n131 = n130 ^ n116 ;
  assign n132 = ~n115 & n131 ;
  assign n133 = n132 ^ n126 ;
  assign n134 = n133 ^ n130 ;
  assign n135 = n134 ^ n111 ;
  assign n136 = n135 ^ n116 ;
  assign n137 = n136 ^ x4 ;
  assign n138 = n137 ^ x4 ;
  assign n139 = ~n74 & ~n138 ;
  assign n140 = ~x7 & ~n139 ;
  assign y0 = n140 ;
endmodule
