module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 ;
  assign n38 = x3 & x4 ;
  assign n39 = ~x2 & n38 ;
  assign n40 = x2 & ~x3 ;
  assign n42 = n40 ^ x4 ;
  assign n41 = n40 ^ x0 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = n43 ^ x3 ;
  assign n45 = n44 ^ n43 ;
  assign n46 = n45 ^ n40 ;
  assign n47 = n43 ^ n41 ;
  assign n48 = n47 ^ n40 ;
  assign n49 = n48 ^ n41 ;
  assign n50 = n49 ^ n40 ;
  assign n51 = n50 ^ n48 ;
  assign n52 = n46 & n51 ;
  assign n53 = n52 ^ n45 ;
  assign n54 = n43 ^ x5 ;
  assign n55 = n54 ^ n44 ;
  assign n56 = n43 ^ x6 ;
  assign n57 = n56 ^ n44 ;
  assign n58 = n55 & n57 ;
  assign n59 = n58 ^ n45 ;
  assign n60 = n53 ^ n48 ;
  assign n61 = n59 & ~n60 ;
  assign n62 = n61 ^ n50 ;
  assign n63 = n62 ^ n48 ;
  assign n64 = n53 & n63 ;
  assign n65 = n64 ^ n45 ;
  assign n66 = n65 ^ n46 ;
  assign n67 = n66 ^ x0 ;
  assign n68 = n67 ^ n40 ;
  assign n69 = ~n39 & n68 ;
  assign n11 = x3 ^ x0 ;
  assign n8 = ~x5 & ~x6 ;
  assign n9 = ~x4 & n8 ;
  assign n12 = n11 ^ n9 ;
  assign n10 = n9 ^ x3 ;
  assign n17 = n12 ^ n10 ;
  assign n18 = n17 ^ x2 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = ~x3 & ~x4 ;
  assign n21 = ~x5 & n20 ;
  assign n22 = n21 ^ n12 ;
  assign n23 = n22 ^ x2 ;
  assign n24 = ~n19 & ~n23 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = n13 ^ n10 ;
  assign n15 = n14 ^ x2 ;
  assign n16 = n10 & ~n15 ;
  assign n25 = n24 ^ n16 ;
  assign n26 = n25 ^ n10 ;
  assign n27 = n16 ^ x2 ;
  assign n28 = n27 ^ n18 ;
  assign n29 = ~x2 & ~n28 ;
  assign n30 = n29 ^ n16 ;
  assign n31 = n26 & n30 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ n10 ;
  assign n35 = n34 ^ x2 ;
  assign n36 = n35 ^ n18 ;
  assign n37 = n36 ^ x0 ;
  assign n70 = n69 ^ n37 ;
  assign n71 = ~x1 & n70 ;
  assign n72 = n71 ^ n37 ;
  assign y0 = ~n72 ;
endmodule
