module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 ;
  assign n17 = ~x0 & ~x4 ;
  assign n18 = ~x3 & n17 ;
  assign n19 = ~x1 & ~x2 ;
  assign n20 = n18 & n19 ;
  assign n21 = x6 & n20 ;
  assign n22 = x9 ^ x8 ;
  assign n23 = x7 & n22 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = ~x10 & ~x11 ;
  assign n28 = n27 ^ x7 ;
  assign n29 = ~n27 & ~n28 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n26 & n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = n21 & ~n34 ;
  assign n36 = n35 ^ n21 ;
  assign y0 = n36 ;
endmodule
