module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n9 = ~x1 & x3 ;
  assign n10 = ~x5 & ~n9 ;
  assign n11 = ~x4 & ~n10 ;
  assign n12 = ~x6 & ~n11 ;
  assign n13 = ~x0 & x7 ;
  assign n14 = x5 ^ x1 ;
  assign n15 = n14 ^ x6 ;
  assign n16 = x3 ^ x2 ;
  assign n17 = x6 ^ x5 ;
  assign n18 = x4 ^ x3 ;
  assign n19 = n18 ^ x3 ;
  assign n20 = ~n17 & ~n19 ;
  assign n21 = n20 ^ x3 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = ~n16 & n22 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n15 & ~n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = x6 & n26 ;
  assign n28 = n27 ^ x6 ;
  assign n29 = n13 & ~n28 ;
  assign n30 = ~n12 & n29 ;
  assign y0 = n30 ;
endmodule
