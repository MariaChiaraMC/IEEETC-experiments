module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n7 = ~x2 & ~x3 ;
  assign n8 = x4 & x5 ;
  assign n9 = ~x3 & ~n8 ;
  assign n10 = x0 & ~n9 ;
  assign n11 = ~n7 & ~n10 ;
  assign n12 = x1 & ~n11 ;
  assign n13 = n8 ^ x0 ;
  assign n14 = n13 ^ n7 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = ~x2 & ~x5 ;
  assign n18 = x3 & ~n17 ;
  assign n19 = ~x4 & ~n18 ;
  assign n20 = ~x1 & ~n19 ;
  assign n21 = n20 ^ x0 ;
  assign n22 = ~x0 & ~n21 ;
  assign n23 = n22 ^ n13 ;
  assign n24 = n23 ^ x0 ;
  assign n25 = n16 & n24 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = n26 ^ x0 ;
  assign n28 = ~n12 & ~n27 ;
  assign n29 = n28 ^ n12 ;
  assign y0 = n29 ;
endmodule
