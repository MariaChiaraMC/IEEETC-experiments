module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 ;
  assign n13 = ~x8 & x11 ;
  assign n14 = x4 & x5 ;
  assign n15 = x1 & n14 ;
  assign n16 = n13 & n15 ;
  assign n17 = ~x3 & ~x5 ;
  assign n18 = x4 & n17 ;
  assign n19 = x8 & x10 ;
  assign n20 = ~x9 & n19 ;
  assign n21 = n18 & n20 ;
  assign n22 = ~x5 & x10 ;
  assign n23 = ~x3 & ~x9 ;
  assign n24 = x1 & n23 ;
  assign n25 = n22 & n24 ;
  assign n26 = ~n21 & ~n25 ;
  assign n27 = ~x4 & x9 ;
  assign n28 = ~x1 & ~n27 ;
  assign n29 = x5 & x11 ;
  assign n30 = x3 & ~x8 ;
  assign n31 = n29 & n30 ;
  assign n32 = ~n28 & n31 ;
  assign n33 = n26 & ~n32 ;
  assign n34 = x0 & ~n33 ;
  assign n35 = x3 & x4 ;
  assign n36 = ~x5 & n35 ;
  assign n37 = n20 & n36 ;
  assign n38 = ~x3 & x5 ;
  assign n39 = n13 & n38 ;
  assign n40 = n27 & n39 ;
  assign n41 = ~n37 & ~n40 ;
  assign n42 = ~x6 & ~n41 ;
  assign n43 = x1 & ~x4 ;
  assign n44 = ~x5 & ~x9 ;
  assign n45 = n43 & n44 ;
  assign n46 = x10 & n45 ;
  assign n47 = ~n42 & ~n46 ;
  assign n48 = ~n34 & n47 ;
  assign n49 = ~n16 & n48 ;
  assign n50 = ~x5 & x9 ;
  assign n51 = ~x10 & n50 ;
  assign n52 = ~x4 & n51 ;
  assign n53 = n30 & n52 ;
  assign n54 = x8 & ~x11 ;
  assign n55 = n14 & n54 ;
  assign n56 = n23 & n55 ;
  assign n57 = ~x6 & ~n56 ;
  assign n58 = ~n53 & n57 ;
  assign n59 = x5 & x8 ;
  assign n60 = n59 ^ x10 ;
  assign n61 = n59 ^ n50 ;
  assign n62 = n61 ^ n50 ;
  assign n63 = n50 ^ n35 ;
  assign n64 = n62 & ~n63 ;
  assign n65 = n64 ^ n50 ;
  assign n66 = ~n60 & ~n65 ;
  assign n67 = n66 ^ x10 ;
  assign n68 = ~x11 & ~n67 ;
  assign n69 = ~x3 & n51 ;
  assign n70 = n69 ^ x1 ;
  assign n71 = n69 ^ x4 ;
  assign n72 = n71 ^ x4 ;
  assign n73 = x3 & x5 ;
  assign n74 = n54 & n73 ;
  assign n75 = n74 ^ x4 ;
  assign n76 = ~n72 & n75 ;
  assign n77 = n76 ^ x4 ;
  assign n78 = ~n70 & ~n77 ;
  assign n79 = n78 ^ x1 ;
  assign n80 = ~n68 & n79 ;
  assign n81 = n80 ^ x0 ;
  assign n82 = n81 ^ n58 ;
  assign n83 = ~n52 & ~n55 ;
  assign n84 = n83 ^ x6 ;
  assign n85 = ~n80 & n84 ;
  assign n86 = n85 ^ n83 ;
  assign n87 = ~n82 & ~n86 ;
  assign n88 = n87 ^ n85 ;
  assign n89 = n88 ^ n83 ;
  assign n90 = n89 ^ n80 ;
  assign n91 = ~n58 & n90 ;
  assign n144 = ~x6 & ~n30 ;
  assign n175 = ~n23 & n144 ;
  assign n176 = x0 & ~x6 ;
  assign n177 = ~x10 & ~n176 ;
  assign n178 = ~x11 & n177 ;
  assign n179 = ~n175 & n178 ;
  assign n180 = ~x5 & ~x10 ;
  assign n92 = ~x1 & ~x4 ;
  assign n93 = ~x9 & n92 ;
  assign n107 = ~x1 & x4 ;
  assign n143 = ~x8 & n107 ;
  assign n181 = ~n93 & ~n143 ;
  assign n182 = ~x1 & x6 ;
  assign n94 = x1 & x4 ;
  assign n183 = n23 & ~n94 ;
  assign n184 = ~n182 & ~n183 ;
  assign n185 = ~x0 & ~n184 ;
  assign n186 = n181 & ~n185 ;
  assign n187 = n180 & ~n186 ;
  assign n188 = ~n179 & ~n187 ;
  assign n189 = x11 ^ x0 ;
  assign n190 = x6 & n35 ;
  assign n191 = n181 & ~n190 ;
  assign n192 = n191 ^ n189 ;
  assign n193 = n192 ^ x11 ;
  assign n194 = n193 ^ n192 ;
  assign n132 = x6 & ~x11 ;
  assign n195 = ~n24 & ~n132 ;
  assign n196 = x4 & ~n195 ;
  assign n197 = n196 ^ n192 ;
  assign n198 = n197 ^ n189 ;
  assign n199 = ~n194 & n198 ;
  assign n200 = n199 ^ n196 ;
  assign n201 = n30 & ~n43 ;
  assign n202 = ~n182 & ~n201 ;
  assign n203 = ~n196 & n202 ;
  assign n204 = n203 ^ n189 ;
  assign n205 = ~n200 & ~n204 ;
  assign n206 = n205 ^ n203 ;
  assign n207 = ~n189 & n206 ;
  assign n208 = n207 ^ n199 ;
  assign n209 = n208 ^ x0 ;
  assign n210 = n209 ^ n196 ;
  assign n211 = n210 ^ x5 ;
  assign n212 = n211 ^ n210 ;
  assign n95 = ~x3 & x6 ;
  assign n133 = ~n95 & ~n132 ;
  assign n145 = ~x0 & ~n144 ;
  assign n213 = n133 & ~n145 ;
  assign n214 = n43 & ~n213 ;
  assign n215 = n214 ^ n210 ;
  assign n216 = ~n212 & n215 ;
  assign n217 = n216 ^ n210 ;
  assign n218 = n188 & ~n217 ;
  assign n96 = ~x10 & n95 ;
  assign n97 = x1 & x10 ;
  assign n98 = ~x0 & ~n97 ;
  assign n99 = ~x6 & ~n23 ;
  assign n100 = n98 & ~n99 ;
  assign n101 = ~n96 & ~n100 ;
  assign n102 = ~n94 & ~n101 ;
  assign n103 = ~n93 & ~n102 ;
  assign n104 = n103 ^ x8 ;
  assign n105 = n104 ^ n103 ;
  assign n106 = n105 ^ x5 ;
  assign n108 = ~x6 & x9 ;
  assign n109 = ~n107 & n108 ;
  assign n110 = x10 & ~n28 ;
  assign n111 = x0 & n110 ;
  assign n112 = ~n109 & ~n111 ;
  assign n113 = ~x3 & ~n112 ;
  assign n114 = ~n97 & ~n108 ;
  assign n115 = ~n98 & ~n114 ;
  assign n116 = ~x4 & n115 ;
  assign n117 = n116 ^ n113 ;
  assign n118 = ~n113 & n117 ;
  assign n119 = n118 ^ n103 ;
  assign n120 = n119 ^ n113 ;
  assign n121 = ~n106 & ~n120 ;
  assign n122 = n121 ^ n118 ;
  assign n123 = n122 ^ n113 ;
  assign n124 = x5 & ~n123 ;
  assign n125 = n124 ^ x5 ;
  assign n126 = n125 ^ x5 ;
  assign n127 = x1 & x11 ;
  assign n128 = x4 & n127 ;
  assign n129 = ~x6 & x8 ;
  assign n130 = x3 & n129 ;
  assign n131 = ~n92 & n130 ;
  assign n134 = x4 & x8 ;
  assign n135 = x3 & n127 ;
  assign n136 = ~n134 & ~n135 ;
  assign n137 = x0 & ~n136 ;
  assign n138 = n133 & n137 ;
  assign n139 = ~n131 & ~n138 ;
  assign n140 = ~n128 & n139 ;
  assign n141 = n140 ^ x9 ;
  assign n142 = n141 ^ n140 ;
  assign n146 = n145 ^ x11 ;
  assign n147 = n146 ^ n43 ;
  assign n148 = x3 & x6 ;
  assign n149 = n148 ^ x1 ;
  assign n150 = n149 ^ n146 ;
  assign n151 = ~n145 & ~n150 ;
  assign n152 = n151 ^ x1 ;
  assign n153 = n152 ^ n145 ;
  assign n154 = n153 ^ n146 ;
  assign n155 = n154 ^ n43 ;
  assign n156 = n147 & ~n155 ;
  assign n157 = n156 ^ n151 ;
  assign n158 = n157 ^ x1 ;
  assign n159 = n158 ^ n146 ;
  assign n160 = ~n43 & ~n159 ;
  assign n161 = n160 ^ n43 ;
  assign n162 = n161 ^ n43 ;
  assign n163 = ~n143 & ~n162 ;
  assign n164 = n163 ^ n140 ;
  assign n165 = n142 & n164 ;
  assign n166 = n165 ^ n140 ;
  assign n167 = n166 ^ n125 ;
  assign n168 = n126 & n167 ;
  assign n169 = n168 ^ n165 ;
  assign n170 = n169 ^ n140 ;
  assign n171 = n170 ^ x5 ;
  assign n172 = ~n125 & n171 ;
  assign n173 = n172 ^ n125 ;
  assign n174 = n173 ^ n125 ;
  assign n219 = n218 ^ n174 ;
  assign n220 = ~x2 & n219 ;
  assign n221 = n220 ^ n218 ;
  assign n222 = ~n91 & n221 ;
  assign n223 = ~x7 & ~n222 ;
  assign n224 = n223 ^ n49 ;
  assign n225 = n17 & n97 ;
  assign n226 = n73 & n127 ;
  assign n227 = ~n225 & ~n226 ;
  assign n230 = x10 & n27 ;
  assign n228 = x11 & ~n180 ;
  assign n229 = ~n96 & n228 ;
  assign n231 = n230 ^ n229 ;
  assign n232 = n229 ^ n134 ;
  assign n233 = n232 ^ n134 ;
  assign n234 = ~x5 & ~n148 ;
  assign n235 = n234 ^ n134 ;
  assign n236 = ~n233 & ~n235 ;
  assign n237 = n236 ^ n134 ;
  assign n238 = n231 & n237 ;
  assign n239 = n238 ^ n230 ;
  assign n240 = n227 & ~n239 ;
  assign n241 = ~x7 & n182 ;
  assign n242 = x5 ^ x3 ;
  assign n243 = n241 & ~n242 ;
  assign n244 = n134 ^ n27 ;
  assign n245 = n27 ^ x3 ;
  assign n246 = n245 ^ n27 ;
  assign n247 = n246 ^ n243 ;
  assign n248 = n244 & ~n247 ;
  assign n249 = n248 ^ n134 ;
  assign n250 = n243 & n249 ;
  assign n251 = n240 & ~n250 ;
  assign n252 = x0 & ~n251 ;
  assign n253 = n17 & n109 ;
  assign n254 = ~n127 & ~n253 ;
  assign n255 = x10 & ~n254 ;
  assign n256 = x1 & n176 ;
  assign n257 = ~x7 & ~n256 ;
  assign n258 = x9 & n129 ;
  assign n259 = n257 & ~n258 ;
  assign n260 = n259 ^ n29 ;
  assign n261 = n259 ^ n22 ;
  assign n262 = n261 ^ n22 ;
  assign n263 = ~n94 & ~n131 ;
  assign n264 = n263 ^ n22 ;
  assign n265 = n262 & n264 ;
  assign n266 = n265 ^ n22 ;
  assign n267 = ~n260 & n266 ;
  assign n268 = n267 ^ n29 ;
  assign n269 = ~n255 & ~n268 ;
  assign n270 = ~n252 & n269 ;
  assign n271 = n270 ^ x2 ;
  assign n272 = n271 ^ n270 ;
  assign n273 = ~n50 & ~n59 ;
  assign n274 = ~n257 & n273 ;
  assign n275 = n274 ^ n270 ;
  assign n276 = ~n272 & ~n275 ;
  assign n277 = n276 ^ n270 ;
  assign n278 = n277 ^ n49 ;
  assign n279 = ~n224 & n278 ;
  assign n280 = n279 ^ n276 ;
  assign n281 = n280 ^ n270 ;
  assign n282 = n281 ^ n223 ;
  assign n283 = n49 & ~n282 ;
  assign n284 = n283 ^ n49 ;
  assign y0 = ~n284 ;
endmodule
