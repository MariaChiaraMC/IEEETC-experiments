module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 ;
  assign n17 = x9 & x10 ;
  assign n18 = x8 & n17 ;
  assign n12 = ~x9 & ~x10 ;
  assign n13 = ~x3 & x4 ;
  assign n14 = n12 & n13 ;
  assign n15 = x1 & x2 ;
  assign n16 = n14 & n15 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = n18 ^ x8 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = n20 & ~n22 ;
  assign n24 = n23 ^ n18 ;
  assign n25 = ~x6 & n24 ;
  assign n26 = n25 ^ n18 ;
  assign n27 = ~x5 & n26 ;
  assign n28 = n27 ^ x7 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = x6 ^ x5 ;
  assign n31 = n30 ^ x6 ;
  assign n32 = ~x6 & ~x8 ;
  assign n33 = ~n17 & n32 ;
  assign n34 = n33 ^ x6 ;
  assign n35 = n31 & n34 ;
  assign n36 = n35 ^ x6 ;
  assign n37 = ~n18 & n36 ;
  assign n38 = n37 ^ n27 ;
  assign n39 = n29 & n38 ;
  assign n40 = n39 ^ n27 ;
  assign n41 = ~x0 & n40 ;
  assign y0 = n41 ;
endmodule
