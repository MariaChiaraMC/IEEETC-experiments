// Benchmark "./pla/m3.pla_2" written by ABC on Mon Apr 20 15:44:08 2020

module \./pla/m3.pla_2  ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z0  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z0;
  assign z0 = ~x0;
endmodule


