module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 ;
  assign n7 = x1 ^ x0 ;
  assign n8 = ~x2 & x3 ;
  assign n9 = x2 & x4 ;
  assign n10 = ~x3 & n9 ;
  assign n11 = x5 & n10 ;
  assign n12 = ~n8 & ~n11 ;
  assign n13 = n12 ^ x1 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = ~x4 & x5 ;
  assign n16 = n8 & n15 ;
  assign n17 = ~n10 & ~n16 ;
  assign n18 = n17 ^ n12 ;
  assign n19 = ~n14 & n18 ;
  assign n20 = n19 ^ n12 ;
  assign n21 = ~n7 & ~n20 ;
  assign y0 = n21 ;
endmodule
