// Benchmark "./rd53.pla" written by ABC on Thu Apr 23 11:00:01 2020

module \./rd53.pla  ( 
    x0, x1, x2, x3, x4,
    z2  );
  input  x0, x1, x2, x3, x4;
  output z2;
  assign z2 = 1'b1;
endmodule


