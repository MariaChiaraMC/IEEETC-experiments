module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
  assign n9 = x4 ^ x3 ;
  assign n8 = x3 ^ x0 ;
  assign n10 = n9 ^ n8 ;
  assign n11 = n10 ^ n8 ;
  assign n15 = x3 ^ x2 ;
  assign n16 = n15 ^ n8 ;
  assign n17 = ~n8 & n16 ;
  assign n12 = x4 ^ x1 ;
  assign n13 = x3 & ~n12 ;
  assign n20 = n17 ^ n13 ;
  assign n14 = n13 ^ n11 ;
  assign n18 = n17 ^ n8 ;
  assign n19 = n14 & ~n18 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = n11 & n21 ;
  assign n23 = n22 ^ n17 ;
  assign n24 = n23 ^ n19 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = x6 & n25 ;
  assign n27 = n26 ^ x6 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = x3 & x4 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n30 ^ n26 ;
  assign n32 = n28 & ~n31 ;
  assign n33 = n32 ^ n26 ;
  assign n34 = x5 & ~n33 ;
  assign n35 = n34 ^ n26 ;
  assign y0 = ~n35 ;
endmodule
