module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n13 = x1 & x4 ;
  assign n14 = x0 & x9 ;
  assign n15 = x8 & ~x10 ;
  assign n16 = n14 & n15 ;
  assign n17 = n13 & n16 ;
  assign n18 = x7 & n17 ;
  assign n19 = ~x5 & ~x11 ;
  assign n20 = x6 & n19 ;
  assign n21 = ~x3 & n20 ;
  assign n22 = n21 ^ x2 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = x5 & ~x6 ;
  assign n25 = x11 & n24 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = ~n23 & n26 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = n18 & n28 ;
  assign y0 = n29 ;
endmodule
