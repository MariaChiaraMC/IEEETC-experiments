module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n8 = x2 & x6 ;
  assign n9 = ~x4 & x5 ;
  assign n10 = n8 & n9 ;
  assign n11 = x3 & n10 ;
  assign n12 = x1 & n11 ;
  assign n13 = x2 & ~x4 ;
  assign n14 = x1 & ~x6 ;
  assign n15 = n13 & ~n14 ;
  assign n16 = n15 ^ x5 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n17 ^ x3 ;
  assign n19 = ~x1 & ~n13 ;
  assign n20 = x4 & ~n8 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = ~n19 & n21 ;
  assign n23 = n22 ^ n15 ;
  assign n24 = n23 ^ n19 ;
  assign n25 = ~n18 & n24 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = n26 ^ n19 ;
  assign n28 = ~x3 & ~n27 ;
  assign n29 = n28 ^ x3 ;
  assign n30 = ~n12 & n29 ;
  assign n31 = ~x0 & ~n30 ;
  assign y0 = n31 ;
endmodule
