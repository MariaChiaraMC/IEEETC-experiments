// Benchmark "./m1.pla" written by ABC on Thu Apr 23 10:59:54 2020

module \./m1.pla  ( 
    x0, x1, x2, x3, x4, x5,
    z1  );
  input  x0, x1, x2, x3, x4, x5;
  output z1;
  assign z1 = 1'b1;
endmodule


