module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n7 = ~x4 & ~x5 ;
  assign n8 = x3 & ~n7 ;
  assign n9 = ~x2 & ~n8 ;
  assign n10 = x2 & x3 ;
  assign n11 = ~x1 & ~n10 ;
  assign n12 = ~n9 & n11 ;
  assign n13 = ~x0 & n12 ;
  assign n14 = x2 ^ x1 ;
  assign n15 = n14 ^ x1 ;
  assign n16 = n15 ^ x0 ;
  assign n17 = x5 ^ x1 ;
  assign n18 = x3 ^ x1 ;
  assign n19 = x4 ^ x1 ;
  assign n20 = n18 & n19 ;
  assign n21 = n20 ^ x0 ;
  assign n22 = n17 & ~n21 ;
  assign n23 = n22 ^ x1 ;
  assign n24 = n16 & n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = ~x0 & n25 ;
  assign n27 = n26 ^ n22 ;
  assign n28 = n27 ^ n24 ;
  assign n29 = ~n13 & ~n28 ;
  assign y0 = ~n29 ;
endmodule
