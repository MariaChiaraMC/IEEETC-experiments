module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ;
  assign n7 = x0 & x1 ;
  assign n8 = x4 ^ x2 ;
  assign n9 = n7 & ~n8 ;
  assign n10 = x3 & ~n9 ;
  assign n11 = x4 ^ x1 ;
  assign n12 = n11 ^ x3 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = ~n12 & n14 ;
  assign n16 = n15 ^ n11 ;
  assign n17 = ~x1 & ~x2 ;
  assign n18 = n17 ^ n12 ;
  assign n19 = x1 ^ x0 ;
  assign n20 = n19 ^ n11 ;
  assign n21 = n19 ^ n12 ;
  assign n22 = ~n20 & ~n21 ;
  assign n23 = n22 ^ x1 ;
  assign n24 = n23 ^ n12 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = ~n18 & n25 ;
  assign n27 = n26 ^ n12 ;
  assign n28 = n27 ^ x5 ;
  assign n29 = ~n16 & ~n28 ;
  assign n30 = n29 ^ n15 ;
  assign n31 = n30 ^ n11 ;
  assign n32 = ~n10 & ~n31 ;
  assign n33 = ~x0 & ~x1 ;
  assign n34 = x5 & n33 ;
  assign n35 = x2 & x4 ;
  assign n36 = x3 & ~n35 ;
  assign n37 = ~n8 & ~n36 ;
  assign n38 = n34 & n37 ;
  assign n39 = ~n32 & ~n38 ;
  assign y0 = ~n39 ;
endmodule
