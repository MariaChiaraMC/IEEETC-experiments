module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 ;
  assign n17 = x5 ^ x1 ;
  assign n18 = x7 ^ x5 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = ~x11 & ~x15 ;
  assign n21 = x14 & n20 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = ~x5 & n22 ;
  assign n24 = n23 ^ x4 ;
  assign n25 = ~n19 & n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n26 ^ x4 ;
  assign n28 = n27 ^ x5 ;
  assign n29 = n17 & ~n28 ;
  assign n30 = n29 ^ x1 ;
  assign n31 = ~x2 & n30 ;
  assign n32 = ~x0 & ~n31 ;
  assign n33 = x5 & ~n21 ;
  assign n34 = ~x12 & ~x13 ;
  assign n35 = ~x8 & n34 ;
  assign n36 = x10 ^ x9 ;
  assign n37 = n36 ^ x7 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = x10 ^ x6 ;
  assign n40 = ~x7 & ~n39 ;
  assign n41 = n40 ^ x6 ;
  assign n42 = ~n38 & n41 ;
  assign n43 = n42 ^ n40 ;
  assign n44 = n43 ^ x6 ;
  assign n45 = n44 ^ x7 ;
  assign n46 = n35 & ~n45 ;
  assign n47 = ~n33 & n46 ;
  assign n48 = x1 & ~n47 ;
  assign n49 = x6 ^ x0 ;
  assign n50 = n49 ^ x3 ;
  assign n51 = ~x4 & x5 ;
  assign n52 = n51 ^ x1 ;
  assign n53 = ~x0 & ~n52 ;
  assign n54 = n53 ^ x1 ;
  assign n55 = n50 & ~n54 ;
  assign n56 = n55 ^ n53 ;
  assign n57 = n56 ^ x1 ;
  assign n58 = n57 ^ x0 ;
  assign n59 = ~x3 & n58 ;
  assign n60 = ~n48 & n59 ;
  assign n61 = ~n32 & n60 ;
  assign y0 = n61 ;
endmodule
