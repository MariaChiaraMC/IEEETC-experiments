// Benchmark "./spla.pla" written by ABC on Thu Apr 23 11:00:01 2020

module \./spla.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15,
    z14  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15;
  output z14;
  assign z14 = 1'b1;
endmodule


