module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;
  assign n9 = x5 ^ x2 ;
  assign n8 = x3 ^ x1 ;
  assign n10 = n9 ^ n8 ;
  assign n11 = n10 ^ x5 ;
  assign n17 = n11 ^ x3 ;
  assign n12 = n9 ^ x5 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n11 ^ n9 ;
  assign n15 = n13 & n14 ;
  assign n16 = n15 ^ n9 ;
  assign n18 = n17 ^ n16 ;
  assign n20 = x4 ^ x2 ;
  assign n21 = n20 ^ x5 ;
  assign n22 = n21 ^ x3 ;
  assign n19 = n17 ^ n14 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = ~n17 & n23 ;
  assign n25 = n24 ^ n9 ;
  assign n26 = n25 ^ n11 ;
  assign n27 = n20 ^ x6 ;
  assign n28 = n27 ^ n20 ;
  assign n29 = n28 ^ n9 ;
  assign n30 = n29 ^ n11 ;
  assign n31 = n12 & n30 ;
  assign n32 = n31 ^ n9 ;
  assign n33 = n32 ^ n11 ;
  assign n34 = n33 ^ n17 ;
  assign n35 = n34 ^ n22 ;
  assign n36 = n26 & n35 ;
  assign n37 = n36 ^ n9 ;
  assign n38 = n37 ^ n12 ;
  assign n39 = n38 ^ n22 ;
  assign n40 = ~n18 & ~n39 ;
  assign n41 = n40 ^ n11 ;
  assign n42 = n41 ^ n17 ;
  assign n43 = ~x0 & ~n42 ;
  assign y0 = n43 ;
endmodule
