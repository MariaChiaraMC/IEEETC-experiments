module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n18 = x14 ^ x12 ;
  assign n19 = x13 & x15 ;
  assign n20 = x16 & n19 ;
  assign n21 = n20 ^ x14 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = ~x3 & ~x5 ;
  assign n24 = ~x2 & x4 ;
  assign n25 = n23 & n24 ;
  assign n26 = ~x15 & ~x16 ;
  assign n27 = x1 & ~x13 ;
  assign n28 = n26 & n27 ;
  assign n29 = n25 & n28 ;
  assign n30 = n29 ^ n20 ;
  assign n31 = ~n22 & n30 ;
  assign n32 = n31 ^ n20 ;
  assign n33 = ~n18 & n32 ;
  assign n34 = n33 ^ x12 ;
  assign y0 = n34 ;
endmodule
