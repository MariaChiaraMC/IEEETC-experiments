module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 ;
  assign n7 = x3 ^ x1 ;
  assign n8 = x5 ^ x3 ;
  assign n9 = x5 ^ x2 ;
  assign n10 = x5 & ~n9 ;
  assign n11 = n10 ^ x5 ;
  assign n12 = n8 & n11 ;
  assign n13 = n12 ^ n10 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = n14 ^ x2 ;
  assign n16 = n7 & ~n15 ;
  assign n17 = n16 ^ x1 ;
  assign n18 = x0 & ~n17 ;
  assign n25 = n9 ^ n8 ;
  assign n19 = n8 ^ x0 ;
  assign n20 = n19 ^ n9 ;
  assign n21 = n9 ^ x5 ;
  assign n22 = n21 ^ x0 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n20 & ~n23 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n26 ^ n20 ;
  assign n28 = n9 ^ x4 ;
  assign n29 = n24 ^ n20 ;
  assign n30 = n28 & n29 ;
  assign n31 = n30 ^ n9 ;
  assign n32 = ~n27 & n31 ;
  assign n33 = n32 ^ n9 ;
  assign n34 = n33 ^ n9 ;
  assign n35 = x1 & n34 ;
  assign n36 = ~n18 & ~n35 ;
  assign y0 = ~n36 ;
endmodule
