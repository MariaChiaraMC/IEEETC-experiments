module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 ;
  assign n16 = x10 & ~x13 ;
  assign n23 = x9 & n16 ;
  assign n24 = n23 ^ x14 ;
  assign n98 = n24 ^ x14 ;
  assign n99 = n98 ^ x14 ;
  assign n100 = n98 & ~n99 ;
  assign n26 = ~x4 & x5 ;
  assign n27 = x7 & ~x9 ;
  assign n28 = ~x0 & ~x1 ;
  assign n29 = n27 & n28 ;
  assign n30 = n26 & n29 ;
  assign n31 = x9 & x13 ;
  assign n32 = ~x1 & x7 ;
  assign n33 = x2 & ~x6 ;
  assign n34 = ~n32 & ~n33 ;
  assign n35 = x3 & ~n34 ;
  assign n36 = ~x6 & n28 ;
  assign n37 = ~x0 & ~x7 ;
  assign n38 = n37 ^ x3 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = x4 & x7 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n41 ^ n37 ;
  assign n43 = ~n39 & n42 ;
  assign n44 = n43 ^ n37 ;
  assign n45 = x2 & n44 ;
  assign n46 = n45 ^ n37 ;
  assign n47 = ~n36 & ~n46 ;
  assign n48 = ~n35 & n47 ;
  assign n49 = x5 & ~n48 ;
  assign n50 = ~x3 & ~n26 ;
  assign n52 = x5 & x7 ;
  assign n53 = x4 & ~n52 ;
  assign n51 = x2 & ~x5 ;
  assign n54 = n53 ^ n51 ;
  assign n55 = x6 & ~n54 ;
  assign n56 = n55 ^ n53 ;
  assign n57 = n50 & n56 ;
  assign n58 = x2 & ~x3 ;
  assign n59 = ~x0 & ~n58 ;
  assign n60 = ~x5 & n37 ;
  assign n61 = ~x4 & n60 ;
  assign n62 = ~n59 & ~n61 ;
  assign n63 = ~n57 & n62 ;
  assign n64 = x1 & ~n63 ;
  assign n65 = x4 & n51 ;
  assign n66 = ~n58 & ~n65 ;
  assign n67 = x0 & ~n66 ;
  assign n68 = ~x13 & ~n67 ;
  assign n69 = x3 & n26 ;
  assign n70 = ~x2 & n69 ;
  assign n71 = x9 ^ x0 ;
  assign n18 = ~x2 & ~x3 ;
  assign n72 = ~x4 & n18 ;
  assign n73 = n72 ^ x9 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = n74 ^ n71 ;
  assign n76 = x3 ^ x1 ;
  assign n77 = x3 & ~n76 ;
  assign n78 = n77 ^ n72 ;
  assign n79 = n78 ^ x3 ;
  assign n80 = ~n75 & n79 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n81 ^ x3 ;
  assign n83 = n71 & n82 ;
  assign n84 = n83 ^ x9 ;
  assign n85 = ~n70 & ~n84 ;
  assign n86 = n68 & n85 ;
  assign n87 = ~n64 & n86 ;
  assign n88 = ~n49 & n87 ;
  assign n89 = ~n31 & ~n88 ;
  assign n90 = ~x10 & ~n89 ;
  assign n91 = ~n30 & n90 ;
  assign n17 = x0 & ~x1 ;
  assign n19 = n17 & ~n18 ;
  assign n20 = x14 & ~n19 ;
  assign n21 = n16 & ~n20 ;
  assign n22 = n21 ^ x14 ;
  assign n25 = n24 ^ n22 ;
  assign n92 = n91 ^ n25 ;
  assign n93 = n92 ^ n25 ;
  assign n94 = n25 ^ n24 ;
  assign n95 = n94 ^ x14 ;
  assign n96 = ~n93 & ~n95 ;
  assign n103 = n100 ^ n96 ;
  assign n97 = n96 ^ x11 ;
  assign n101 = n100 ^ n98 ;
  assign n102 = n97 & n101 ;
  assign n104 = n103 ^ n102 ;
  assign n105 = x11 & n104 ;
  assign n106 = n105 ^ n96 ;
  assign n107 = n106 ^ n100 ;
  assign n108 = n107 ^ n102 ;
  assign n109 = n108 ^ n23 ;
  assign y0 = n109 ;
endmodule
