module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 ;
  assign n11 = ~x3 & ~x6 ;
  assign n12 = x5 & x8 ;
  assign n13 = ~x0 & x2 ;
  assign n14 = n12 & n13 ;
  assign n15 = n11 & n14 ;
  assign n16 = ~x5 & ~x8 ;
  assign n17 = ~x6 & n16 ;
  assign n18 = x3 & n17 ;
  assign n19 = n13 & n18 ;
  assign n20 = x3 & x6 ;
  assign n21 = ~n11 & ~n20 ;
  assign n22 = ~x0 & ~n21 ;
  assign n23 = ~x2 & n22 ;
  assign n24 = ~x5 & x8 ;
  assign n25 = n23 & n24 ;
  assign n26 = ~n19 & ~n25 ;
  assign n27 = ~n15 & n26 ;
  assign n28 = x1 & x4 ;
  assign n29 = ~n27 & n28 ;
  assign n30 = ~x0 & ~x6 ;
  assign n31 = ~x1 & ~x2 ;
  assign n32 = x5 & ~x8 ;
  assign n33 = n32 ^ n17 ;
  assign n34 = ~x0 & n33 ;
  assign n35 = n34 ^ n17 ;
  assign n36 = n31 & n35 ;
  assign n37 = ~n30 & n36 ;
  assign n38 = ~n29 & ~n37 ;
  assign n39 = n16 ^ n12 ;
  assign n40 = ~x6 & n39 ;
  assign n41 = n40 ^ n12 ;
  assign n42 = x3 ^ x0 ;
  assign n44 = n42 ^ x2 ;
  assign n50 = n44 ^ n42 ;
  assign n46 = x0 & n17 ;
  assign n43 = n42 ^ x3 ;
  assign n45 = n44 ^ n43 ;
  assign n47 = n46 ^ n45 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = n48 ^ n42 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = n45 ^ n44 ;
  assign n53 = n52 ^ n42 ;
  assign n54 = n53 ^ n42 ;
  assign n55 = n48 & ~n54 ;
  assign n56 = n55 ^ n48 ;
  assign n57 = ~n53 & n56 ;
  assign n58 = n57 ^ n42 ;
  assign n59 = n51 & n58 ;
  assign n60 = n59 ^ n55 ;
  assign n61 = n60 ^ n42 ;
  assign n62 = n61 ^ x2 ;
  assign n63 = n62 ^ n50 ;
  assign n64 = n41 & n63 ;
  assign n65 = ~n15 & ~n64 ;
  assign n66 = n65 ^ x1 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = x2 & n16 ;
  assign n69 = n68 ^ x8 ;
  assign n70 = x6 ^ x3 ;
  assign n71 = ~x2 & x5 ;
  assign n72 = n71 ^ x6 ;
  assign n73 = n70 & n72 ;
  assign n74 = ~x0 & n73 ;
  assign n75 = ~n69 & n74 ;
  assign n76 = n75 ^ n65 ;
  assign n77 = n67 & ~n76 ;
  assign n78 = n77 ^ n65 ;
  assign n79 = ~x4 & ~n78 ;
  assign n80 = n38 & ~n79 ;
  assign n81 = n80 ^ x7 ;
  assign n82 = n81 ^ n80 ;
  assign n83 = x8 ^ x5 ;
  assign n84 = x4 & n83 ;
  assign n85 = n84 ^ x5 ;
  assign n86 = n23 ^ n16 ;
  assign n87 = n86 ^ n23 ;
  assign n88 = x0 & x6 ;
  assign n89 = n88 ^ n23 ;
  assign n90 = n87 & n89 ;
  assign n91 = n90 ^ n23 ;
  assign n92 = ~n85 & n91 ;
  assign n93 = x1 & n92 ;
  assign n94 = x1 & ~x4 ;
  assign n95 = ~n21 & n94 ;
  assign n96 = ~x1 & x4 ;
  assign n97 = ~x3 & n96 ;
  assign n98 = x6 & n97 ;
  assign n99 = ~n95 & ~n98 ;
  assign n100 = n14 & ~n99 ;
  assign n101 = n20 & n96 ;
  assign n102 = x4 ^ x3 ;
  assign n103 = n102 ^ n88 ;
  assign n104 = n88 ^ x4 ;
  assign n105 = n104 ^ x4 ;
  assign n106 = n105 ^ n103 ;
  assign n107 = x4 ^ x1 ;
  assign n108 = n107 ^ n30 ;
  assign n109 = n30 & n108 ;
  assign n110 = n109 ^ x4 ;
  assign n111 = n110 ^ n30 ;
  assign n112 = ~n106 & ~n111 ;
  assign n113 = n112 ^ n109 ;
  assign n114 = n113 ^ n30 ;
  assign n115 = n103 & n114 ;
  assign n116 = n115 ^ n88 ;
  assign n117 = ~n101 & ~n116 ;
  assign n118 = n68 & ~n117 ;
  assign n119 = ~n100 & ~n118 ;
  assign n120 = ~n93 & n119 ;
  assign n121 = n120 ^ n80 ;
  assign n122 = ~n82 & n121 ;
  assign n123 = n122 ^ n80 ;
  assign n124 = ~x9 & ~n123 ;
  assign y0 = n124 ;
endmodule
