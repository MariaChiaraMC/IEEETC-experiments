module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 ;
  assign n10 = ~x1 & ~x2 ;
  assign n11 = x8 ^ x7 ;
  assign n12 = n10 & n11 ;
  assign n13 = ~x3 & n12 ;
  assign n14 = x0 & ~n13 ;
  assign n15 = ~x7 & ~x8 ;
  assign n16 = x4 ^ x1 ;
  assign n17 = ~x5 & ~x6 ;
  assign n18 = n17 ^ x4 ;
  assign n19 = ~n16 & ~n18 ;
  assign n20 = n19 ^ x4 ;
  assign n21 = n15 & n20 ;
  assign n22 = x3 & n21 ;
  assign n33 = x7 & ~x8 ;
  assign n23 = x8 ^ x4 ;
  assign n24 = x8 ^ x5 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = x5 & x6 ;
  assign n27 = n26 ^ x5 ;
  assign n28 = n25 & ~n27 ;
  assign n29 = n28 ^ x5 ;
  assign n30 = ~n23 & n29 ;
  assign n31 = n30 ^ x4 ;
  assign n32 = ~x3 & ~n31 ;
  assign n34 = n33 ^ n32 ;
  assign n35 = n34 ^ x1 ;
  assign n47 = n35 ^ n34 ;
  assign n36 = ~x1 & ~x7 ;
  assign n37 = x6 & ~x8 ;
  assign n38 = ~x4 & ~x5 ;
  assign n39 = ~n37 & n38 ;
  assign n40 = n36 & n39 ;
  assign n41 = n40 ^ n35 ;
  assign n42 = n41 ^ n34 ;
  assign n43 = n40 ^ n32 ;
  assign n44 = n43 ^ n40 ;
  assign n45 = n44 ^ n42 ;
  assign n46 = n42 & n45 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = n48 ^ n42 ;
  assign n50 = n34 ^ x7 ;
  assign n51 = n46 ^ n42 ;
  assign n52 = ~n50 & n51 ;
  assign n53 = n52 ^ n34 ;
  assign n54 = ~n49 & n53 ;
  assign n55 = n54 ^ n34 ;
  assign n56 = n55 ^ n32 ;
  assign n57 = n56 ^ n34 ;
  assign n58 = ~n22 & ~n57 ;
  assign n59 = ~x0 & ~x2 ;
  assign n60 = ~n58 & n59 ;
  assign n61 = ~x7 & x8 ;
  assign n62 = x2 & ~n61 ;
  assign n63 = ~x4 & ~n26 ;
  assign n64 = n36 & ~n63 ;
  assign n65 = n64 ^ x3 ;
  assign n66 = n65 ^ n64 ;
  assign n67 = n66 ^ n62 ;
  assign n68 = ~x8 & ~n17 ;
  assign n69 = x1 & ~x4 ;
  assign n70 = x8 & ~n26 ;
  assign n71 = ~n69 & ~n70 ;
  assign n72 = ~x1 & x4 ;
  assign n73 = ~n15 & ~n72 ;
  assign n74 = ~n71 & n73 ;
  assign n75 = n74 ^ n68 ;
  assign n76 = ~n68 & ~n75 ;
  assign n77 = n76 ^ n64 ;
  assign n78 = n77 ^ n68 ;
  assign n79 = ~n67 & ~n78 ;
  assign n80 = n79 ^ n76 ;
  assign n81 = n80 ^ n68 ;
  assign n82 = n62 & ~n81 ;
  assign n83 = n82 ^ n62 ;
  assign n84 = ~n60 & ~n83 ;
  assign n85 = x3 & x4 ;
  assign n86 = ~n17 & n85 ;
  assign n87 = n33 & n86 ;
  assign n88 = x1 & n87 ;
  assign n89 = ~n84 & ~n88 ;
  assign n90 = ~n14 & ~n89 ;
  assign y0 = n90 ;
endmodule
