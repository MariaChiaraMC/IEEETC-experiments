module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n11 = ~x3 & ~x6 ;
  assign n12 = ~x0 & ~x2 ;
  assign n13 = ~x8 & n12 ;
  assign n14 = ~n11 & ~n13 ;
  assign n15 = x9 ^ x8 ;
  assign n16 = x7 & ~n15 ;
  assign n17 = ~n14 & ~n16 ;
  assign n18 = x3 & x6 ;
  assign n19 = ~x1 & ~x5 ;
  assign n20 = ~n18 & n19 ;
  assign n21 = x2 ^ x0 ;
  assign n22 = n11 ^ x0 ;
  assign n23 = n11 ^ x4 ;
  assign n24 = ~n11 & n23 ;
  assign n25 = n24 ^ n11 ;
  assign n26 = n22 & ~n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n27 ^ n11 ;
  assign n29 = n28 ^ x4 ;
  assign n30 = ~n21 & n29 ;
  assign n31 = n30 ^ x4 ;
  assign n32 = n20 & ~n31 ;
  assign n33 = n17 & n32 ;
  assign y0 = n33 ;
endmodule
