module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 ;
  assign n10 = x7 & x8 ;
  assign n11 = ~x3 & n10 ;
  assign n12 = x2 & ~x4 ;
  assign n13 = ~x7 & n12 ;
  assign n14 = ~n11 & ~n13 ;
  assign n15 = x5 & x6 ;
  assign n16 = ~n14 & n15 ;
  assign n17 = ~x6 & ~x8 ;
  assign n18 = n17 ^ x4 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = ~x4 & ~x7 ;
  assign n21 = n20 ^ x4 ;
  assign n22 = n19 & n21 ;
  assign n23 = n22 ^ x4 ;
  assign n24 = x3 & n23 ;
  assign n25 = ~n10 & n24 ;
  assign n26 = n25 ^ x5 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = ~x6 & x7 ;
  assign n29 = ~x4 & ~x8 ;
  assign n30 = x6 & n29 ;
  assign n31 = ~n28 & ~n30 ;
  assign n32 = x3 & ~n31 ;
  assign n33 = x2 & x4 ;
  assign n34 = ~x6 & ~x7 ;
  assign n35 = n34 ^ x8 ;
  assign n36 = ~x3 & n35 ;
  assign n37 = n36 ^ x8 ;
  assign n38 = n33 & n37 ;
  assign n41 = ~x2 & n29 ;
  assign n42 = ~n10 & ~n41 ;
  assign n39 = ~x2 & x4 ;
  assign n40 = ~x8 & n39 ;
  assign n43 = n42 ^ n40 ;
  assign n44 = x6 & ~n43 ;
  assign n45 = n44 ^ n42 ;
  assign n46 = ~n38 & n45 ;
  assign n47 = ~n32 & n46 ;
  assign n48 = n47 ^ n25 ;
  assign n49 = ~n27 & ~n48 ;
  assign n50 = n49 ^ n25 ;
  assign n51 = ~n16 & ~n50 ;
  assign n52 = x1 & ~n51 ;
  assign n53 = x3 & x8 ;
  assign n56 = n15 & n53 ;
  assign n57 = ~x5 & ~x8 ;
  assign n58 = ~x4 & n57 ;
  assign n59 = ~n56 & ~n58 ;
  assign n54 = ~x5 & x6 ;
  assign n55 = n53 & n54 ;
  assign n60 = n59 ^ n55 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = n59 ^ x4 ;
  assign n63 = n62 ^ n59 ;
  assign n64 = n61 & ~n63 ;
  assign n65 = n64 ^ n59 ;
  assign n66 = x2 & ~n65 ;
  assign n67 = n66 ^ n59 ;
  assign n68 = x7 & ~n67 ;
  assign n69 = x4 & x7 ;
  assign n70 = x2 & x6 ;
  assign n71 = ~n69 & ~n70 ;
  assign n72 = x2 & x7 ;
  assign n73 = x5 & ~x8 ;
  assign n74 = ~n72 & n73 ;
  assign n75 = ~n71 & n74 ;
  assign n76 = ~n17 & n20 ;
  assign n77 = ~n73 & ~n76 ;
  assign n78 = ~x2 & ~n15 ;
  assign n79 = ~n77 & n78 ;
  assign n80 = x7 & n15 ;
  assign n81 = ~n69 & ~n80 ;
  assign n82 = n33 & ~n57 ;
  assign n83 = ~n81 & ~n82 ;
  assign n84 = ~x5 & x8 ;
  assign n85 = ~x5 & ~x7 ;
  assign n86 = ~x6 & n85 ;
  assign n87 = ~n10 & ~n86 ;
  assign n88 = x2 & ~n87 ;
  assign n89 = ~n84 & n88 ;
  assign n90 = ~n83 & ~n89 ;
  assign n91 = ~n79 & n90 ;
  assign n92 = x3 & ~n91 ;
  assign n93 = ~n75 & ~n92 ;
  assign n94 = ~x1 & ~n93 ;
  assign n95 = n94 ^ n68 ;
  assign n96 = ~x7 & n39 ;
  assign n97 = n73 & n96 ;
  assign n98 = n97 ^ x3 ;
  assign n99 = n98 ^ n97 ;
  assign n102 = n69 ^ x4 ;
  assign n100 = n69 ^ x2 ;
  assign n103 = n102 ^ n100 ;
  assign n104 = n103 ^ n100 ;
  assign n114 = n104 ^ n69 ;
  assign n106 = n69 ^ x5 ;
  assign n107 = n106 ^ n100 ;
  assign n108 = n107 ^ x8 ;
  assign n109 = n108 ^ n107 ;
  assign n110 = n109 ^ n103 ;
  assign n111 = n110 ^ n100 ;
  assign n112 = n111 ^ n69 ;
  assign n115 = n114 ^ n112 ;
  assign n101 = n100 ^ n69 ;
  assign n105 = n101 & ~n104 ;
  assign n113 = n112 ^ n105 ;
  assign n116 = n115 ^ n113 ;
  assign n117 = n103 ^ n85 ;
  assign n118 = n117 ^ n107 ;
  assign n119 = n118 ^ n107 ;
  assign n120 = n115 ^ n112 ;
  assign n121 = n119 & n120 ;
  assign n122 = n121 ^ n118 ;
  assign n123 = n122 ^ n119 ;
  assign n124 = ~n115 & ~n123 ;
  assign n125 = n124 ^ n121 ;
  assign n126 = n116 & n125 ;
  assign n127 = n126 ^ n105 ;
  assign n128 = n127 ^ x2 ;
  assign n129 = n128 ^ n114 ;
  assign n130 = ~x6 & n129 ;
  assign n131 = n33 & n84 ;
  assign n132 = ~x4 & ~n10 ;
  assign n133 = ~n73 & ~n85 ;
  assign n134 = n132 & n133 ;
  assign n135 = ~n131 & ~n134 ;
  assign n136 = ~n130 & n135 ;
  assign n137 = ~x1 & ~n136 ;
  assign n138 = x6 ^ x4 ;
  assign n139 = n138 ^ x6 ;
  assign n140 = n54 ^ x6 ;
  assign n141 = n139 & ~n140 ;
  assign n142 = n141 ^ x6 ;
  assign n143 = n72 & ~n142 ;
  assign n144 = ~x8 & n143 ;
  assign n145 = ~x7 & x8 ;
  assign n146 = n12 & n145 ;
  assign n147 = n17 & n69 ;
  assign n148 = ~x4 & n70 ;
  assign n149 = ~n147 & ~n148 ;
  assign n150 = n149 ^ x5 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = n151 ^ n146 ;
  assign n153 = n40 ^ x7 ;
  assign n154 = ~x7 & ~n153 ;
  assign n155 = n154 ^ n149 ;
  assign n156 = n155 ^ x7 ;
  assign n157 = n152 & n156 ;
  assign n158 = n157 ^ n154 ;
  assign n159 = n158 ^ x7 ;
  assign n160 = ~n146 & ~n159 ;
  assign n161 = n160 ^ n146 ;
  assign n162 = ~n144 & ~n161 ;
  assign n163 = ~n137 & n162 ;
  assign n164 = n163 ^ n97 ;
  assign n165 = ~n99 & ~n164 ;
  assign n166 = n165 ^ n97 ;
  assign n167 = n166 ^ n68 ;
  assign n168 = n95 & n167 ;
  assign n169 = n168 ^ n165 ;
  assign n170 = n169 ^ n97 ;
  assign n171 = n170 ^ n94 ;
  assign n172 = ~n68 & n171 ;
  assign n173 = n172 ^ n68 ;
  assign n174 = ~n52 & ~n173 ;
  assign n175 = ~x0 & ~n174 ;
  assign n176 = ~x1 & ~x3 ;
  assign n177 = n30 & n85 ;
  assign n178 = n139 ^ x7 ;
  assign n179 = x7 ^ x6 ;
  assign n180 = n179 ^ x6 ;
  assign n181 = x8 ^ x6 ;
  assign n182 = n181 ^ x6 ;
  assign n183 = n180 & ~n182 ;
  assign n184 = n183 ^ x6 ;
  assign n185 = n178 & n184 ;
  assign n186 = n185 ^ n138 ;
  assign n187 = n186 ^ x5 ;
  assign n188 = n187 ^ n186 ;
  assign n189 = ~x4 & ~n17 ;
  assign n190 = x4 & ~n145 ;
  assign n191 = ~n28 & n190 ;
  assign n192 = ~n189 & ~n191 ;
  assign n193 = n192 ^ n186 ;
  assign n194 = n188 & ~n193 ;
  assign n195 = n194 ^ n186 ;
  assign n196 = x0 & ~n195 ;
  assign n197 = ~n177 & ~n196 ;
  assign n198 = n176 & ~n197 ;
  assign n199 = ~x2 & n198 ;
  assign n200 = ~n175 & ~n199 ;
  assign y0 = ~n200 ;
endmodule
