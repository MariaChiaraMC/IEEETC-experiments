module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 ;
  assign n16 = ~x9 & ~x14 ;
  assign n17 = x6 ^ x4 ;
  assign n18 = x8 ^ x4 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = n17 & n19 ;
  assign n21 = n20 ^ x4 ;
  assign n22 = ~x4 & ~x7 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = ~n21 & n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n16 & n25 ;
  assign n27 = n26 ^ n16 ;
  assign n28 = x3 & ~n27 ;
  assign n29 = ~x0 & ~x2 ;
  assign n30 = ~x11 & n29 ;
  assign n31 = ~x10 & n30 ;
  assign n32 = ~x12 & n31 ;
  assign n33 = ~n28 & n32 ;
  assign n34 = ~x7 & ~x8 ;
  assign n35 = ~x6 & n34 ;
  assign n36 = ~x3 & ~n35 ;
  assign n37 = x8 ^ x6 ;
  assign n38 = ~x7 & ~n37 ;
  assign n39 = n38 ^ x6 ;
  assign n40 = x4 & n39 ;
  assign n41 = ~x1 & ~x5 ;
  assign n42 = x14 ^ x13 ;
  assign n43 = n41 & ~n42 ;
  assign n44 = ~n40 & n43 ;
  assign n45 = ~n36 & n44 ;
  assign n46 = n45 ^ x9 ;
  assign n47 = n46 ^ n45 ;
  assign n48 = x4 & n34 ;
  assign n49 = ~x13 & x14 ;
  assign n50 = x1 & x5 ;
  assign n51 = x6 & n50 ;
  assign n52 = n49 & n51 ;
  assign n53 = n48 & n52 ;
  assign n54 = n53 ^ n45 ;
  assign n55 = n47 & n54 ;
  assign n56 = n55 ^ n45 ;
  assign n57 = n33 & n56 ;
  assign y0 = n57 ;
endmodule
