module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 ;
  assign n9 = ~x4 & x5 ;
  assign n10 = ~x1 & ~x3 ;
  assign n11 = ~x0 & ~x7 ;
  assign n12 = n10 & n11 ;
  assign n13 = n9 & n12 ;
  assign n24 = x6 & x7 ;
  assign n68 = x1 & n24 ;
  assign n53 = x0 & ~x3 ;
  assign n69 = n9 & n53 ;
  assign n70 = n68 & n69 ;
  assign n35 = ~x5 & ~x6 ;
  assign n36 = ~x0 & n35 ;
  assign n116 = ~x4 & n36 ;
  assign n73 = x6 ^ x5 ;
  assign n71 = x4 ^ x0 ;
  assign n72 = n71 ^ x6 ;
  assign n84 = n73 ^ n72 ;
  assign n80 = n73 ^ x3 ;
  assign n81 = n80 ^ x4 ;
  assign n85 = n84 ^ n81 ;
  assign n86 = n85 ^ n81 ;
  assign n75 = n73 ^ x0 ;
  assign n76 = n75 ^ x6 ;
  assign n87 = n76 ^ n73 ;
  assign n88 = n87 ^ n81 ;
  assign n89 = ~n86 & n88 ;
  assign n74 = n73 ^ x6 ;
  assign n77 = n76 ^ n74 ;
  assign n78 = n77 ^ n73 ;
  assign n79 = n78 ^ n72 ;
  assign n82 = n81 ^ n79 ;
  assign n83 = n72 & n82 ;
  assign n90 = n89 ^ n83 ;
  assign n91 = n90 ^ n72 ;
  assign n92 = n83 ^ n81 ;
  assign n93 = n92 ^ n85 ;
  assign n94 = n81 & ~n93 ;
  assign n95 = n94 ^ n83 ;
  assign n96 = n91 & n95 ;
  assign n97 = n96 ^ n89 ;
  assign n98 = n97 ^ n94 ;
  assign n99 = n98 ^ n72 ;
  assign n100 = n99 ^ n81 ;
  assign n101 = n100 ^ n85 ;
  assign n102 = n101 ^ x3 ;
  assign n103 = n102 ^ n101 ;
  assign n104 = ~x0 & x6 ;
  assign n105 = x0 & ~x6 ;
  assign n106 = n9 & ~n105 ;
  assign n107 = ~n104 & n106 ;
  assign n108 = x0 & n35 ;
  assign n109 = ~n107 & ~n108 ;
  assign n110 = n109 ^ n101 ;
  assign n111 = n110 ^ n101 ;
  assign n112 = n103 & ~n111 ;
  assign n113 = n112 ^ n101 ;
  assign n114 = x1 & ~n113 ;
  assign n115 = n114 ^ n101 ;
  assign n117 = n116 ^ n115 ;
  assign n118 = n117 ^ x7 ;
  assign n125 = n118 ^ n117 ;
  assign n119 = n118 ^ n10 ;
  assign n120 = n119 ^ n117 ;
  assign n121 = n116 ^ n10 ;
  assign n122 = n121 ^ n10 ;
  assign n123 = n122 ^ n120 ;
  assign n124 = n120 & n123 ;
  assign n126 = n125 ^ n124 ;
  assign n127 = n126 ^ n120 ;
  assign n34 = x1 & x3 ;
  assign n128 = n117 ^ n34 ;
  assign n129 = n124 ^ n120 ;
  assign n130 = n128 & n129 ;
  assign n131 = n130 ^ n117 ;
  assign n132 = ~n127 & ~n131 ;
  assign n133 = n132 ^ n117 ;
  assign n134 = n133 ^ n116 ;
  assign n135 = n134 ^ n117 ;
  assign n136 = ~n70 & ~n135 ;
  assign n14 = x5 & x6 ;
  assign n15 = n12 & n14 ;
  assign n16 = x3 & ~x5 ;
  assign n17 = ~x0 & x1 ;
  assign n18 = x7 ^ x6 ;
  assign n19 = ~x7 & n18 ;
  assign n20 = ~x3 & n19 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n17 & n21 ;
  assign n23 = x0 & x3 ;
  assign n25 = ~x6 & x7 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = x1 & n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n23 & n28 ;
  assign n30 = ~n22 & ~n29 ;
  assign n31 = ~n16 & ~n30 ;
  assign n32 = n31 ^ x4 ;
  assign n33 = n32 ^ n31 ;
  assign n37 = n34 & n36 ;
  assign n38 = x0 & n21 ;
  assign n39 = ~n16 & n38 ;
  assign n40 = n39 ^ n24 ;
  assign n41 = n40 ^ x1 ;
  assign n50 = n41 ^ n40 ;
  assign n42 = ~x3 & n17 ;
  assign n43 = x5 & n42 ;
  assign n44 = n43 ^ n41 ;
  assign n45 = n44 ^ n40 ;
  assign n46 = n41 ^ n39 ;
  assign n47 = n46 ^ n43 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = ~n45 & ~n48 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = n51 ^ n45 ;
  assign n54 = ~n16 & ~n53 ;
  assign n55 = n54 ^ n40 ;
  assign n56 = n49 ^ n45 ;
  assign n57 = n55 & ~n56 ;
  assign n58 = n57 ^ n40 ;
  assign n59 = ~n52 & n58 ;
  assign n60 = n59 ^ n40 ;
  assign n61 = n60 ^ n24 ;
  assign n62 = n61 ^ n40 ;
  assign n63 = ~n37 & ~n62 ;
  assign n64 = n63 ^ n31 ;
  assign n65 = n33 & ~n64 ;
  assign n66 = n65 ^ n31 ;
  assign n67 = ~n15 & ~n66 ;
  assign n137 = n136 ^ n67 ;
  assign n138 = x2 & n137 ;
  assign n139 = n138 ^ n67 ;
  assign n140 = ~n13 & n139 ;
  assign y0 = ~n140 ;
endmodule
