module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 ;
  assign n8 = x1 & x3 ;
  assign n9 = ~x5 & ~n8 ;
  assign n10 = ~x4 & x6 ;
  assign n11 = ~n9 & n10 ;
  assign n12 = x3 & ~x5 ;
  assign n13 = x3 ^ x2 ;
  assign n14 = x3 ^ x1 ;
  assign n15 = n13 & n14 ;
  assign n16 = n15 ^ x0 ;
  assign n17 = n12 & n16 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = x0 & n18 ;
  assign n20 = n19 ^ x0 ;
  assign n21 = n11 & ~n20 ;
  assign y0 = n21 ;
endmodule
