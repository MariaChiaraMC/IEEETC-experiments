module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 ;
  assign n23 = x17 ^ x3 ;
  assign n35 = n23 ^ x3 ;
  assign n22 = x3 ^ x2 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ x3 ;
  assign n27 = x18 & x19 ;
  assign n28 = ~x17 & n27 ;
  assign n29 = ~x20 & n28 ;
  assign n30 = x1 & ~n29 ;
  assign n31 = n30 ^ n24 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = n32 ^ n26 ;
  assign n34 = n26 & ~n33 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = n36 ^ n26 ;
  assign n38 = x16 ^ x3 ;
  assign n39 = n34 ^ n26 ;
  assign n40 = n38 & n39 ;
  assign n41 = n40 ^ x3 ;
  assign n42 = n37 & ~n41 ;
  assign n43 = n42 ^ x3 ;
  assign n44 = n43 ^ x17 ;
  assign n45 = n44 ^ x3 ;
  assign n46 = ~x15 & n45 ;
  assign n47 = x16 & x20 ;
  assign n48 = n27 & n47 ;
  assign n49 = x3 & ~n48 ;
  assign n50 = ~n46 & ~n49 ;
  assign n51 = ~x0 & ~n50 ;
  assign y0 = n51 ;
endmodule
