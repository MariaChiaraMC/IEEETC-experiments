module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 ;
  assign n9 = ~x3 & ~x4 ;
  assign n10 = ~x2 & x7 ;
  assign n11 = ~x2 & ~x5 ;
  assign n12 = ~n10 & ~n11 ;
  assign n13 = ~x6 & ~n12 ;
  assign n14 = n9 & n13 ;
  assign n18 = x2 & x5 ;
  assign n15 = x6 ^ x4 ;
  assign n16 = n12 & n15 ;
  assign n17 = n16 ^ x3 ;
  assign n19 = n18 ^ n17 ;
  assign n28 = n19 ^ n17 ;
  assign n20 = x4 & ~x6 ;
  assign n21 = n10 & n20 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ n17 ;
  assign n24 = n19 ^ n16 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n23 & ~n26 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = n17 ^ x4 ;
  assign n32 = n27 ^ n23 ;
  assign n33 = n31 & n32 ;
  assign n34 = n33 ^ n17 ;
  assign n35 = ~n30 & n34 ;
  assign n36 = n35 ^ n17 ;
  assign n37 = n36 ^ x3 ;
  assign n38 = n37 ^ n17 ;
  assign n39 = x7 ^ x4 ;
  assign n40 = n39 ^ x7 ;
  assign n44 = ~x3 & ~x5 ;
  assign n41 = n11 ^ x7 ;
  assign n42 = x7 & ~n41 ;
  assign n47 = n44 ^ n42 ;
  assign n43 = n42 ^ x7 ;
  assign n45 = n44 ^ n40 ;
  assign n46 = n43 & n45 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = n40 & n48 ;
  assign n50 = n49 ^ n42 ;
  assign n51 = n50 ^ n46 ;
  assign n52 = ~n38 & ~n51 ;
  assign n53 = ~n14 & n52 ;
  assign n54 = n53 ^ x2 ;
  assign n55 = n54 ^ x1 ;
  assign n68 = n55 ^ n54 ;
  assign n56 = x1 & x7 ;
  assign n57 = x7 ^ x3 ;
  assign n58 = x4 & n57 ;
  assign n59 = ~n56 & ~n58 ;
  assign n60 = x6 & ~n59 ;
  assign n61 = x5 & n60 ;
  assign n62 = n61 ^ n55 ;
  assign n63 = n62 ^ n54 ;
  assign n64 = n55 ^ n53 ;
  assign n65 = n64 ^ n61 ;
  assign n66 = n65 ^ n63 ;
  assign n67 = n63 & n66 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = n69 ^ n63 ;
  assign n71 = n54 ^ n9 ;
  assign n72 = n67 ^ n63 ;
  assign n73 = n71 & n72 ;
  assign n74 = n73 ^ n54 ;
  assign n75 = ~n70 & n74 ;
  assign n76 = n75 ^ n54 ;
  assign n77 = n76 ^ x2 ;
  assign n78 = n77 ^ n54 ;
  assign n79 = ~x0 & ~n78 ;
  assign y0 = n79 ;
endmodule
