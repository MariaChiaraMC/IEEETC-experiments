module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n17 = x5 & ~x7 ;
  assign n18 = x5 & ~x6 ;
  assign n19 = ~x8 & ~x9 ;
  assign n20 = x11 ^ x10 ;
  assign n21 = n19 & n20 ;
  assign n22 = n18 & n21 ;
  assign n23 = ~n17 & ~n22 ;
  assign n24 = x6 ^ x5 ;
  assign n25 = x7 ^ x6 ;
  assign n26 = n25 ^ x7 ;
  assign n27 = ~x10 & ~x11 ;
  assign n28 = n27 ^ x7 ;
  assign n29 = ~n26 & n28 ;
  assign n30 = n29 ^ x7 ;
  assign n31 = n24 & n30 ;
  assign n32 = x9 ^ x8 ;
  assign n33 = n31 & n32 ;
  assign n34 = n23 & ~n33 ;
  assign y0 = ~n34 ;
endmodule
