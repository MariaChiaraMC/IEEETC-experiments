module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 ;
  assign n9 = x4 & x5 ;
  assign n10 = x3 & ~x7 ;
  assign n11 = n9 & n10 ;
  assign n12 = ~x2 & x6 ;
  assign n13 = ~x1 & n12 ;
  assign n14 = n11 & n13 ;
  assign n15 = x1 & ~x2 ;
  assign n16 = x4 ^ x3 ;
  assign n17 = n16 ^ x4 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = x7 ^ x5 ;
  assign n20 = n19 ^ x5 ;
  assign n21 = x5 ^ x4 ;
  assign n22 = n21 ^ x5 ;
  assign n23 = ~n20 & ~n22 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = ~n18 & n24 ;
  assign n26 = n25 ^ n16 ;
  assign n27 = n15 & ~n26 ;
  assign n28 = ~x4 & ~x5 ;
  assign n29 = x7 & n28 ;
  assign n30 = x3 & n29 ;
  assign n31 = ~x4 & ~x7 ;
  assign n32 = ~x5 & n31 ;
  assign n33 = x3 ^ x1 ;
  assign n34 = x3 & ~n33 ;
  assign n35 = n34 ^ x3 ;
  assign n36 = x4 & x7 ;
  assign n37 = n36 ^ x3 ;
  assign n38 = n35 & n37 ;
  assign n39 = n38 ^ n34 ;
  assign n40 = n39 ^ x3 ;
  assign n41 = n40 ^ x1 ;
  assign n42 = ~n32 & ~n41 ;
  assign n43 = n42 ^ x1 ;
  assign n44 = ~n30 & n43 ;
  assign n45 = x2 & ~n44 ;
  assign n46 = ~n27 & ~n45 ;
  assign n47 = x6 & ~n46 ;
  assign n48 = ~n14 & ~n47 ;
  assign n49 = ~x2 & ~x6 ;
  assign n50 = ~n11 & ~n29 ;
  assign n51 = n50 ^ x1 ;
  assign n52 = n51 ^ n50 ;
  assign n53 = x3 & ~x5 ;
  assign n54 = n31 & ~n53 ;
  assign n55 = n54 ^ n50 ;
  assign n56 = ~n52 & ~n55 ;
  assign n57 = n56 ^ n50 ;
  assign n58 = n49 & ~n57 ;
  assign n59 = n48 & ~n58 ;
  assign n60 = x0 & ~n59 ;
  assign n61 = x2 & ~x6 ;
  assign n62 = x1 & ~x3 ;
  assign n63 = n32 & n62 ;
  assign n64 = n61 & n63 ;
  assign n65 = ~n60 & ~n64 ;
  assign n66 = n13 & n30 ;
  assign n67 = x5 & ~n31 ;
  assign n68 = n13 & ~n28 ;
  assign n69 = ~n67 & n68 ;
  assign n70 = x4 & x6 ;
  assign n71 = ~x1 & ~n70 ;
  assign n73 = n71 ^ x2 ;
  assign n72 = n71 ^ x6 ;
  assign n74 = n73 ^ n72 ;
  assign n79 = n74 ^ n73 ;
  assign n75 = n74 ^ x4 ;
  assign n76 = n75 ^ n71 ;
  assign n77 = n76 ^ x5 ;
  assign n78 = n77 ^ n73 ;
  assign n80 = n79 ^ n78 ;
  assign n83 = n77 ^ x5 ;
  assign n81 = n71 ^ x5 ;
  assign n82 = n81 ^ n78 ;
  assign n84 = n83 ^ n82 ;
  assign n85 = n80 & ~n84 ;
  assign n86 = n85 ^ n77 ;
  assign n87 = n86 ^ n81 ;
  assign n88 = n87 ^ n83 ;
  assign n89 = n82 ^ n79 ;
  assign n90 = ~n86 & n89 ;
  assign n91 = n90 ^ n77 ;
  assign n92 = n91 ^ n78 ;
  assign n93 = n92 ^ n79 ;
  assign n94 = ~n88 & ~n93 ;
  assign n95 = x7 & n94 ;
  assign n96 = ~x3 & ~n95 ;
  assign n97 = ~n69 & n96 ;
  assign n98 = x6 ^ x2 ;
  assign n99 = x7 ^ x4 ;
  assign n100 = ~n98 & n99 ;
  assign n101 = n100 ^ x2 ;
  assign n102 = n101 ^ n100 ;
  assign n103 = n100 ^ n70 ;
  assign n104 = n103 ^ n100 ;
  assign n105 = ~n102 & n104 ;
  assign n106 = n105 ^ n100 ;
  assign n107 = x1 & n106 ;
  assign n108 = n107 ^ n100 ;
  assign n109 = n108 ^ x5 ;
  assign n110 = n109 ^ n108 ;
  assign n111 = n110 ^ x3 ;
  assign n112 = n49 ^ n31 ;
  assign n113 = n31 & n112 ;
  assign n114 = n113 ^ n108 ;
  assign n115 = n114 ^ n31 ;
  assign n116 = ~n111 & n115 ;
  assign n117 = n116 ^ n113 ;
  assign n118 = n117 ^ n31 ;
  assign n119 = x3 & n118 ;
  assign n120 = n119 ^ x3 ;
  assign n121 = ~x0 & ~n120 ;
  assign n122 = ~n97 & n121 ;
  assign n123 = ~n66 & ~n122 ;
  assign n124 = n65 & n123 ;
  assign y0 = ~n124 ;
endmodule
