module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n8 = x6 ^ x4 ;
  assign n9 = x6 ^ x5 ;
  assign n10 = n9 ^ n8 ;
  assign n11 = ~x1 & ~x2 ;
  assign n12 = ~x0 & n11 ;
  assign n13 = x3 & ~n12 ;
  assign n14 = n13 ^ x6 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = x1 & x2 ;
  assign n17 = ~x3 & ~n16 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = n15 & n18 ;
  assign n20 = n19 ^ n13 ;
  assign n21 = n20 ^ n8 ;
  assign n22 = ~n10 & n21 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n23 ^ n13 ;
  assign n25 = n24 ^ n9 ;
  assign n26 = ~n8 & ~n25 ;
  assign n27 = n26 ^ n8 ;
  assign n28 = n27 ^ n9 ;
  assign y0 = ~n28 ;
endmodule
