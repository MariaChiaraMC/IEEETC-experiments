module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n11 = x8 ^ x7 ;
  assign n15 = n11 ^ x8 ;
  assign n13 = x8 ^ x1 ;
  assign n12 = n11 ^ x3 ;
  assign n14 = n13 ^ n12 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n15 ^ x8 ;
  assign n18 = ~n16 & ~n17 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = n19 ^ x8 ;
  assign n22 = n14 ^ n13 ;
  assign n23 = n22 ^ x8 ;
  assign n24 = ~n22 & ~n23 ;
  assign n21 = ~x0 & ~x2 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ n13 ;
  assign n27 = n26 ^ n14 ;
  assign n28 = ~n15 & ~n27 ;
  assign n29 = n28 ^ n21 ;
  assign n30 = n29 ^ x8 ;
  assign n31 = ~n20 & n30 ;
  assign n32 = n31 ^ n21 ;
  assign n33 = n32 ^ n24 ;
  assign n34 = n33 ^ n28 ;
  assign n35 = n34 ^ n13 ;
  assign n36 = n35 ^ n14 ;
  assign n37 = n36 ^ x7 ;
  assign n38 = n37 ^ x8 ;
  assign y0 = ~n38 ;
endmodule
