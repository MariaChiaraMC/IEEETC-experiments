module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 ;
  assign n17 = ~x0 & ~x2 ;
  assign n18 = n17 ^ x1 ;
  assign n19 = ~x9 & ~x10 ;
  assign n20 = x9 & x10 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = ~x6 & ~x8 ;
  assign n23 = x6 & x11 ;
  assign n24 = x4 & n23 ;
  assign n25 = ~n22 & ~n24 ;
  assign n26 = ~x8 & x11 ;
  assign n27 = ~x12 & x13 ;
  assign n28 = n26 & ~n27 ;
  assign n29 = ~n25 & ~n28 ;
  assign n30 = ~x14 & x15 ;
  assign n31 = ~n27 & ~n30 ;
  assign n32 = ~x1 & ~n31 ;
  assign n33 = x5 & x7 ;
  assign n34 = ~x4 & ~x11 ;
  assign n35 = n27 & ~n34 ;
  assign n36 = n33 & ~n35 ;
  assign n37 = n32 & n36 ;
  assign n38 = n29 & n37 ;
  assign n39 = ~x14 & ~x15 ;
  assign n40 = x4 & ~x12 ;
  assign n41 = ~x5 & ~x7 ;
  assign n42 = ~x6 & ~x13 ;
  assign n43 = n41 & n42 ;
  assign n44 = x8 & ~x11 ;
  assign n45 = x1 & n44 ;
  assign n46 = n43 & n45 ;
  assign n47 = n40 & n46 ;
  assign n48 = n39 & n47 ;
  assign n49 = ~n38 & ~n48 ;
  assign n50 = n21 & ~n49 ;
  assign n51 = x8 & ~x9 ;
  assign n52 = ~x8 & x9 ;
  assign n53 = ~n51 & ~n52 ;
  assign n54 = x6 & ~n53 ;
  assign n55 = x7 & ~n54 ;
  assign n56 = x7 & ~n27 ;
  assign n57 = n32 & ~n56 ;
  assign n58 = ~x6 & n52 ;
  assign n59 = x13 & x15 ;
  assign n60 = ~x7 & n59 ;
  assign n61 = ~n58 & ~n60 ;
  assign n62 = ~x12 & ~x14 ;
  assign n63 = ~n61 & n62 ;
  assign n64 = ~x10 & ~n63 ;
  assign n65 = n57 & n64 ;
  assign n66 = ~n55 & n65 ;
  assign n67 = ~x12 & ~n19 ;
  assign n68 = ~x7 & n22 ;
  assign n69 = n67 & n68 ;
  assign n70 = ~x13 & ~n30 ;
  assign n71 = ~x10 & ~n70 ;
  assign n72 = ~x1 & ~n71 ;
  assign n73 = n72 ^ n69 ;
  assign n74 = n39 ^ x13 ;
  assign n75 = n74 ^ n39 ;
  assign n76 = x14 & x15 ;
  assign n77 = ~n39 & ~n76 ;
  assign n78 = n77 ^ n39 ;
  assign n79 = ~n75 & n78 ;
  assign n80 = n79 ^ n39 ;
  assign n81 = n80 ^ n69 ;
  assign n82 = ~n73 & n81 ;
  assign n83 = n82 ^ n79 ;
  assign n84 = n83 ^ n39 ;
  assign n85 = n84 ^ n72 ;
  assign n86 = n69 & ~n85 ;
  assign n87 = n86 ^ n69 ;
  assign n88 = ~n66 & ~n87 ;
  assign n89 = ~x11 & ~n88 ;
  assign n90 = ~x5 & n89 ;
  assign n91 = ~x6 & x7 ;
  assign n92 = ~x5 & n91 ;
  assign n93 = x1 & n92 ;
  assign n94 = ~n90 & ~n93 ;
  assign n95 = x4 & ~n94 ;
  assign n96 = ~n50 & ~n95 ;
  assign n97 = n96 ^ n18 ;
  assign n98 = n97 ^ n17 ;
  assign n99 = n98 ^ n97 ;
  assign n100 = x0 & x4 ;
  assign n101 = ~x5 & n100 ;
  assign n102 = n101 ^ n97 ;
  assign n103 = n102 ^ n18 ;
  assign n104 = n99 & n103 ;
  assign n105 = n104 ^ n101 ;
  assign n106 = ~x10 & ~x11 ;
  assign n107 = n41 & ~n106 ;
  assign n108 = ~n92 & ~n107 ;
  assign n109 = ~n30 & ~n108 ;
  assign n110 = ~x15 & ~n106 ;
  assign n111 = x6 & ~n110 ;
  assign n112 = n33 & ~n111 ;
  assign n113 = ~x7 & x10 ;
  assign n114 = ~n106 & ~n113 ;
  assign n115 = x5 & x6 ;
  assign n116 = n76 & n115 ;
  assign n117 = n114 & n116 ;
  assign n118 = ~n112 & ~n117 ;
  assign n119 = ~n109 & n118 ;
  assign n120 = n27 & ~n119 ;
  assign n121 = x12 & n106 ;
  assign n122 = x13 & ~n121 ;
  assign n123 = n41 & n122 ;
  assign n124 = x13 & ~n92 ;
  assign n125 = ~n108 & ~n124 ;
  assign n126 = x11 & ~n21 ;
  assign n127 = ~n26 & ~n27 ;
  assign n128 = ~n126 & n127 ;
  assign n129 = n128 ^ x6 ;
  assign n130 = n129 ^ n128 ;
  assign n131 = n51 ^ x11 ;
  assign n132 = n51 ^ x10 ;
  assign n133 = n132 ^ x10 ;
  assign n134 = n19 ^ x10 ;
  assign n135 = ~n133 & n134 ;
  assign n136 = n135 ^ x10 ;
  assign n137 = n131 & n136 ;
  assign n138 = n137 ^ x11 ;
  assign n139 = ~n27 & n138 ;
  assign n140 = n139 ^ n128 ;
  assign n141 = ~n130 & ~n140 ;
  assign n142 = n141 ^ n128 ;
  assign n143 = n33 & ~n142 ;
  assign n144 = ~n125 & ~n143 ;
  assign n145 = ~n123 & n144 ;
  assign n146 = n30 & ~n145 ;
  assign n147 = x15 ^ x14 ;
  assign n148 = n113 & n115 ;
  assign n149 = ~x13 & n148 ;
  assign n150 = x12 & n149 ;
  assign n151 = ~x6 & ~n20 ;
  assign n152 = n151 ^ x5 ;
  assign n153 = n152 ^ n56 ;
  assign n154 = n53 ^ x5 ;
  assign n155 = n154 ^ x10 ;
  assign n156 = ~x10 & n155 ;
  assign n157 = n156 ^ x5 ;
  assign n158 = n157 ^ x10 ;
  assign n159 = ~n153 & ~n158 ;
  assign n160 = n159 ^ n156 ;
  assign n161 = n160 ^ x10 ;
  assign n162 = n56 & ~n161 ;
  assign n163 = ~n150 & ~n162 ;
  assign n164 = n163 ^ x15 ;
  assign n165 = n164 ^ n163 ;
  assign n166 = n165 ^ n147 ;
  assign n167 = n148 ^ n27 ;
  assign n168 = n148 & n167 ;
  assign n169 = n168 ^ n163 ;
  assign n170 = n169 ^ n148 ;
  assign n171 = ~n166 & ~n170 ;
  assign n172 = n171 ^ n168 ;
  assign n173 = n172 ^ n148 ;
  assign n174 = n147 & n173 ;
  assign n175 = ~x11 & n174 ;
  assign n176 = ~n146 & ~n175 ;
  assign n177 = ~n120 & n176 ;
  assign n178 = x4 & ~n177 ;
  assign n193 = x6 & x7 ;
  assign n194 = n51 & n193 ;
  assign n195 = ~x4 & n194 ;
  assign n179 = x13 ^ x7 ;
  assign n180 = n179 ^ x13 ;
  assign n181 = n106 ^ x13 ;
  assign n182 = n180 & n181 ;
  assign n183 = n182 ^ x13 ;
  assign n184 = x6 & n183 ;
  assign n185 = n184 ^ x7 ;
  assign n186 = ~x4 & ~n185 ;
  assign n187 = ~n26 & ~n44 ;
  assign n188 = ~x13 & n19 ;
  assign n189 = ~n187 & n188 ;
  assign n190 = n91 & n189 ;
  assign n191 = ~n186 & ~n190 ;
  assign n192 = n30 & ~n191 ;
  assign n196 = n195 ^ n192 ;
  assign n197 = n196 ^ n195 ;
  assign n198 = x6 & ~x11 ;
  assign n199 = ~n30 & n198 ;
  assign n200 = ~x9 & ~n187 ;
  assign n201 = x7 & ~n200 ;
  assign n202 = ~n40 & ~n193 ;
  assign n203 = ~n201 & n202 ;
  assign n204 = ~n199 & ~n203 ;
  assign n205 = ~x6 & n30 ;
  assign n206 = ~x7 & n205 ;
  assign n207 = ~x7 & ~n23 ;
  assign n208 = n207 ^ x4 ;
  assign n209 = ~x10 & n208 ;
  assign n210 = n208 ^ n207 ;
  assign n211 = x11 & x12 ;
  assign n212 = n211 ^ n209 ;
  assign n213 = n210 & n212 ;
  assign n214 = n213 ^ n211 ;
  assign n215 = n209 & n214 ;
  assign n216 = n215 ^ x4 ;
  assign n217 = ~n206 & ~n216 ;
  assign n218 = x12 & ~n30 ;
  assign n219 = x7 & x10 ;
  assign n220 = ~n218 & ~n219 ;
  assign n221 = x13 & n220 ;
  assign n222 = n217 & n221 ;
  assign n223 = ~n204 & n222 ;
  assign n224 = n223 ^ n195 ;
  assign n225 = n224 ^ n195 ;
  assign n226 = ~n197 & ~n225 ;
  assign n227 = n226 ^ n195 ;
  assign n228 = x5 & ~n227 ;
  assign n229 = n228 ^ n195 ;
  assign n230 = ~n178 & ~n229 ;
  assign n231 = ~n101 & n230 ;
  assign n232 = n231 ^ n18 ;
  assign n233 = ~n105 & n232 ;
  assign n234 = n233 ^ n231 ;
  assign n235 = n18 & n234 ;
  assign n236 = n235 ^ n104 ;
  assign n237 = n236 ^ x1 ;
  assign n238 = n237 ^ n101 ;
  assign n239 = ~x3 & n238 ;
  assign y0 = n239 ;
endmodule
