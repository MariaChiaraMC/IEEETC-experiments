module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 ;
  assign n9 = x3 ^ x2 ;
  assign n10 = n9 ^ x5 ;
  assign n11 = x6 ^ x5 ;
  assign n12 = n11 ^ x6 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n11 ^ x3 ;
  assign n15 = ~n13 & n14 ;
  assign n16 = n15 ^ n11 ;
  assign n17 = ~x7 & n11 ;
  assign n18 = n17 ^ n10 ;
  assign n19 = n16 & ~n18 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = ~n10 & n20 ;
  assign n22 = n21 ^ x3 ;
  assign n23 = n22 ^ n10 ;
  assign n24 = ~x4 & ~n23 ;
  assign n25 = ~x2 & ~x5 ;
  assign n26 = n25 ^ x3 ;
  assign n27 = n26 ^ x4 ;
  assign n28 = x6 ^ x3 ;
  assign n29 = x4 ^ x3 ;
  assign n30 = x7 ^ x5 ;
  assign n31 = ~n29 & ~n30 ;
  assign n32 = n31 ^ x5 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n28 & n33 ;
  assign n35 = n34 ^ x3 ;
  assign n36 = n27 & ~n35 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = x4 & n37 ;
  assign n39 = ~n24 & ~n38 ;
  assign n40 = ~x1 & ~n39 ;
  assign y0 = ~n40 ;
endmodule
