module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 ;
  output y0 ;
  wire n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 ;
  assign n23 = x1 ^ x0 ;
  assign n24 = x2 ^ x1 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = x5 ^ x3 ;
  assign n28 = x5 ^ x1 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = ~n27 & ~n29 ;
  assign n31 = n30 ^ x5 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = n26 & ~n32 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ n27 ;
  assign n36 = n23 & ~n35 ;
  assign n37 = ~x4 & n36 ;
  assign n38 = ~x19 & ~x20 ;
  assign n39 = n38 ^ x18 ;
  assign n40 = n39 ^ x18 ;
  assign n41 = x1 & x2 ;
  assign n42 = x11 & x13 ;
  assign n43 = ~x8 & ~x10 ;
  assign n44 = ~x9 & n43 ;
  assign n45 = n42 & n44 ;
  assign n46 = ~x6 & ~x7 ;
  assign n47 = ~x8 & n46 ;
  assign n48 = x8 & x10 ;
  assign n49 = x9 & n48 ;
  assign n50 = ~n47 & ~n49 ;
  assign n51 = n50 ^ x12 ;
  assign n53 = ~x9 & ~x10 ;
  assign n52 = x11 & n47 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = n54 ^ n52 ;
  assign n56 = ~x11 & ~x13 ;
  assign n57 = n56 ^ n52 ;
  assign n58 = ~n55 & n57 ;
  assign n59 = n58 ^ n52 ;
  assign n60 = n59 ^ n50 ;
  assign n61 = n51 & ~n60 ;
  assign n62 = n61 ^ n58 ;
  assign n63 = n62 ^ n52 ;
  assign n64 = n63 ^ x12 ;
  assign n65 = ~n50 & ~n64 ;
  assign n66 = n65 ^ n50 ;
  assign n67 = ~n45 & n66 ;
  assign n68 = ~n41 & n67 ;
  assign n69 = x3 & ~n68 ;
  assign n70 = ~x12 & ~x13 ;
  assign n71 = x9 & n70 ;
  assign n72 = x0 & n71 ;
  assign n73 = ~n69 & ~n72 ;
  assign n74 = ~x4 & ~n73 ;
  assign n77 = x12 ^ x1 ;
  assign n78 = n77 ^ x1 ;
  assign n75 = x4 ^ x1 ;
  assign n76 = n75 ^ x1 ;
  assign n79 = n78 ^ n76 ;
  assign n80 = x13 ^ x1 ;
  assign n81 = n80 ^ x1 ;
  assign n82 = n81 ^ n78 ;
  assign n83 = ~n78 & ~n82 ;
  assign n84 = n83 ^ n78 ;
  assign n85 = ~n79 & ~n84 ;
  assign n86 = n85 ^ n83 ;
  assign n87 = n86 ^ x1 ;
  assign n88 = n87 ^ n78 ;
  assign n89 = ~x3 & n88 ;
  assign n90 = n89 ^ x1 ;
  assign n91 = n90 ^ x3 ;
  assign n92 = n91 ^ x2 ;
  assign n161 = n92 ^ n91 ;
  assign n94 = x16 & ~x17 ;
  assign n95 = n43 & n94 ;
  assign n96 = n46 ^ x11 ;
  assign n97 = x15 ^ x13 ;
  assign n98 = n97 ^ x15 ;
  assign n99 = x15 ^ x12 ;
  assign n100 = ~n98 & n99 ;
  assign n101 = n100 ^ x15 ;
  assign n102 = n101 ^ n46 ;
  assign n103 = n96 & ~n102 ;
  assign n104 = n103 ^ n100 ;
  assign n105 = n104 ^ x15 ;
  assign n106 = n105 ^ x11 ;
  assign n107 = n46 & ~n106 ;
  assign n108 = n107 ^ n46 ;
  assign n109 = n95 & n108 ;
  assign n110 = ~x1 & n109 ;
  assign n111 = n110 ^ x9 ;
  assign n112 = n111 ^ x2 ;
  assign n113 = n112 ^ n110 ;
  assign n125 = n113 ^ n111 ;
  assign n126 = n125 ^ n110 ;
  assign n127 = n126 ^ n110 ;
  assign n128 = ~x0 & x1 ;
  assign n129 = n128 ^ n111 ;
  assign n130 = n129 ^ n111 ;
  assign n131 = n130 ^ n110 ;
  assign n132 = ~n127 & ~n131 ;
  assign n114 = x13 & n43 ;
  assign n115 = ~x11 & n114 ;
  assign n116 = x11 & ~x12 ;
  assign n117 = ~x1 & n43 ;
  assign n118 = n117 ^ x10 ;
  assign n119 = n116 & n118 ;
  assign n120 = ~n115 & ~n119 ;
  assign n121 = n120 ^ n111 ;
  assign n122 = n121 ^ n113 ;
  assign n123 = n122 ^ n110 ;
  assign n124 = n113 & ~n123 ;
  assign n133 = n132 ^ n124 ;
  assign n134 = n133 ^ n113 ;
  assign n135 = n124 ^ n110 ;
  assign n136 = n135 ^ n126 ;
  assign n137 = n110 & ~n136 ;
  assign n138 = n137 ^ n124 ;
  assign n139 = n134 & n138 ;
  assign n140 = n139 ^ n132 ;
  assign n141 = n140 ^ n137 ;
  assign n142 = n141 ^ n113 ;
  assign n143 = n142 ^ n110 ;
  assign n144 = n143 ^ n126 ;
  assign n145 = n144 ^ x9 ;
  assign n146 = n145 ^ x0 ;
  assign n147 = n145 ^ x13 ;
  assign n148 = n145 ^ x4 ;
  assign n149 = n145 & n148 ;
  assign n150 = n149 ^ n145 ;
  assign n151 = n147 & n150 ;
  assign n152 = n151 ^ n149 ;
  assign n153 = n152 ^ n145 ;
  assign n154 = n153 ^ x4 ;
  assign n155 = ~n146 & n154 ;
  assign n156 = n155 ^ x0 ;
  assign n93 = n92 ^ n90 ;
  assign n157 = n156 ^ n93 ;
  assign n158 = n156 ^ n92 ;
  assign n159 = n158 ^ n91 ;
  assign n160 = n157 & n159 ;
  assign n162 = n161 ^ n160 ;
  assign n163 = ~x1 & x21 ;
  assign n164 = ~x4 & n163 ;
  assign n165 = n164 ^ n92 ;
  assign n166 = ~n161 & ~n165 ;
  assign n167 = n166 ^ n164 ;
  assign n168 = ~n162 & n167 ;
  assign n169 = n168 ^ n160 ;
  assign n170 = n169 ^ n92 ;
  assign n171 = n170 ^ x3 ;
  assign n172 = n171 ^ n91 ;
  assign n173 = ~n74 & ~n172 ;
  assign n174 = x5 & ~n173 ;
  assign n187 = x2 & ~x4 ;
  assign n188 = ~x11 & n47 ;
  assign n189 = ~n53 & n188 ;
  assign n190 = ~x11 & n48 ;
  assign n191 = ~x10 & x11 ;
  assign n192 = x8 & n191 ;
  assign n193 = n46 & n192 ;
  assign n194 = ~n190 & ~n193 ;
  assign n195 = x9 & ~n194 ;
  assign n196 = ~n189 & ~n195 ;
  assign n197 = n187 & ~n196 ;
  assign n198 = n70 & n197 ;
  assign n176 = x3 & ~x5 ;
  assign n175 = x4 ^ x3 ;
  assign n177 = n176 ^ n175 ;
  assign n178 = n177 ^ x4 ;
  assign n199 = n198 ^ n178 ;
  assign n203 = n199 ^ n177 ;
  assign n204 = n203 ^ n175 ;
  assign n179 = n178 ^ n177 ;
  assign n180 = n179 ^ n175 ;
  assign n181 = n180 ^ n175 ;
  assign n182 = x2 & x11 ;
  assign n183 = n44 & n182 ;
  assign n184 = n183 ^ n177 ;
  assign n185 = n184 ^ n175 ;
  assign n186 = ~n181 & n185 ;
  assign n200 = n199 ^ n186 ;
  assign n201 = n200 ^ n175 ;
  assign n202 = n180 & n201 ;
  assign n205 = n204 ^ n202 ;
  assign n206 = n205 ^ n180 ;
  assign n207 = n175 ^ x1 ;
  assign n208 = n204 ^ n201 ;
  assign n209 = n208 ^ n180 ;
  assign n210 = ~n207 & n209 ;
  assign n211 = n210 ^ n175 ;
  assign n212 = n206 & ~n211 ;
  assign n213 = n212 ^ n210 ;
  assign n214 = n213 ^ n175 ;
  assign n215 = n214 ^ x3 ;
  assign n216 = x0 & n215 ;
  assign n217 = ~x3 & ~x5 ;
  assign n218 = n198 & n217 ;
  assign n219 = ~x0 & x2 ;
  assign n220 = ~n176 & ~n219 ;
  assign n221 = x4 & ~n220 ;
  assign n222 = ~n218 & ~n221 ;
  assign n223 = x1 & ~n222 ;
  assign n224 = x1 & ~n193 ;
  assign n225 = n195 & ~n224 ;
  assign n226 = ~n188 & ~n225 ;
  assign n227 = x1 & ~x9 ;
  assign n228 = ~n53 & n70 ;
  assign n229 = ~n227 & n228 ;
  assign n230 = ~n226 & n229 ;
  assign n231 = x3 & ~n230 ;
  assign n232 = x2 & ~n193 ;
  assign n233 = ~x1 & x3 ;
  assign n234 = x9 & n233 ;
  assign n235 = ~x2 & ~x5 ;
  assign n236 = ~x0 & n235 ;
  assign n237 = ~n234 & ~n236 ;
  assign n238 = ~x4 & ~n237 ;
  assign n239 = ~n232 & n238 ;
  assign n240 = ~n231 & n239 ;
  assign n241 = ~n223 & ~n240 ;
  assign n242 = ~n216 & n241 ;
  assign n243 = ~n174 & n242 ;
  assign n244 = n243 ^ x18 ;
  assign n245 = n40 & n244 ;
  assign n246 = n245 ^ x18 ;
  assign n247 = x14 & n246 ;
  assign n248 = ~n37 & n247 ;
  assign y0 = ~n248 ;
endmodule
