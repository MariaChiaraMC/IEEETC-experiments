module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 ;
  assign n11 = ~x5 & ~x7 ;
  assign n12 = x8 & ~x9 ;
  assign n13 = x2 & x3 ;
  assign n14 = n12 & n13 ;
  assign n15 = n11 & n14 ;
  assign n16 = x5 & x8 ;
  assign n17 = x7 & ~x9 ;
  assign n18 = x2 & n17 ;
  assign n19 = ~x3 & ~x6 ;
  assign n20 = n18 & n19 ;
  assign n21 = ~x2 & x6 ;
  assign n22 = ~x1 & ~x9 ;
  assign n23 = n21 & ~n22 ;
  assign n24 = n17 ^ x3 ;
  assign n25 = n23 & n24 ;
  assign n26 = ~n20 & ~n25 ;
  assign n27 = n16 & ~n26 ;
  assign n28 = ~n15 & ~n27 ;
  assign n29 = x4 & ~n28 ;
  assign n30 = x0 & n29 ;
  assign n31 = n16 & n18 ;
  assign n32 = x3 & x6 ;
  assign n33 = n32 ^ n19 ;
  assign n34 = x0 & n33 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = n31 & n35 ;
  assign n37 = x3 & x5 ;
  assign n38 = x2 & ~x3 ;
  assign n39 = n11 & n38 ;
  assign n40 = ~n37 & ~n39 ;
  assign n41 = ~x0 & ~x8 ;
  assign n42 = x9 & n41 ;
  assign n43 = ~x6 & n42 ;
  assign n44 = ~n40 & n43 ;
  assign n45 = ~x0 & x7 ;
  assign n46 = ~x8 & ~x9 ;
  assign n47 = ~x5 & n46 ;
  assign n48 = x9 & n16 ;
  assign n49 = ~n47 & ~n48 ;
  assign n50 = n49 ^ x3 ;
  assign n57 = n50 ^ n49 ;
  assign n51 = n50 ^ x5 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = x6 ^ x5 ;
  assign n54 = n53 ^ x5 ;
  assign n55 = n54 ^ n52 ;
  assign n56 = n52 & ~n55 ;
  assign n58 = n57 ^ n56 ;
  assign n59 = n58 ^ n52 ;
  assign n60 = n49 ^ n12 ;
  assign n61 = n56 ^ n52 ;
  assign n62 = ~n60 & n61 ;
  assign n63 = n62 ^ n49 ;
  assign n64 = n59 & ~n63 ;
  assign n65 = n64 ^ n49 ;
  assign n66 = n65 ^ n49 ;
  assign n67 = n45 & n66 ;
  assign n68 = ~x5 & ~x6 ;
  assign n69 = ~x8 & x9 ;
  assign n70 = x3 & n69 ;
  assign n71 = n68 & n70 ;
  assign n72 = x5 & n32 ;
  assign n73 = x9 & n72 ;
  assign n74 = ~x3 & x5 ;
  assign n75 = ~x6 & n46 ;
  assign n76 = n74 & n75 ;
  assign n77 = n32 & n47 ;
  assign n78 = ~n76 & ~n77 ;
  assign n79 = ~n73 & n78 ;
  assign n80 = ~x7 & ~n79 ;
  assign n81 = ~n71 & ~n80 ;
  assign n82 = n81 ^ x0 ;
  assign n83 = n82 ^ n81 ;
  assign n84 = n83 ^ n67 ;
  assign n85 = ~x6 & ~x7 ;
  assign n86 = x3 & ~n47 ;
  assign n87 = ~n49 & ~n86 ;
  assign n88 = n87 ^ n85 ;
  assign n89 = n85 & n88 ;
  assign n90 = n89 ^ n81 ;
  assign n91 = n90 ^ n85 ;
  assign n92 = n84 & ~n91 ;
  assign n93 = n92 ^ n89 ;
  assign n94 = n93 ^ n85 ;
  assign n95 = ~n67 & n94 ;
  assign n96 = n95 ^ n67 ;
  assign n97 = ~x2 & n96 ;
  assign n98 = x7 & n68 ;
  assign n99 = ~x2 & x3 ;
  assign n100 = n98 & n99 ;
  assign n101 = n12 & n100 ;
  assign n102 = ~n97 & ~n101 ;
  assign n103 = ~n44 & n102 ;
  assign n104 = n103 ^ x4 ;
  assign n105 = n104 ^ n103 ;
  assign n106 = n37 & n85 ;
  assign n107 = x0 & x2 ;
  assign n108 = n106 & n107 ;
  assign n109 = n69 & n108 ;
  assign n110 = x6 & x7 ;
  assign n111 = ~x0 & n110 ;
  assign n112 = x9 & n111 ;
  assign n113 = x5 ^ x3 ;
  assign n114 = ~x8 & n113 ;
  assign n115 = n114 ^ x3 ;
  assign n116 = n112 & n115 ;
  assign n117 = x0 & n11 ;
  assign n118 = n12 & n32 ;
  assign n119 = n117 & n118 ;
  assign n120 = n45 & n74 ;
  assign n121 = x0 & ~x3 ;
  assign n122 = ~x5 & n121 ;
  assign n123 = ~n120 & ~n122 ;
  assign n124 = n75 & ~n123 ;
  assign n125 = ~n119 & ~n124 ;
  assign n126 = ~n116 & n125 ;
  assign n127 = ~x2 & ~n126 ;
  assign n128 = x2 & x5 ;
  assign n129 = n128 ^ x7 ;
  assign n130 = n129 ^ n118 ;
  assign n131 = n130 ^ n128 ;
  assign n132 = n131 ^ n130 ;
  assign n133 = n130 ^ n71 ;
  assign n134 = n133 ^ n129 ;
  assign n135 = n132 & ~n134 ;
  assign n136 = n135 ^ n71 ;
  assign n137 = x6 & x9 ;
  assign n138 = ~x3 & ~x8 ;
  assign n139 = n137 & n138 ;
  assign n140 = ~n71 & ~n139 ;
  assign n141 = n140 ^ n129 ;
  assign n142 = ~n136 & n141 ;
  assign n143 = n142 ^ n140 ;
  assign n144 = n129 & n143 ;
  assign n145 = n144 ^ n135 ;
  assign n146 = n145 ^ x7 ;
  assign n147 = n146 ^ n71 ;
  assign n148 = ~x0 & n147 ;
  assign n149 = ~n127 & ~n148 ;
  assign n150 = ~n109 & n149 ;
  assign n151 = n150 ^ n103 ;
  assign n152 = ~n105 & n151 ;
  assign n153 = n152 ^ n103 ;
  assign n154 = ~n36 & n153 ;
  assign n155 = n154 ^ x1 ;
  assign n156 = n155 ^ n154 ;
  assign n157 = n14 & n117 ;
  assign n158 = n13 & n98 ;
  assign n159 = ~x5 & n33 ;
  assign n160 = n159 ^ n32 ;
  assign n161 = ~x2 & n160 ;
  assign n162 = ~n158 & ~n161 ;
  assign n163 = ~x0 & n12 ;
  assign n164 = ~n162 & n163 ;
  assign n165 = ~x0 & ~n32 ;
  assign n166 = ~x3 & x7 ;
  assign n167 = n128 & ~n166 ;
  assign n168 = ~n85 & n167 ;
  assign n169 = n165 & n168 ;
  assign n170 = n32 & n117 ;
  assign n171 = n74 & n110 ;
  assign n172 = n107 & n171 ;
  assign n173 = ~n108 & ~n172 ;
  assign n174 = ~n170 & n173 ;
  assign n175 = ~n169 & n174 ;
  assign n176 = n46 & ~n175 ;
  assign n185 = ~x2 & ~x8 ;
  assign n186 = ~n107 & ~n185 ;
  assign n187 = ~x5 & x9 ;
  assign n188 = n85 & n187 ;
  assign n189 = ~n186 & n188 ;
  assign n177 = x6 & x8 ;
  assign n178 = n177 ^ x2 ;
  assign n179 = n178 ^ n177 ;
  assign n180 = ~x6 & ~x8 ;
  assign n181 = n180 ^ n177 ;
  assign n182 = ~n179 & n181 ;
  assign n183 = n182 ^ n177 ;
  assign n184 = n117 & n183 ;
  assign n190 = n189 ^ n184 ;
  assign n191 = n190 ^ n189 ;
  assign n192 = ~n21 & n45 ;
  assign n193 = n48 & n192 ;
  assign n194 = n193 ^ n189 ;
  assign n195 = n194 ^ n189 ;
  assign n196 = ~n191 & ~n195 ;
  assign n197 = n196 ^ n189 ;
  assign n198 = x3 & ~n197 ;
  assign n199 = n198 ^ n189 ;
  assign n200 = ~n176 & ~n199 ;
  assign n201 = ~n164 & n200 ;
  assign n202 = n201 ^ x4 ;
  assign n203 = n202 ^ n201 ;
  assign n210 = x8 ^ x3 ;
  assign n204 = x7 ^ x6 ;
  assign n205 = n204 ^ x8 ;
  assign n206 = n205 ^ x8 ;
  assign n207 = n206 ^ x0 ;
  assign n208 = n207 ^ x0 ;
  assign n209 = n208 ^ n205 ;
  assign n211 = n210 ^ n209 ;
  assign n212 = n211 ^ x0 ;
  assign n213 = n212 ^ n210 ;
  assign n214 = n213 ^ n211 ;
  assign n215 = x7 ^ x2 ;
  assign n216 = n215 ^ x2 ;
  assign n217 = n216 ^ n215 ;
  assign n218 = n217 ^ n212 ;
  assign n219 = n218 ^ n211 ;
  assign n220 = ~n214 & n219 ;
  assign n221 = n220 ^ n212 ;
  assign n222 = n221 ^ n211 ;
  assign n223 = n217 ^ n211 ;
  assign n224 = n210 ^ n205 ;
  assign n225 = n224 ^ n217 ;
  assign n226 = n225 ^ n211 ;
  assign n227 = ~n223 & n226 ;
  assign n228 = n227 ^ n205 ;
  assign n229 = n228 ^ n210 ;
  assign n230 = n229 ^ n212 ;
  assign n231 = n230 ^ n217 ;
  assign n232 = n231 ^ n211 ;
  assign n233 = n216 ^ n205 ;
  assign n234 = n233 ^ n210 ;
  assign n235 = n234 ^ n212 ;
  assign n236 = n235 ^ n217 ;
  assign n237 = ~n211 & n236 ;
  assign n238 = n237 ^ n216 ;
  assign n239 = n238 ^ n205 ;
  assign n240 = n239 ^ n217 ;
  assign n241 = n240 ^ n211 ;
  assign n242 = ~n232 & ~n241 ;
  assign n243 = n242 ^ n205 ;
  assign n244 = n222 & n243 ;
  assign n245 = ~x5 & ~n244 ;
  assign n246 = n41 & n110 ;
  assign n247 = x0 & ~x7 ;
  assign n248 = x8 ^ x6 ;
  assign n249 = n247 & ~n248 ;
  assign n250 = ~n246 & ~n249 ;
  assign n251 = n38 & ~n250 ;
  assign n252 = ~x0 & n85 ;
  assign n253 = x8 & n99 ;
  assign n254 = n252 & n253 ;
  assign n255 = x5 & ~n254 ;
  assign n256 = n19 & n185 ;
  assign n257 = ~x0 & n256 ;
  assign n258 = n255 & ~n257 ;
  assign n259 = ~n251 & n258 ;
  assign n260 = ~x9 & ~n259 ;
  assign n261 = ~n245 & n260 ;
  assign n262 = ~x7 & n13 ;
  assign n263 = n41 & n262 ;
  assign n264 = n120 & n185 ;
  assign n265 = ~x8 & n38 ;
  assign n266 = ~n37 & ~n265 ;
  assign n267 = x5 & ~x8 ;
  assign n268 = x0 & ~n267 ;
  assign n269 = ~n266 & n268 ;
  assign n270 = x7 & n269 ;
  assign n271 = ~n264 & ~n270 ;
  assign n272 = ~n263 & n271 ;
  assign n273 = n137 & ~n272 ;
  assign n274 = x0 & ~n166 ;
  assign n275 = x9 & n68 ;
  assign n276 = n275 ^ x2 ;
  assign n277 = n276 ^ n275 ;
  assign n278 = n275 ^ n106 ;
  assign n279 = n278 ^ n275 ;
  assign n280 = ~n277 & n279 ;
  assign n281 = n280 ^ n275 ;
  assign n282 = ~x8 & n281 ;
  assign n283 = n282 ^ n275 ;
  assign n284 = n274 & n283 ;
  assign n285 = ~n13 & n284 ;
  assign n286 = ~n273 & ~n285 ;
  assign n287 = ~n261 & n286 ;
  assign n288 = n287 ^ n201 ;
  assign n289 = n203 & n288 ;
  assign n290 = n289 ^ n201 ;
  assign n291 = ~n157 & n290 ;
  assign n292 = n291 ^ n154 ;
  assign n293 = ~n156 & n292 ;
  assign n294 = n293 ^ n154 ;
  assign n295 = ~n30 & n294 ;
  assign y0 = ~n295 ;
endmodule
