module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 ;
  assign n9 = x2 & x3 ;
  assign n10 = x1 & ~x4 ;
  assign n11 = ~n9 & ~n10 ;
  assign n12 = x6 & x7 ;
  assign n13 = ~x5 & n12 ;
  assign n14 = ~n11 & n13 ;
  assign n15 = x5 & ~x6 ;
  assign n16 = ~x3 & ~x7 ;
  assign n17 = n16 ^ x1 ;
  assign n18 = x2 & ~n17 ;
  assign n19 = n18 ^ x1 ;
  assign n20 = n15 & ~n19 ;
  assign n21 = ~x6 & ~x7 ;
  assign n22 = x3 & ~n21 ;
  assign n23 = ~x2 & ~x6 ;
  assign n24 = ~n21 & ~n23 ;
  assign n25 = ~n22 & ~n24 ;
  assign n26 = x2 & x6 ;
  assign n27 = ~n16 & n26 ;
  assign n28 = ~x1 & ~n27 ;
  assign n29 = ~n25 & ~n28 ;
  assign n30 = x5 & ~n29 ;
  assign n31 = ~x4 & n30 ;
  assign n32 = ~n20 & ~n31 ;
  assign n33 = ~n14 & n32 ;
  assign n34 = x0 & ~n33 ;
  assign n35 = ~x5 & ~n26 ;
  assign n36 = n22 & ~n35 ;
  assign n37 = x2 & n12 ;
  assign n38 = x2 & x5 ;
  assign n39 = ~n37 & ~n38 ;
  assign n40 = ~x0 & n39 ;
  assign n41 = ~n36 & n40 ;
  assign n42 = n16 ^ x5 ;
  assign n43 = x6 & ~n42 ;
  assign n44 = n43 ^ x5 ;
  assign n45 = ~x2 & ~n44 ;
  assign n46 = ~n41 & ~n45 ;
  assign n47 = x1 & ~n46 ;
  assign n50 = x3 & x7 ;
  assign n48 = x5 ^ x2 ;
  assign n49 = n48 ^ x6 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = n51 ^ x5 ;
  assign n54 = n52 ^ x1 ;
  assign n53 = n52 ^ n50 ;
  assign n55 = n54 ^ n53 ;
  assign n56 = n55 ^ n48 ;
  assign n63 = n56 ^ n54 ;
  assign n64 = n63 ^ n48 ;
  assign n57 = n56 ^ n52 ;
  assign n58 = n57 ^ n51 ;
  assign n65 = n64 ^ n58 ;
  assign n66 = n65 ^ n51 ;
  assign n67 = ~n51 & n66 ;
  assign n68 = n67 ^ n56 ;
  assign n69 = n68 ^ n58 ;
  assign n70 = n69 ^ n51 ;
  assign n71 = n70 ^ n48 ;
  assign n72 = n58 ^ n51 ;
  assign n73 = n72 ^ n48 ;
  assign n74 = ~n69 & n73 ;
  assign n75 = n74 ^ n56 ;
  assign n76 = n75 ^ n58 ;
  assign n77 = n76 ^ n51 ;
  assign n78 = n77 ^ n48 ;
  assign n79 = ~n71 & ~n78 ;
  assign n59 = n58 ^ n56 ;
  assign n60 = n59 ^ n51 ;
  assign n61 = n60 ^ n48 ;
  assign n62 = n60 & ~n61 ;
  assign n80 = n79 ^ n62 ;
  assign n81 = n80 ^ n67 ;
  assign n82 = n81 ^ n56 ;
  assign n83 = n82 ^ n58 ;
  assign n84 = n83 ^ n51 ;
  assign n85 = n84 ^ n48 ;
  assign n86 = x0 & ~n85 ;
  assign n87 = x1 & ~x6 ;
  assign n88 = n9 & ~n87 ;
  assign n89 = n12 ^ x5 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = x1 ^ x0 ;
  assign n92 = x5 & ~n91 ;
  assign n93 = n92 ^ x1 ;
  assign n94 = n90 & ~n93 ;
  assign n95 = n94 ^ n92 ;
  assign n96 = n95 ^ x1 ;
  assign n97 = n96 ^ x5 ;
  assign n98 = n88 & ~n97 ;
  assign n99 = ~n86 & ~n98 ;
  assign n100 = ~n47 & n99 ;
  assign n103 = n100 ^ x1 ;
  assign n104 = n103 ^ n100 ;
  assign n101 = n100 ^ x5 ;
  assign n102 = n101 ^ n100 ;
  assign n105 = n104 ^ n102 ;
  assign n106 = ~n23 & n50 ;
  assign n107 = ~n26 & ~n106 ;
  assign n108 = ~x0 & ~n107 ;
  assign n109 = ~n37 & ~n108 ;
  assign n110 = n109 ^ n100 ;
  assign n111 = n110 ^ n100 ;
  assign n112 = n111 ^ n104 ;
  assign n113 = n104 & ~n112 ;
  assign n114 = n113 ^ n104 ;
  assign n115 = n105 & n114 ;
  assign n116 = n115 ^ n113 ;
  assign n117 = n116 ^ n100 ;
  assign n118 = n117 ^ n104 ;
  assign n119 = ~x4 & ~n118 ;
  assign n120 = n119 ^ n100 ;
  assign n121 = ~n34 & n120 ;
  assign y0 = ~n121 ;
endmodule
