module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 ;
  assign n9 = x2 ^ x1 ;
  assign n10 = x6 ^ x3 ;
  assign n11 = x5 ^ x3 ;
  assign n12 = ~n10 & ~n11 ;
  assign n13 = n12 ^ x3 ;
  assign n14 = ~x3 & x7 ;
  assign n15 = n14 ^ x4 ;
  assign n16 = ~n13 & ~n15 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = ~x4 & n17 ;
  assign n19 = n18 ^ x3 ;
  assign n20 = n19 ^ x4 ;
  assign n21 = ~x2 & ~n20 ;
  assign n22 = ~n9 & n21 ;
  assign n23 = n22 ^ n9 ;
  assign y0 = n23 ;
endmodule
