// Benchmark "./b12.pla" written by ABC on Thu Apr 23 10:59:48 2020

module \./b12.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    z1  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14;
  output z1;
  wire new_n17_, new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_;
  assign new_n17_ = x5 & x6;
  assign new_n18_ = x2 & new_n17_;
  assign new_n19_ = x1 & new_n18_;
  assign new_n20_ = x1 & x3;
  assign new_n21_ = ~x2 & ~new_n20_;
  assign new_n22_ = ~x3 & ~x4;
  assign new_n23_ = ~new_n21_ & ~new_n22_;
  assign z1 = ~new_n19_ & new_n23_;
endmodule


