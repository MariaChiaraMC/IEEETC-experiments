module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 ;
  assign n9 = ~x6 & x7 ;
  assign n10 = x3 & x4 ;
  assign n11 = ~x2 & x5 ;
  assign n12 = n10 & n11 ;
  assign n13 = n9 & n12 ;
  assign n14 = x0 & n13 ;
  assign n15 = ~x2 & ~x3 ;
  assign n16 = ~n11 & ~n15 ;
  assign n17 = ~x0 & x7 ;
  assign n18 = n16 & n17 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = ~x3 & x5 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = ~x3 & ~x6 ;
  assign n25 = x5 & ~x7 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n24 & n26 ;
  assign n28 = n27 ^ n20 ;
  assign n29 = n28 ^ n24 ;
  assign n30 = n23 & ~n29 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = ~n19 & n32 ;
  assign n34 = n33 ^ n18 ;
  assign n35 = x4 & n34 ;
  assign n36 = x2 & ~x3 ;
  assign n37 = x4 & ~x5 ;
  assign n38 = x6 & ~x7 ;
  assign n39 = n37 & n38 ;
  assign n40 = n36 & n39 ;
  assign n43 = ~x5 & x7 ;
  assign n41 = ~x4 & ~n38 ;
  assign n42 = ~n16 & n41 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = n42 ^ x3 ;
  assign n46 = n45 ^ n44 ;
  assign n47 = ~x4 & x6 ;
  assign n48 = n47 ^ n9 ;
  assign n49 = x3 & ~n48 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = ~n46 & ~n50 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = n52 ^ n47 ;
  assign n54 = n53 ^ x3 ;
  assign n55 = n44 & ~n54 ;
  assign n56 = n55 ^ n43 ;
  assign n57 = ~n40 & ~n56 ;
  assign n58 = x3 & ~x6 ;
  assign n59 = x2 & n58 ;
  assign n60 = x7 ^ x4 ;
  assign n61 = x7 ^ x5 ;
  assign n62 = n60 & n61 ;
  assign n63 = n59 & n62 ;
  assign n64 = n57 & ~n63 ;
  assign n65 = n64 ^ x0 ;
  assign n66 = n65 ^ n64 ;
  assign n67 = n66 ^ n35 ;
  assign n68 = ~x3 & n47 ;
  assign n69 = ~x7 & n68 ;
  assign n70 = x2 & x7 ;
  assign n71 = ~n10 & n70 ;
  assign n72 = x6 ^ x3 ;
  assign n73 = n71 & n72 ;
  assign n74 = ~n69 & ~n73 ;
  assign n75 = n74 ^ x5 ;
  assign n76 = x5 & ~n75 ;
  assign n77 = n76 ^ n64 ;
  assign n78 = n77 ^ x5 ;
  assign n79 = n67 & ~n78 ;
  assign n80 = n79 ^ n76 ;
  assign n81 = n80 ^ x5 ;
  assign n82 = ~n35 & n81 ;
  assign n83 = n82 ^ n35 ;
  assign n84 = n83 ^ x1 ;
  assign n85 = n84 ^ n83 ;
  assign n86 = x5 ^ x2 ;
  assign n87 = n24 ^ x0 ;
  assign n88 = n87 ^ n86 ;
  assign n89 = x3 & x6 ;
  assign n90 = n89 ^ x5 ;
  assign n91 = ~x0 & ~n90 ;
  assign n92 = n91 ^ x5 ;
  assign n93 = n88 & n92 ;
  assign n94 = n93 ^ n91 ;
  assign n95 = n94 ^ x5 ;
  assign n96 = n95 ^ x0 ;
  assign n97 = ~n86 & ~n96 ;
  assign n98 = n97 ^ x4 ;
  assign n99 = n98 ^ n97 ;
  assign n100 = ~x0 & x5 ;
  assign n101 = ~x2 & n24 ;
  assign n102 = n100 & n101 ;
  assign n103 = n102 ^ n97 ;
  assign n104 = ~n99 & n103 ;
  assign n105 = n104 ^ n97 ;
  assign n106 = ~x7 & n105 ;
  assign n107 = ~n47 & ~n70 ;
  assign n108 = x7 ^ x2 ;
  assign n109 = x4 ^ x2 ;
  assign n110 = n109 ^ x3 ;
  assign n111 = n110 ^ x2 ;
  assign n112 = n108 & ~n111 ;
  assign n113 = n112 ^ x2 ;
  assign n114 = n107 ^ n36 ;
  assign n115 = n113 & n114 ;
  assign n116 = n115 ^ n36 ;
  assign n117 = n107 & n116 ;
  assign n118 = n117 ^ n107 ;
  assign n119 = n118 ^ n107 ;
  assign n120 = x5 & n119 ;
  assign n121 = n37 ^ x6 ;
  assign n122 = n36 ^ x7 ;
  assign n123 = n122 ^ n36 ;
  assign n124 = n36 ^ x3 ;
  assign n125 = ~n123 & n124 ;
  assign n126 = n125 ^ n36 ;
  assign n127 = n126 ^ n37 ;
  assign n128 = ~n121 & n127 ;
  assign n129 = n128 ^ n125 ;
  assign n130 = n129 ^ n36 ;
  assign n131 = n130 ^ x6 ;
  assign n132 = n37 & ~n131 ;
  assign n133 = n132 ^ n37 ;
  assign n134 = ~n120 & ~n133 ;
  assign n135 = n134 ^ x0 ;
  assign n136 = n135 ^ n134 ;
  assign n137 = n136 ^ n106 ;
  assign n138 = ~x5 & x6 ;
  assign n139 = n138 ^ x2 ;
  assign n140 = n139 ^ x4 ;
  assign n141 = n58 ^ x3 ;
  assign n142 = ~x2 & ~n141 ;
  assign n143 = n142 ^ x3 ;
  assign n144 = n140 & n143 ;
  assign n145 = n144 ^ n142 ;
  assign n146 = n145 ^ x3 ;
  assign n147 = n146 ^ x2 ;
  assign n148 = ~x4 & ~n147 ;
  assign n149 = n148 ^ x7 ;
  assign n150 = x7 & n149 ;
  assign n151 = n150 ^ n134 ;
  assign n152 = n151 ^ x7 ;
  assign n153 = n137 & ~n152 ;
  assign n154 = n153 ^ n150 ;
  assign n155 = n154 ^ x7 ;
  assign n156 = ~n106 & n155 ;
  assign n157 = n156 ^ n106 ;
  assign n158 = n157 ^ n83 ;
  assign n159 = n85 & n158 ;
  assign n160 = n159 ^ n83 ;
  assign n161 = ~n14 & ~n160 ;
  assign y0 = ~n161 ;
endmodule
