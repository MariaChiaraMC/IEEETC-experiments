// Benchmark "./pla/amd.pla_20" written by ABC on Mon Apr 20 15:43:51 2020

module \./pla/amd.pla_20  ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    z0  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13;
  output z0;
  wire new_n16_, new_n17_, new_n18_, new_n19_, new_n20_, new_n21_, new_n22_,
    new_n23_, new_n24_, new_n25_;
  assign new_n16_ = x03 & ~x10;
  assign new_n17_ = ~x11 & ~new_n16_;
  assign new_n18_ = ~x05 & ~x13;
  assign new_n19_ = ~x08 & new_n18_;
  assign new_n20_ = ~new_n17_ & new_n19_;
  assign new_n21_ = ~x06 & x10;
  assign new_n22_ = x11 & ~new_n21_;
  assign new_n23_ = ~x09 & ~x12;
  assign new_n24_ = ~x04 & new_n23_;
  assign new_n25_ = ~new_n22_ & new_n24_;
  assign z0 = new_n20_ & new_n25_;
endmodule


