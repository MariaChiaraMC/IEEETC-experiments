module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 ;
  output y0 ;
  wire n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 ;
  assign n14 = ~x3 & ~x5 ;
  assign n15 = x1 & n14 ;
  assign n16 = x3 & x5 ;
  assign n17 = x4 & ~n16 ;
  assign n18 = ~n15 & ~n17 ;
  assign n19 = ~x2 & ~n18 ;
  assign n21 = x4 ^ x3 ;
  assign n20 = x4 ^ x1 ;
  assign n22 = n21 ^ n20 ;
  assign n25 = x6 ^ x1 ;
  assign n23 = x6 ^ x5 ;
  assign n24 = n23 ^ n21 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n25 ^ n20 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = n28 ^ x6 ;
  assign n30 = n29 ^ n22 ;
  assign n31 = n26 & n30 ;
  assign n32 = n31 ^ n21 ;
  assign n33 = n22 & ~n32 ;
  assign n34 = n33 ^ n21 ;
  assign n35 = x6 ^ x2 ;
  assign n36 = n31 ^ n26 ;
  assign n37 = ~n35 & n36 ;
  assign n38 = n37 ^ x6 ;
  assign n39 = ~n34 & n38 ;
  assign n40 = n39 ^ x4 ;
  assign n41 = ~n19 & ~n40 ;
  assign n42 = ~n14 & ~n16 ;
  assign n43 = n42 ^ x1 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = ~x6 & ~n42 ;
  assign n46 = ~x7 & ~x11 ;
  assign n47 = x8 & ~x10 ;
  assign n48 = ~x9 & ~x12 ;
  assign n49 = n16 & n48 ;
  assign n50 = n47 & n49 ;
  assign n51 = n46 & n50 ;
  assign n52 = x4 & ~n51 ;
  assign n53 = ~n45 & ~n52 ;
  assign n54 = n53 ^ n42 ;
  assign n55 = n44 & ~n54 ;
  assign n56 = n55 ^ n42 ;
  assign n57 = x2 & ~n56 ;
  assign n58 = n41 & ~n57 ;
  assign n59 = ~x0 & ~n58 ;
  assign y0 = n59 ;
endmodule
