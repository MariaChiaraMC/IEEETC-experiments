module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 ;
  assign n25 = x1 & x2 ;
  assign n26 = x5 & n25 ;
  assign n27 = ~x0 & n26 ;
  assign n28 = n27 ^ x4 ;
  assign n29 = ~x3 & ~x14 ;
  assign n30 = x3 & x14 ;
  assign n31 = ~n29 & ~n30 ;
  assign n32 = x15 & x16 ;
  assign n33 = ~x18 & x23 ;
  assign n34 = n32 & n33 ;
  assign n35 = ~n31 & n34 ;
  assign n36 = x6 ^ x3 ;
  assign n37 = n36 ^ x6 ;
  assign n38 = x7 ^ x6 ;
  assign n39 = n37 & n38 ;
  assign n40 = n39 ^ x6 ;
  assign n41 = x17 & n40 ;
  assign n42 = ~n35 & ~n41 ;
  assign n43 = n42 ^ n28 ;
  assign n44 = n43 ^ n27 ;
  assign n45 = n44 ^ n43 ;
  assign n46 = ~x17 & x18 ;
  assign n47 = ~n25 & n32 ;
  assign n48 = ~n46 & n47 ;
  assign n58 = ~x1 & ~x2 ;
  assign n49 = x2 ^ x1 ;
  assign n50 = n49 ^ x2 ;
  assign n51 = x11 ^ x2 ;
  assign n52 = n51 ^ x2 ;
  assign n53 = n50 & n52 ;
  assign n54 = n53 ^ x2 ;
  assign n55 = x14 & n54 ;
  assign n56 = n55 ^ x2 ;
  assign n57 = x10 & n56 ;
  assign n59 = n58 ^ n57 ;
  assign n60 = n59 ^ x0 ;
  assign n68 = n60 ^ n59 ;
  assign n61 = ~x9 & n30 ;
  assign n62 = n61 ^ n60 ;
  assign n63 = n62 ^ n59 ;
  assign n64 = n60 ^ n57 ;
  assign n65 = n64 ^ n61 ;
  assign n66 = n65 ^ n63 ;
  assign n67 = n63 & ~n66 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = n69 ^ n63 ;
  assign n71 = n59 ^ n29 ;
  assign n72 = n67 ^ n63 ;
  assign n73 = ~n71 & n72 ;
  assign n74 = n73 ^ n59 ;
  assign n75 = ~n70 & n74 ;
  assign n76 = n75 ^ n59 ;
  assign n77 = n76 ^ n58 ;
  assign n78 = n77 ^ n59 ;
  assign n79 = n48 & n78 ;
  assign n80 = ~x5 & n79 ;
  assign n81 = n80 ^ n43 ;
  assign n82 = n81 ^ n28 ;
  assign n83 = n45 & n82 ;
  assign n84 = n83 ^ n80 ;
  assign n85 = x14 & x18 ;
  assign n86 = n32 & ~n85 ;
  assign n87 = ~n31 & n86 ;
  assign n88 = x14 ^ x3 ;
  assign n89 = x15 ^ x14 ;
  assign n90 = ~n88 & n89 ;
  assign n91 = n90 ^ x14 ;
  assign n92 = x16 & n91 ;
  assign n93 = x17 & ~n92 ;
  assign n94 = ~n87 & ~n93 ;
  assign n95 = ~n80 & n94 ;
  assign n96 = n95 ^ n28 ;
  assign n97 = ~n84 & ~n96 ;
  assign n98 = n97 ^ n95 ;
  assign n99 = ~n28 & n98 ;
  assign n100 = n99 ^ n83 ;
  assign n101 = n100 ^ x4 ;
  assign n102 = n101 ^ n80 ;
  assign n103 = x13 & ~n102 ;
  assign y0 = n103 ;
endmodule
