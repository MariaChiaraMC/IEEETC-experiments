module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 ;
  assign n11 = ~x1 & ~x3 ;
  assign n12 = x2 & x4 ;
  assign n13 = ~x7 & x8 ;
  assign n14 = n12 & n13 ;
  assign n15 = x5 & ~x6 ;
  assign n16 = n14 & n15 ;
  assign n17 = n11 & n16 ;
  assign n18 = ~x2 & x6 ;
  assign n19 = x7 & n18 ;
  assign n20 = ~x1 & ~x4 ;
  assign n21 = x5 & ~x8 ;
  assign n22 = ~x0 & ~x3 ;
  assign n23 = n21 & ~n22 ;
  assign n24 = n20 & n23 ;
  assign n25 = n19 & n24 ;
  assign n26 = x9 & ~n25 ;
  assign n27 = ~n17 & n26 ;
  assign n28 = ~x2 & x4 ;
  assign n29 = ~x5 & n28 ;
  assign n30 = x1 & x3 ;
  assign n31 = x7 & x8 ;
  assign n32 = n30 & n31 ;
  assign n33 = n29 & n32 ;
  assign n34 = ~x1 & ~x5 ;
  assign n35 = x2 & ~x8 ;
  assign n36 = ~x4 & ~x7 ;
  assign n37 = x3 & ~n36 ;
  assign n38 = n35 & n37 ;
  assign n39 = n34 & n38 ;
  assign n40 = ~n33 & ~n39 ;
  assign n41 = n40 ^ x3 ;
  assign n43 = x2 & ~x4 ;
  assign n44 = x5 & x7 ;
  assign n45 = n43 & n44 ;
  assign n42 = ~x2 & ~x7 ;
  assign n46 = n45 ^ n42 ;
  assign n47 = n46 ^ x8 ;
  assign n54 = n47 ^ n46 ;
  assign n48 = n47 ^ n21 ;
  assign n49 = n48 ^ n46 ;
  assign n50 = n42 ^ n21 ;
  assign n51 = n50 ^ n21 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = n49 & n52 ;
  assign n55 = n54 ^ n53 ;
  assign n56 = n55 ^ n49 ;
  assign n57 = ~x4 & ~x5 ;
  assign n58 = n57 ^ n46 ;
  assign n59 = n53 ^ n49 ;
  assign n60 = ~n58 & n59 ;
  assign n61 = n60 ^ n46 ;
  assign n62 = ~n56 & n61 ;
  assign n63 = n62 ^ n46 ;
  assign n64 = n63 ^ n42 ;
  assign n65 = n64 ^ n46 ;
  assign n66 = n65 ^ x1 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = n35 & n36 ;
  assign n69 = x8 ^ x4 ;
  assign n70 = n69 ^ x4 ;
  assign n71 = n28 ^ x4 ;
  assign n72 = ~n70 & ~n71 ;
  assign n73 = n72 ^ x4 ;
  assign n74 = n44 & ~n73 ;
  assign n75 = ~n68 & ~n74 ;
  assign n76 = ~n14 & n75 ;
  assign n77 = n76 ^ n65 ;
  assign n78 = ~n67 & ~n77 ;
  assign n79 = n78 ^ n65 ;
  assign n80 = n79 ^ n40 ;
  assign n81 = ~n41 & n80 ;
  assign n82 = n81 ^ n78 ;
  assign n83 = n82 ^ n65 ;
  assign n84 = n83 ^ x3 ;
  assign n85 = n40 & ~n84 ;
  assign n86 = n85 ^ n40 ;
  assign n87 = n86 ^ n40 ;
  assign n88 = n87 ^ x6 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = n89 ^ x0 ;
  assign n91 = x2 & ~x3 ;
  assign n92 = x1 & x5 ;
  assign n93 = ~n34 & ~n92 ;
  assign n94 = ~x1 & ~x2 ;
  assign n95 = x4 & ~n94 ;
  assign n96 = n93 & n95 ;
  assign n97 = ~n91 & n96 ;
  assign n98 = x2 & ~x5 ;
  assign n99 = ~x4 & n11 ;
  assign n100 = ~n98 & n99 ;
  assign n101 = ~n97 & ~n100 ;
  assign n102 = n13 & ~n101 ;
  assign n103 = ~x3 & ~x8 ;
  assign n104 = n29 & n103 ;
  assign n105 = ~x1 & n104 ;
  assign n106 = n11 & n21 ;
  assign n107 = n12 & n106 ;
  assign n108 = n107 ^ x7 ;
  assign n109 = n108 ^ n107 ;
  assign n110 = n30 & n35 ;
  assign n111 = ~x1 & x8 ;
  assign n112 = x3 ^ x2 ;
  assign n113 = n111 & n112 ;
  assign n114 = ~n110 & ~n113 ;
  assign n115 = n57 & ~n114 ;
  assign n116 = n92 ^ x4 ;
  assign n117 = ~x2 & x3 ;
  assign n118 = n117 ^ n91 ;
  assign n119 = n91 ^ x8 ;
  assign n120 = n119 ^ n91 ;
  assign n121 = n118 & n120 ;
  assign n122 = n121 ^ n91 ;
  assign n123 = n122 ^ n92 ;
  assign n124 = n116 & n123 ;
  assign n125 = n124 ^ n121 ;
  assign n126 = n125 ^ n91 ;
  assign n127 = n126 ^ x4 ;
  assign n128 = n92 & n127 ;
  assign n129 = n128 ^ n92 ;
  assign n130 = ~n115 & ~n129 ;
  assign n131 = ~n104 & n130 ;
  assign n132 = n131 ^ n107 ;
  assign n133 = n109 & ~n132 ;
  assign n134 = n133 ^ n107 ;
  assign n135 = ~n105 & ~n134 ;
  assign n136 = n135 ^ n102 ;
  assign n137 = ~n102 & ~n136 ;
  assign n138 = n137 ^ n87 ;
  assign n139 = n138 ^ n102 ;
  assign n140 = ~n90 & ~n139 ;
  assign n141 = n140 ^ n137 ;
  assign n142 = n141 ^ n102 ;
  assign n143 = ~x0 & ~n142 ;
  assign n144 = n143 ^ x0 ;
  assign n145 = n27 & n144 ;
  assign n146 = x8 ^ x1 ;
  assign n147 = x7 ^ x2 ;
  assign n148 = n147 ^ n146 ;
  assign n149 = x7 ^ x6 ;
  assign n150 = n149 ^ x7 ;
  assign n151 = x8 ^ x7 ;
  assign n152 = n151 ^ x7 ;
  assign n153 = ~n150 & n152 ;
  assign n154 = n153 ^ x7 ;
  assign n155 = n154 ^ n146 ;
  assign n156 = ~n148 & ~n155 ;
  assign n157 = n156 ^ n153 ;
  assign n158 = n157 ^ x7 ;
  assign n159 = n158 ^ n147 ;
  assign n160 = ~n146 & n159 ;
  assign n161 = n160 ^ n146 ;
  assign n162 = n57 & ~n161 ;
  assign n166 = ~x2 & n44 ;
  assign n163 = x1 & x2 ;
  assign n164 = x6 & n163 ;
  assign n165 = n31 & n164 ;
  assign n167 = n166 ^ n165 ;
  assign n168 = n167 ^ n165 ;
  assign n169 = n111 ^ x8 ;
  assign n170 = ~x6 & ~n169 ;
  assign n171 = n170 ^ x8 ;
  assign n172 = n171 ^ n165 ;
  assign n173 = n172 ^ n165 ;
  assign n174 = n168 & ~n173 ;
  assign n175 = n174 ^ n165 ;
  assign n176 = ~x4 & n175 ;
  assign n177 = n176 ^ n165 ;
  assign n178 = ~n162 & ~n177 ;
  assign n179 = n178 ^ x3 ;
  assign n180 = n179 ^ n178 ;
  assign n181 = n180 ^ x0 ;
  assign n182 = x1 & x8 ;
  assign n183 = n29 & n182 ;
  assign n184 = ~x4 & n92 ;
  assign n185 = x6 ^ x2 ;
  assign n186 = n184 & ~n185 ;
  assign n187 = ~n183 & ~n186 ;
  assign n188 = x8 & n57 ;
  assign n189 = ~x6 & n188 ;
  assign n190 = ~n163 & n189 ;
  assign n191 = n187 & ~n190 ;
  assign n192 = x7 & ~n191 ;
  assign n193 = x4 & x5 ;
  assign n194 = x2 & x6 ;
  assign n195 = x4 & ~n194 ;
  assign n196 = ~n193 & ~n195 ;
  assign n197 = ~n164 & n196 ;
  assign n198 = ~x7 & ~n57 ;
  assign n199 = ~x1 & n185 ;
  assign n200 = n198 & ~n199 ;
  assign n201 = n197 & n200 ;
  assign n202 = ~x6 & n44 ;
  assign n203 = n163 & n202 ;
  assign n204 = x4 & n203 ;
  assign n205 = ~n201 & ~n204 ;
  assign n206 = ~x8 & ~n205 ;
  assign n207 = n206 ^ n192 ;
  assign n208 = ~n192 & n207 ;
  assign n209 = n208 ^ n178 ;
  assign n210 = n209 ^ n192 ;
  assign n211 = ~n181 & ~n210 ;
  assign n212 = n211 ^ n208 ;
  assign n213 = n212 ^ n192 ;
  assign n214 = x0 & ~n213 ;
  assign n215 = n214 ^ x0 ;
  assign n216 = n145 & ~n215 ;
  assign n217 = n30 & n57 ;
  assign n218 = x0 & x6 ;
  assign n219 = n42 & n218 ;
  assign n220 = n217 & n219 ;
  assign n221 = ~x9 & ~n220 ;
  assign n222 = x3 & ~n194 ;
  assign n223 = ~x0 & ~n222 ;
  assign n224 = n186 & n223 ;
  assign n225 = x0 & ~x6 ;
  assign n226 = ~x5 & n225 ;
  assign n227 = n43 & n226 ;
  assign n228 = n11 & n227 ;
  assign n229 = ~x2 & ~x3 ;
  assign n230 = ~x0 & ~x5 ;
  assign n231 = x6 & n230 ;
  assign n232 = n231 ^ x4 ;
  assign n233 = n232 ^ x1 ;
  assign n240 = n233 ^ n232 ;
  assign n235 = ~n93 & n225 ;
  assign n234 = n233 ^ n231 ;
  assign n236 = n235 ^ n234 ;
  assign n237 = n235 ^ n233 ;
  assign n238 = n237 ^ n232 ;
  assign n239 = n236 & ~n238 ;
  assign n241 = n240 ^ n239 ;
  assign n242 = x5 & x6 ;
  assign n243 = ~x0 & n242 ;
  assign n244 = n243 ^ n233 ;
  assign n245 = n240 & n244 ;
  assign n246 = n245 ^ n243 ;
  assign n247 = n241 & n246 ;
  assign n248 = n247 ^ n239 ;
  assign n249 = n248 ^ n233 ;
  assign n250 = n249 ^ x4 ;
  assign n251 = n250 ^ n232 ;
  assign n252 = n229 & n251 ;
  assign n253 = ~n228 & ~n252 ;
  assign n254 = ~n224 & n253 ;
  assign n255 = x7 & ~n254 ;
  assign n256 = ~x0 & n193 ;
  assign n257 = ~x6 & ~x7 ;
  assign n258 = n94 & n257 ;
  assign n259 = n256 & n258 ;
  assign n260 = n259 ^ x3 ;
  assign n261 = n19 & n230 ;
  assign n262 = ~x5 & ~x7 ;
  assign n263 = x2 & n262 ;
  assign n264 = ~n166 & ~n263 ;
  assign n265 = ~x4 & n225 ;
  assign n266 = ~n264 & n265 ;
  assign n267 = ~n261 & ~n266 ;
  assign n268 = n267 ^ x1 ;
  assign n269 = n268 ^ n267 ;
  assign n270 = x0 & ~x2 ;
  assign n271 = n262 & n270 ;
  assign n272 = ~n45 & ~n271 ;
  assign n273 = x6 & ~n272 ;
  assign n274 = ~x7 & n242 ;
  assign n275 = ~n226 & ~n274 ;
  assign n276 = x0 & ~x7 ;
  assign n277 = ~n28 & ~n276 ;
  assign n278 = ~n43 & n277 ;
  assign n279 = ~n275 & n278 ;
  assign n280 = ~n273 & ~n279 ;
  assign n281 = n280 ^ n267 ;
  assign n282 = n269 & n281 ;
  assign n283 = n282 ^ n267 ;
  assign n284 = n283 ^ n259 ;
  assign n285 = ~n260 & n284 ;
  assign n286 = n285 ^ n282 ;
  assign n287 = n286 ^ n267 ;
  assign n288 = n287 ^ x3 ;
  assign n289 = ~n259 & ~n288 ;
  assign n290 = n289 ^ n259 ;
  assign n291 = n290 ^ n259 ;
  assign n292 = ~n255 & n291 ;
  assign n293 = n292 ^ x8 ;
  assign n294 = n293 ^ n292 ;
  assign n295 = x4 ^ x2 ;
  assign n296 = n262 ^ x4 ;
  assign n297 = n296 ^ n262 ;
  assign n298 = n262 ^ n202 ;
  assign n299 = n297 & n298 ;
  assign n300 = n299 ^ n262 ;
  assign n301 = n295 & n300 ;
  assign n302 = ~x0 & n301 ;
  assign n303 = n43 & n274 ;
  assign n304 = ~n302 & ~n303 ;
  assign n305 = n30 & ~n304 ;
  assign n306 = x3 & ~x4 ;
  assign n307 = ~n218 & n262 ;
  assign n308 = n306 & n307 ;
  assign n309 = x4 ^ x3 ;
  assign n310 = ~n44 & ~n262 ;
  assign n311 = n310 ^ n309 ;
  assign n312 = x4 ^ x0 ;
  assign n313 = x5 ^ x4 ;
  assign n314 = n312 & n313 ;
  assign n315 = n314 ^ x4 ;
  assign n316 = n315 ^ n309 ;
  assign n317 = n311 & n316 ;
  assign n318 = n317 ^ n314 ;
  assign n319 = n318 ^ x4 ;
  assign n320 = n319 ^ n310 ;
  assign n321 = n309 & n320 ;
  assign n322 = n321 ^ n309 ;
  assign n323 = x6 & n322 ;
  assign n324 = ~n308 & ~n323 ;
  assign n325 = n94 & ~n324 ;
  assign n326 = ~x3 & x4 ;
  assign n327 = n274 & n326 ;
  assign n328 = n270 & n327 ;
  assign n329 = ~n325 & ~n328 ;
  assign n330 = ~n305 & n329 ;
  assign n331 = ~x0 & ~x1 ;
  assign n332 = n91 & n331 ;
  assign n333 = x6 & ~n310 ;
  assign n334 = n333 ^ x4 ;
  assign n335 = n334 ^ n333 ;
  assign n336 = n333 ^ n202 ;
  assign n337 = n335 & n336 ;
  assign n338 = n337 ^ n333 ;
  assign n339 = n332 & n338 ;
  assign n340 = n330 & ~n339 ;
  assign n341 = n340 ^ n292 ;
  assign n342 = n294 & n341 ;
  assign n343 = n342 ^ n292 ;
  assign n344 = n221 & n343 ;
  assign n345 = ~n216 & ~n344 ;
  assign n346 = ~x8 & n42 ;
  assign n347 = ~x1 & x3 ;
  assign n348 = n256 & n347 ;
  assign n349 = n348 ^ x0 ;
  assign n350 = n349 ^ n348 ;
  assign n351 = n11 & n193 ;
  assign n352 = ~n217 & ~n351 ;
  assign n353 = n352 ^ n348 ;
  assign n354 = n353 ^ n348 ;
  assign n355 = n350 & ~n354 ;
  assign n356 = n355 ^ n348 ;
  assign n357 = x6 & n356 ;
  assign n358 = n357 ^ n348 ;
  assign n359 = n346 & n358 ;
  assign n360 = ~n345 & ~n359 ;
  assign y0 = ~n360 ;
endmodule
