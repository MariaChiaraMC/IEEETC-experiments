module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 ;
  assign n11 = ~x3 & ~x4 ;
  assign n12 = x2 & ~n11 ;
  assign n13 = ~x1 & ~n12 ;
  assign n14 = ~x7 & ~n13 ;
  assign n15 = ~x6 & x8 ;
  assign n16 = x6 & ~x8 ;
  assign n17 = ~n15 & ~n16 ;
  assign n18 = ~n14 & n17 ;
  assign n19 = ~x5 & n18 ;
  assign n20 = ~x1 & x7 ;
  assign n21 = x4 ^ x0 ;
  assign n22 = x3 ^ x0 ;
  assign n23 = n21 & n22 ;
  assign n24 = n23 ^ x0 ;
  assign n25 = x2 ^ x0 ;
  assign n26 = n25 ^ x0 ;
  assign n27 = n26 ^ n20 ;
  assign n28 = n24 & n27 ;
  assign n29 = n28 ^ n23 ;
  assign n30 = n20 & n29 ;
  assign n31 = n30 ^ x0 ;
  assign n32 = n19 & n31 ;
  assign n48 = x1 & ~n11 ;
  assign n35 = x2 & ~x5 ;
  assign n34 = ~x2 & x5 ;
  assign n72 = n16 & ~n34 ;
  assign n73 = ~n35 & n72 ;
  assign n74 = ~x3 & ~n15 ;
  assign n75 = ~x3 & ~n34 ;
  assign n76 = ~n74 & ~n75 ;
  assign n77 = ~n73 & ~n76 ;
  assign n78 = n48 & ~n77 ;
  assign n79 = ~x1 & x2 ;
  assign n80 = x5 ^ x4 ;
  assign n63 = n16 ^ n15 ;
  assign n81 = n15 ^ x5 ;
  assign n82 = n81 ^ n15 ;
  assign n83 = n63 & n82 ;
  assign n84 = n83 ^ n15 ;
  assign n85 = n80 & n84 ;
  assign n86 = n79 & n85 ;
  assign n87 = ~n78 & ~n86 ;
  assign n88 = x6 ^ x4 ;
  assign n89 = n88 ^ x8 ;
  assign n90 = n34 ^ x8 ;
  assign n91 = n90 ^ x6 ;
  assign n92 = n91 ^ n34 ;
  assign n93 = n92 ^ n89 ;
  assign n94 = n35 ^ x6 ;
  assign n95 = n35 & ~n94 ;
  assign n96 = n95 ^ n34 ;
  assign n97 = n96 ^ n35 ;
  assign n98 = n93 & n97 ;
  assign n99 = n98 ^ n95 ;
  assign n100 = n99 ^ n35 ;
  assign n101 = n89 & n100 ;
  assign n102 = x1 & n101 ;
  assign n103 = x3 & ~n102 ;
  assign n104 = ~n87 & ~n103 ;
  assign n33 = x4 ^ x1 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = n35 ^ x4 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n37 & ~n39 ;
  assign n41 = n40 ^ n35 ;
  assign n42 = n33 & n41 ;
  assign n43 = n42 ^ n35 ;
  assign n44 = n17 ^ n15 ;
  assign n45 = x3 & n44 ;
  assign n46 = n45 ^ n15 ;
  assign n47 = n43 & n46 ;
  assign n49 = n16 ^ x2 ;
  assign n50 = n49 ^ x5 ;
  assign n51 = n50 ^ x1 ;
  assign n60 = n51 ^ n16 ;
  assign n52 = n16 ^ x5 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n53 ^ n51 ;
  assign n55 = n54 ^ n16 ;
  assign n56 = n53 ^ x1 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = ~n55 & n58 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = n61 ^ n55 ;
  assign n64 = n59 ^ n55 ;
  assign n65 = n63 & ~n64 ;
  assign n66 = n65 ^ n16 ;
  assign n67 = ~n62 & n66 ;
  assign n68 = n67 ^ n16 ;
  assign n69 = n68 ^ n16 ;
  assign n70 = ~n48 & n69 ;
  assign n71 = ~n47 & ~n70 ;
  assign n105 = n104 ^ n71 ;
  assign n106 = ~x7 & ~n105 ;
  assign n107 = n106 ^ n104 ;
  assign n108 = ~x0 & n107 ;
  assign n109 = ~n32 & ~n108 ;
  assign n110 = x9 & ~n109 ;
  assign y0 = n110 ;
endmodule
