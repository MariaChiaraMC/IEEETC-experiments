// Benchmark "./br1.pla" written by ABC on Thu Apr 23 10:59:48 2020

module \./br1.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11,
    z3  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11;
  output z3;
  assign z3 = ~x2 | ~x3;
endmodule


