module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 ;
  assign n16 = x6 & ~x11 ;
  assign n17 = ~x0 & ~x2 ;
  assign n18 = x13 & ~x14 ;
  assign n19 = ~x1 & ~x7 ;
  assign n20 = n18 & n19 ;
  assign n21 = n17 & n20 ;
  assign n22 = x3 & ~x5 ;
  assign n23 = x8 & x9 ;
  assign n24 = ~x4 & x10 ;
  assign n25 = n23 & n24 ;
  assign n26 = ~n22 & n25 ;
  assign n27 = n21 & n26 ;
  assign n28 = ~x13 & x14 ;
  assign n29 = n22 & n28 ;
  assign n30 = ~x4 & x9 ;
  assign n31 = ~x7 & ~n30 ;
  assign n32 = n29 & ~n31 ;
  assign n33 = x0 & x2 ;
  assign n34 = n33 ^ x4 ;
  assign n35 = n33 ^ x1 ;
  assign n36 = n35 ^ x1 ;
  assign n37 = x10 ^ x1 ;
  assign n38 = n36 & n37 ;
  assign n39 = n38 ^ x1 ;
  assign n40 = n34 & ~n39 ;
  assign n41 = n40 ^ x4 ;
  assign n42 = n32 & n41 ;
  assign n43 = x9 ^ x8 ;
  assign n44 = x9 & x10 ;
  assign n45 = n43 & n44 ;
  assign n46 = n45 ^ n43 ;
  assign n47 = x4 & ~n46 ;
  assign n48 = n47 ^ x1 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = x10 & n17 ;
  assign n51 = x4 & ~n50 ;
  assign n52 = x7 & n23 ;
  assign n53 = n52 ^ x8 ;
  assign n54 = ~n51 & n53 ;
  assign n55 = n54 ^ n47 ;
  assign n56 = n49 & n55 ;
  assign n57 = n56 ^ n47 ;
  assign n58 = n42 & n57 ;
  assign n59 = ~n27 & ~n58 ;
  assign n60 = n59 ^ x12 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = ~x5 & n18 ;
  assign n63 = ~x4 & n62 ;
  assign n64 = ~x8 & ~x9 ;
  assign n65 = ~x10 & n64 ;
  assign n66 = x3 ^ x2 ;
  assign n67 = ~x3 & n66 ;
  assign n68 = x1 & n67 ;
  assign n69 = n68 ^ n66 ;
  assign n70 = n65 & ~n69 ;
  assign n71 = x0 & x7 ;
  assign n72 = n70 & n71 ;
  assign n73 = n63 & n72 ;
  assign n74 = n73 ^ n59 ;
  assign n75 = n61 & ~n74 ;
  assign n76 = n75 ^ n59 ;
  assign n77 = n16 & ~n76 ;
  assign y0 = n77 ;
endmodule
