module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 ;
  assign n11 = x4 & x5 ;
  assign n12 = ~x2 & ~n11 ;
  assign n13 = ~x0 & n12 ;
  assign n14 = ~x4 & ~x5 ;
  assign n15 = n14 ^ x3 ;
  assign n16 = n14 ^ x1 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = n17 ^ n15 ;
  assign n22 = x7 & ~x8 ;
  assign n23 = x8 & x9 ;
  assign n24 = ~n22 & ~n23 ;
  assign n19 = x9 ^ x8 ;
  assign n20 = x7 & ~n19 ;
  assign n21 = n20 ^ x8 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = ~n14 & ~n25 ;
  assign n27 = n26 ^ n21 ;
  assign n28 = n18 & n27 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = n29 ^ n21 ;
  assign n31 = n30 ^ n14 ;
  assign n32 = ~n15 & ~n31 ;
  assign n33 = n32 ^ x3 ;
  assign n34 = ~x7 & x8 ;
  assign n35 = x1 & ~n22 ;
  assign n36 = ~n34 & n35 ;
  assign n37 = ~x1 & ~x3 ;
  assign n38 = n14 & n37 ;
  assign n39 = n38 ^ x6 ;
  assign n40 = n39 ^ x6 ;
  assign n41 = n19 ^ x8 ;
  assign n42 = n22 ^ x8 ;
  assign n43 = ~n41 & n42 ;
  assign n44 = n43 ^ x8 ;
  assign n45 = x6 & n44 ;
  assign n46 = n45 ^ x6 ;
  assign n47 = n40 & ~n46 ;
  assign n48 = n47 ^ x6 ;
  assign n49 = ~n36 & ~n48 ;
  assign n50 = ~n33 & n49 ;
  assign n51 = n13 & n50 ;
  assign y0 = n51 ;
endmodule
