// Benchmark "./pla/l8err.pla_dbb_orig_0NonExact" written by ABC on Fri Nov 20 10:23:10 2020

module \./pla/l8err.pla_dbb_orig_0NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = 1'b1;
endmodule


