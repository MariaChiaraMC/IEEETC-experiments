module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 ;
  assign n17 = x8 & x10 ;
  assign n18 = ~x8 & ~x10 ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = ~x2 & x6 ;
  assign n21 = ~x0 & x1 ;
  assign n22 = ~x5 & ~x7 ;
  assign n23 = n21 & n22 ;
  assign n24 = x0 & ~x1 ;
  assign n25 = x5 & x7 ;
  assign n26 = n24 & n25 ;
  assign n27 = ~n23 & ~n26 ;
  assign n28 = x3 & x11 ;
  assign n29 = x9 & n28 ;
  assign n30 = ~x4 & n29 ;
  assign n31 = ~x3 & ~x4 ;
  assign n32 = ~x12 & n31 ;
  assign n33 = ~x14 & x15 ;
  assign n34 = x9 & x11 ;
  assign n35 = ~x13 & n34 ;
  assign n36 = n33 & n35 ;
  assign n37 = n32 & n36 ;
  assign n38 = ~x12 & x13 ;
  assign n39 = ~x9 & ~x11 ;
  assign n40 = n38 & n39 ;
  assign n41 = x3 & x4 ;
  assign n42 = x14 & x15 ;
  assign n43 = x14 & ~n42 ;
  assign n44 = n41 & ~n43 ;
  assign n45 = n40 & n44 ;
  assign n46 = ~n37 & ~n45 ;
  assign n47 = ~n30 & n46 ;
  assign n48 = ~n27 & ~n47 ;
  assign n49 = x12 & x13 ;
  assign n50 = ~x0 & x3 ;
  assign n51 = n49 & n50 ;
  assign n52 = ~x9 & n25 ;
  assign n53 = x4 & ~x11 ;
  assign n54 = n52 & n53 ;
  assign n55 = n51 & n54 ;
  assign n56 = ~n48 & ~n55 ;
  assign n57 = x1 & n22 ;
  assign n58 = ~x0 & ~x12 ;
  assign n59 = n34 & n41 ;
  assign n60 = n58 & n59 ;
  assign n61 = x0 & x13 ;
  assign n62 = x12 & x14 ;
  assign n63 = ~x3 & x15 ;
  assign n64 = n62 & n63 ;
  assign n65 = n39 & n64 ;
  assign n66 = x3 & x9 ;
  assign n67 = x11 & ~x12 ;
  assign n68 = n66 & n67 ;
  assign n69 = ~n65 & ~n68 ;
  assign n70 = n61 & ~n69 ;
  assign n71 = x4 & x15 ;
  assign n72 = ~x14 & n58 ;
  assign n73 = x3 & ~x9 ;
  assign n74 = ~x11 & ~x13 ;
  assign n75 = n73 & n74 ;
  assign n76 = n72 & n75 ;
  assign n77 = ~x0 & ~x14 ;
  assign n78 = x0 & x14 ;
  assign n79 = ~n77 & ~n78 ;
  assign n80 = ~x3 & n79 ;
  assign n81 = x12 & n34 ;
  assign n82 = ~x13 & ~n50 ;
  assign n83 = n81 & n82 ;
  assign n84 = ~n80 & n83 ;
  assign n85 = x0 & x3 ;
  assign n86 = ~x12 & ~x14 ;
  assign n87 = ~n62 & ~n86 ;
  assign n88 = ~x11 & x13 ;
  assign n89 = ~x9 & n88 ;
  assign n90 = ~n87 & n89 ;
  assign n91 = n85 & n90 ;
  assign n92 = ~n84 & ~n91 ;
  assign n93 = ~n76 & n92 ;
  assign n94 = n71 & ~n93 ;
  assign n95 = ~n70 & ~n94 ;
  assign n96 = ~n60 & n95 ;
  assign n97 = n57 & ~n96 ;
  assign n98 = x4 & x7 ;
  assign n99 = ~x11 & ~x12 ;
  assign n100 = ~x3 & x5 ;
  assign n101 = x0 & ~x9 ;
  assign n102 = n100 & n101 ;
  assign n103 = ~n99 & n102 ;
  assign n104 = ~x0 & x5 ;
  assign n105 = n34 & n104 ;
  assign n106 = ~x3 & n105 ;
  assign n107 = x0 & ~x5 ;
  assign n108 = n73 & ~n107 ;
  assign n109 = ~x11 & n38 ;
  assign n110 = x5 & x11 ;
  assign n111 = ~x0 & ~n110 ;
  assign n112 = ~n109 & n111 ;
  assign n113 = n108 & ~n112 ;
  assign n114 = ~n106 & ~n113 ;
  assign n115 = ~n103 & n114 ;
  assign n116 = n98 & ~n115 ;
  assign n117 = ~x0 & ~x3 ;
  assign n118 = ~x5 & n34 ;
  assign n119 = x4 & x13 ;
  assign n120 = ~x12 & n119 ;
  assign n121 = x7 & n49 ;
  assign n122 = ~n120 & ~n121 ;
  assign n123 = n118 & ~n122 ;
  assign n124 = n117 & n123 ;
  assign n125 = ~n116 & ~n124 ;
  assign n126 = n125 ^ x1 ;
  assign n127 = n126 ^ n125 ;
  assign n128 = n127 ^ n97 ;
  assign n129 = x3 & x5 ;
  assign n130 = ~x7 & n129 ;
  assign n131 = n38 & n130 ;
  assign n132 = ~x0 & ~x5 ;
  assign n133 = x12 & ~x13 ;
  assign n134 = ~n38 & ~n133 ;
  assign n135 = ~x7 & n33 ;
  assign n136 = ~n38 & ~n135 ;
  assign n137 = ~n134 & ~n136 ;
  assign n138 = n137 ^ x7 ;
  assign n139 = n138 ^ n137 ;
  assign n140 = x13 & x15 ;
  assign n141 = n140 ^ n137 ;
  assign n142 = n141 ^ n137 ;
  assign n143 = ~n139 & n142 ;
  assign n144 = n143 ^ n137 ;
  assign n145 = ~x3 & n144 ;
  assign n146 = n145 ^ n137 ;
  assign n147 = n132 & n146 ;
  assign n148 = x0 & x7 ;
  assign n149 = x3 & ~x5 ;
  assign n150 = n38 & n149 ;
  assign n151 = ~n100 & ~n150 ;
  assign n152 = n148 & ~n151 ;
  assign n153 = ~x12 & ~x13 ;
  assign n154 = n25 & n117 ;
  assign n155 = ~n153 & n154 ;
  assign n156 = ~n152 & ~n155 ;
  assign n157 = ~n147 & n156 ;
  assign n158 = ~n131 & n157 ;
  assign n159 = n34 & ~n158 ;
  assign n160 = x15 & n49 ;
  assign n161 = x14 & n49 ;
  assign n162 = ~n160 & ~n161 ;
  assign n163 = n39 & n154 ;
  assign n164 = ~n162 & n163 ;
  assign n165 = x0 & x5 ;
  assign n166 = x7 & n165 ;
  assign n167 = ~x9 & ~x12 ;
  assign n168 = ~x11 & n140 ;
  assign n169 = n167 & n168 ;
  assign n170 = n166 & n169 ;
  assign n171 = ~x3 & n170 ;
  assign n172 = ~n164 & ~n171 ;
  assign n173 = ~n159 & n172 ;
  assign n174 = n173 ^ x4 ;
  assign n175 = x4 & ~n174 ;
  assign n176 = n175 ^ n125 ;
  assign n177 = n176 ^ x4 ;
  assign n178 = n128 & ~n177 ;
  assign n179 = n178 ^ n175 ;
  assign n180 = n179 ^ x4 ;
  assign n181 = ~n97 & n180 ;
  assign n182 = n181 ^ n97 ;
  assign n183 = n56 & ~n182 ;
  assign n184 = n20 & ~n183 ;
  assign n185 = x1 & ~x7 ;
  assign n186 = n39 & n140 ;
  assign n187 = n100 & n186 ;
  assign n188 = n185 & n187 ;
  assign n189 = ~x1 & x7 ;
  assign n190 = ~x5 & x15 ;
  assign n191 = x3 & n39 ;
  assign n192 = x13 & n191 ;
  assign n193 = n190 & n192 ;
  assign n194 = x5 & ~x13 ;
  assign n195 = ~x3 & n34 ;
  assign n196 = n194 & n195 ;
  assign n197 = ~n193 & ~n196 ;
  assign n198 = n189 & ~n197 ;
  assign n199 = x3 & n185 ;
  assign n200 = ~x5 & ~x13 ;
  assign n201 = n34 & n200 ;
  assign n202 = n199 & n201 ;
  assign n203 = ~n198 & ~n202 ;
  assign n204 = ~n188 & n203 ;
  assign n205 = ~x0 & x6 ;
  assign n206 = ~x4 & n205 ;
  assign n207 = ~x2 & x4 ;
  assign n208 = ~x6 & n207 ;
  assign n209 = ~n206 & ~n208 ;
  assign n210 = ~x0 & ~x2 ;
  assign n211 = n87 & ~n210 ;
  assign n212 = ~n209 & n211 ;
  assign n213 = ~n204 & n212 ;
  assign n214 = x9 & x13 ;
  assign n215 = x11 & x12 ;
  assign n216 = n214 & n215 ;
  assign n217 = ~x5 & x7 ;
  assign n218 = ~x2 & n41 ;
  assign n219 = n217 & n218 ;
  assign n220 = n24 & n219 ;
  assign n221 = x1 & ~x2 ;
  assign n222 = x4 & x5 ;
  assign n223 = n117 & n222 ;
  assign n224 = ~n31 & ~n41 ;
  assign n225 = n107 & n224 ;
  assign n226 = ~n223 & ~n225 ;
  assign n227 = n221 & ~n226 ;
  assign n228 = x2 & x4 ;
  assign n229 = ~x0 & n228 ;
  assign n230 = ~x3 & ~x5 ;
  assign n231 = ~n129 & ~n230 ;
  assign n232 = ~x1 & n231 ;
  assign n233 = n229 & n232 ;
  assign n234 = x2 & n21 ;
  assign n235 = x3 & ~x4 ;
  assign n236 = ~x5 & n235 ;
  assign n237 = n234 & n236 ;
  assign n238 = ~n233 & ~n237 ;
  assign n239 = ~n227 & n238 ;
  assign n240 = ~x7 & ~n239 ;
  assign n241 = ~n220 & ~n240 ;
  assign n242 = n216 & ~n241 ;
  assign n243 = ~n213 & ~n242 ;
  assign n244 = x0 & ~x12 ;
  assign n245 = ~x0 & x12 ;
  assign n246 = ~n244 & ~n245 ;
  assign n247 = x2 & ~x4 ;
  assign n248 = ~n207 & ~n247 ;
  assign n249 = ~x4 & ~x6 ;
  assign n250 = ~x4 & x14 ;
  assign n251 = ~n249 & ~n250 ;
  assign n252 = x4 & x6 ;
  assign n253 = x4 & ~x14 ;
  assign n254 = ~n252 & ~n253 ;
  assign n255 = n251 & n254 ;
  assign n256 = ~n248 & n255 ;
  assign n257 = ~x7 & x9 ;
  assign n258 = ~x1 & x5 ;
  assign n259 = x11 & ~x13 ;
  assign n260 = n258 & n259 ;
  assign n261 = n257 & n260 ;
  assign n262 = n256 & n261 ;
  assign n263 = x1 & ~x5 ;
  assign n264 = x7 & ~x9 ;
  assign n265 = n88 & n264 ;
  assign n266 = ~x2 & ~x4 ;
  assign n267 = x6 & x14 ;
  assign n268 = n266 & n267 ;
  assign n269 = ~x6 & ~x14 ;
  assign n270 = n228 & n269 ;
  assign n271 = ~n268 & ~n270 ;
  assign n272 = n265 & ~n271 ;
  assign n273 = n263 & n272 ;
  assign n274 = ~n262 & ~n273 ;
  assign n275 = ~n246 & ~n274 ;
  assign n276 = ~n185 & ~n189 ;
  assign n277 = ~x6 & x12 ;
  assign n278 = ~x0 & x4 ;
  assign n279 = n277 & n278 ;
  assign n280 = ~x2 & x5 ;
  assign n281 = x13 & x14 ;
  assign n282 = n39 & n281 ;
  assign n283 = n280 & n282 ;
  assign n284 = ~x13 & ~x14 ;
  assign n285 = x11 & n284 ;
  assign n286 = x2 & x9 ;
  assign n287 = ~x5 & n286 ;
  assign n288 = n285 & n287 ;
  assign n289 = ~n283 & ~n288 ;
  assign n290 = n279 & ~n289 ;
  assign n291 = ~x4 & x6 ;
  assign n292 = ~x2 & x14 ;
  assign n293 = n201 & n292 ;
  assign n294 = x13 & ~x14 ;
  assign n295 = x2 & x5 ;
  assign n296 = n39 & n295 ;
  assign n297 = n294 & n296 ;
  assign n298 = ~n293 & ~n297 ;
  assign n299 = n244 & ~n298 ;
  assign n300 = n291 & n299 ;
  assign n301 = ~n290 & ~n300 ;
  assign n302 = ~n276 & ~n301 ;
  assign n303 = ~n275 & ~n302 ;
  assign n304 = ~x3 & ~x15 ;
  assign n305 = ~n303 & ~n304 ;
  assign n306 = x6 & n228 ;
  assign n307 = ~x0 & ~x9 ;
  assign n308 = x1 & x3 ;
  assign n309 = n22 & n308 ;
  assign n310 = ~x14 & n140 ;
  assign n311 = n99 & n310 ;
  assign n312 = n309 & n311 ;
  assign n313 = ~x1 & x3 ;
  assign n314 = ~x11 & x12 ;
  assign n315 = n313 & ~n314 ;
  assign n316 = ~x3 & n25 ;
  assign n317 = n99 ^ n25 ;
  assign n318 = ~x1 & ~x13 ;
  assign n319 = n42 & n318 ;
  assign n320 = ~n140 & ~n294 ;
  assign n321 = ~x1 & ~n140 ;
  assign n322 = ~n320 & ~n321 ;
  assign n323 = ~n319 & ~n322 ;
  assign n324 = n323 ^ n316 ;
  assign n325 = n317 & n324 ;
  assign n326 = n325 ^ n323 ;
  assign n327 = n316 & n326 ;
  assign n328 = n327 ^ n25 ;
  assign n329 = ~n315 & n328 ;
  assign n330 = ~n312 & ~n329 ;
  assign n331 = n307 & ~n330 ;
  assign n332 = ~x0 & n118 ;
  assign n333 = ~x1 & ~x7 ;
  assign n334 = n42 & n133 ;
  assign n335 = n333 & n334 ;
  assign n336 = x3 & n335 ;
  assign n337 = x1 & ~x12 ;
  assign n338 = ~x3 & x7 ;
  assign n339 = n337 & n338 ;
  assign n340 = n339 ^ x13 ;
  assign n341 = n340 ^ n339 ;
  assign n342 = n341 ^ n336 ;
  assign n343 = x12 & x15 ;
  assign n344 = n343 ^ n199 ;
  assign n345 = n199 & n344 ;
  assign n346 = n345 ^ n339 ;
  assign n347 = n346 ^ n199 ;
  assign n348 = n342 & n347 ;
  assign n349 = n348 ^ n345 ;
  assign n350 = n349 ^ n199 ;
  assign n351 = ~n336 & n350 ;
  assign n352 = n351 ^ n336 ;
  assign n353 = n332 & n352 ;
  assign n354 = ~x1 & ~x3 ;
  assign n355 = ~n308 & ~n354 ;
  assign n356 = x13 & n215 ;
  assign n357 = x0 & x9 ;
  assign n358 = n22 & n357 ;
  assign n359 = n356 & n358 ;
  assign n360 = n355 & n359 ;
  assign n361 = n39 & n49 ;
  assign n362 = n309 & n361 ;
  assign n363 = n39 & n308 ;
  assign n364 = x1 & x9 ;
  assign n365 = ~x3 & n364 ;
  assign n366 = n259 & n365 ;
  assign n367 = ~n363 & ~n366 ;
  assign n368 = n22 & ~n367 ;
  assign n369 = ~x1 & ~x11 ;
  assign n370 = n52 & n369 ;
  assign n371 = ~x3 & n370 ;
  assign n372 = x3 & n318 ;
  assign n373 = n22 & n34 ;
  assign n374 = n372 & n373 ;
  assign n375 = ~n371 & ~n374 ;
  assign n376 = ~n368 & n375 ;
  assign n377 = n244 & ~n376 ;
  assign n378 = ~n362 & ~n377 ;
  assign n379 = ~n360 & n378 ;
  assign n380 = n42 & ~n379 ;
  assign n381 = ~n353 & ~n380 ;
  assign n382 = ~n331 & n381 ;
  assign n383 = n306 & ~n382 ;
  assign n384 = ~x3 & x9 ;
  assign n385 = n259 & n384 ;
  assign n386 = n385 ^ n192 ;
  assign n387 = n386 ^ n192 ;
  assign n388 = n192 ^ x15 ;
  assign n389 = n388 ^ n192 ;
  assign n390 = n387 & n389 ;
  assign n391 = n390 ^ n192 ;
  assign n392 = ~x5 & n391 ;
  assign n393 = n392 ^ n192 ;
  assign n403 = x6 & x12 ;
  assign n404 = ~x4 & n403 ;
  assign n394 = x4 & ~x6 ;
  assign n395 = ~x12 & n394 ;
  assign n396 = ~x1 & x2 ;
  assign n397 = x7 & ~x14 ;
  assign n398 = n396 & n397 ;
  assign n399 = ~x7 & x14 ;
  assign n400 = n221 & n399 ;
  assign n401 = ~n398 & ~n400 ;
  assign n402 = n395 & ~n401 ;
  assign n405 = n404 ^ n402 ;
  assign n406 = n405 ^ n402 ;
  assign n407 = x2 ^ x1 ;
  assign n409 = ~x7 & ~x14 ;
  assign n408 = x7 & x14 ;
  assign n410 = n409 ^ n408 ;
  assign n411 = n409 ^ x2 ;
  assign n412 = n411 ^ n409 ;
  assign n413 = n410 & ~n412 ;
  assign n414 = n413 ^ n409 ;
  assign n415 = ~n407 & n414 ;
  assign n416 = n415 ^ n402 ;
  assign n417 = n416 ^ n402 ;
  assign n418 = n406 & n417 ;
  assign n419 = n418 ^ n402 ;
  assign n420 = ~x0 & n419 ;
  assign n421 = n420 ^ n402 ;
  assign n422 = n393 & n421 ;
  assign n423 = ~n383 & ~n422 ;
  assign n424 = ~n305 & n423 ;
  assign n425 = x6 & x13 ;
  assign n426 = ~x1 & x12 ;
  assign n427 = n338 & n426 ;
  assign n428 = n332 & n427 ;
  assign n429 = ~x0 & ~x7 ;
  assign n430 = n313 & n314 ;
  assign n431 = ~x5 & ~x9 ;
  assign n432 = n42 & n431 ;
  assign n433 = n430 & n432 ;
  assign n434 = x5 & x12 ;
  assign n435 = ~n149 & ~n434 ;
  assign n436 = x3 & x12 ;
  assign n437 = x11 & n364 ;
  assign n438 = ~n436 & n437 ;
  assign n439 = ~n435 & n438 ;
  assign n440 = ~n433 & ~n439 ;
  assign n441 = n429 & ~n440 ;
  assign n442 = n26 & n65 ;
  assign n443 = ~n441 & ~n442 ;
  assign n444 = ~n428 & n443 ;
  assign n445 = n425 & ~n444 ;
  assign n446 = x2 & n445 ;
  assign n447 = n424 & ~n446 ;
  assign n448 = n243 & n447 ;
  assign n449 = ~n184 & n448 ;
  assign n450 = x0 & x1 ;
  assign n451 = ~x3 & ~x7 ;
  assign n452 = n216 & n451 ;
  assign n453 = ~x3 & n217 ;
  assign n454 = n34 & n38 ;
  assign n455 = n453 & n454 ;
  assign n456 = ~n452 & ~n455 ;
  assign n457 = ~n73 & ~n384 ;
  assign n458 = n457 ^ x11 ;
  assign n459 = n458 ^ n457 ;
  assign n460 = ~x9 & n49 ;
  assign n461 = n460 ^ n457 ;
  assign n462 = ~n459 & ~n461 ;
  assign n463 = n462 ^ n457 ;
  assign n464 = n25 & ~n463 ;
  assign n465 = n456 & ~n464 ;
  assign n466 = x3 & ~x7 ;
  assign n467 = n186 & n466 ;
  assign n468 = x7 & n39 ;
  assign n469 = ~x3 & x13 ;
  assign n470 = ~x14 & ~x15 ;
  assign n471 = n469 & ~n470 ;
  assign n472 = n468 & n471 ;
  assign n473 = x7 & x11 ;
  assign n474 = n384 & n473 ;
  assign n475 = ~x13 & x15 ;
  assign n476 = ~n284 & ~n475 ;
  assign n477 = n28 & n257 ;
  assign n478 = ~n476 & n477 ;
  assign n479 = ~n474 & ~n478 ;
  assign n480 = ~n472 & n479 ;
  assign n483 = n480 ^ x3 ;
  assign n484 = n483 ^ n480 ;
  assign n481 = n480 ^ n33 ;
  assign n482 = n481 ^ n480 ;
  assign n485 = n484 ^ n482 ;
  assign n486 = n257 & n259 ;
  assign n487 = ~n265 & ~n486 ;
  assign n488 = n487 ^ n480 ;
  assign n489 = n488 ^ n480 ;
  assign n490 = n489 ^ n484 ;
  assign n491 = n484 & ~n490 ;
  assign n492 = n491 ^ n484 ;
  assign n493 = n485 & n492 ;
  assign n494 = n493 ^ n491 ;
  assign n495 = n494 ^ n480 ;
  assign n496 = n495 ^ n484 ;
  assign n497 = ~x12 & ~n496 ;
  assign n498 = n497 ^ n480 ;
  assign n499 = ~n467 & n498 ;
  assign n500 = n499 ^ x5 ;
  assign n501 = n500 ^ n499 ;
  assign n502 = n501 ^ n465 ;
  assign n503 = x12 & ~x14 ;
  assign n504 = ~n343 & ~n503 ;
  assign n505 = ~n192 & ~n385 ;
  assign n506 = ~n504 & ~n505 ;
  assign n507 = ~x3 & ~x9 ;
  assign n508 = n168 & n507 ;
  assign n509 = ~n506 & ~n508 ;
  assign n510 = n509 ^ x7 ;
  assign n511 = ~x7 & n510 ;
  assign n512 = n511 ^ n499 ;
  assign n513 = n512 ^ x7 ;
  assign n514 = n502 & n513 ;
  assign n515 = n514 ^ n511 ;
  assign n516 = n515 ^ x7 ;
  assign n517 = n465 & ~n516 ;
  assign n518 = n517 ^ n465 ;
  assign n519 = n450 & ~n518 ;
  assign n520 = n217 & n313 ;
  assign n521 = n216 & n520 ;
  assign n522 = x3 & x7 ;
  assign n523 = n165 & n522 ;
  assign n524 = n40 & n523 ;
  assign n525 = x1 & n231 ;
  assign n526 = x5 & n313 ;
  assign n527 = ~n525 & ~n526 ;
  assign n528 = ~x13 & x14 ;
  assign n529 = ~n38 & ~n528 ;
  assign n530 = n39 & n529 ;
  assign n531 = ~n527 & n530 ;
  assign n532 = ~x1 & ~x12 ;
  assign n533 = ~x14 & n532 ;
  assign n534 = n35 & n533 ;
  assign n535 = n231 & n534 ;
  assign n536 = ~n531 & ~n535 ;
  assign n537 = x15 & ~n536 ;
  assign n538 = ~x1 & x11 ;
  assign n539 = n66 & n538 ;
  assign n540 = n73 & n99 ;
  assign n541 = ~n195 & ~n540 ;
  assign n542 = x1 & ~n541 ;
  assign n543 = ~n539 & ~n542 ;
  assign n544 = x5 & ~n543 ;
  assign n545 = ~n537 & ~n544 ;
  assign n546 = n429 & ~n545 ;
  assign n547 = ~n524 & ~n546 ;
  assign n548 = ~n521 & n547 ;
  assign n549 = ~x0 & x7 ;
  assign n550 = x1 & ~x3 ;
  assign n551 = x5 & ~x9 ;
  assign n552 = n88 & n551 ;
  assign n553 = ~n201 & ~n552 ;
  assign n554 = n550 & ~n553 ;
  assign n555 = n62 & n554 ;
  assign n556 = x3 & ~x12 ;
  assign n557 = n201 & ~n556 ;
  assign n558 = ~n313 & ~n550 ;
  assign n559 = ~n62 & ~n558 ;
  assign n560 = n557 & n559 ;
  assign n561 = ~x14 & n49 ;
  assign n562 = n39 & n526 ;
  assign n563 = n561 & n562 ;
  assign n564 = ~n560 & ~n563 ;
  assign n565 = ~n100 & ~n149 ;
  assign n566 = n34 & n153 ;
  assign n567 = n39 & n161 ;
  assign n568 = ~n566 & ~n567 ;
  assign n569 = ~x1 & ~n568 ;
  assign n570 = ~x9 & x12 ;
  assign n571 = x1 & ~x11 ;
  assign n572 = n570 & n571 ;
  assign n573 = n294 & n572 ;
  assign n574 = ~n569 & ~n573 ;
  assign n575 = ~n565 & ~n574 ;
  assign n576 = n564 & ~n575 ;
  assign n577 = x15 & ~n576 ;
  assign n578 = n308 & n551 ;
  assign n579 = n62 & n539 ;
  assign n580 = n200 & n579 ;
  assign n581 = ~n578 & ~n580 ;
  assign n582 = ~n577 & n581 ;
  assign n583 = ~n555 & n582 ;
  assign n584 = n549 & ~n583 ;
  assign n585 = ~x13 & n33 ;
  assign n586 = ~x7 & x12 ;
  assign n587 = x7 & ~x12 ;
  assign n588 = ~n586 & ~n587 ;
  assign n589 = n585 & ~n588 ;
  assign n590 = n149 & n589 ;
  assign n591 = x7 & x12 ;
  assign n592 = x15 & n22 ;
  assign n593 = ~n591 & ~n592 ;
  assign n594 = n469 & ~n593 ;
  assign n595 = ~n150 & ~n594 ;
  assign n596 = ~n590 & n595 ;
  assign n597 = n34 & ~n596 ;
  assign n598 = x12 & ~x15 ;
  assign n599 = n192 & n409 ;
  assign n600 = n474 & n528 ;
  assign n601 = ~n599 & ~n600 ;
  assign n602 = ~n598 & ~n601 ;
  assign n603 = x9 & x12 ;
  assign n604 = n284 & n603 ;
  assign n605 = x11 & n604 ;
  assign n606 = ~n186 & ~n605 ;
  assign n607 = n338 & ~n606 ;
  assign n608 = ~x7 & ~x12 ;
  assign n609 = ~n281 & ~n284 ;
  assign n610 = x15 & n39 ;
  assign n611 = ~n609 & n610 ;
  assign n612 = ~n34 & ~n611 ;
  assign n613 = n608 & ~n612 ;
  assign n614 = n613 ^ x3 ;
  assign n615 = n614 ^ n613 ;
  assign n616 = n615 ^ n607 ;
  assign n617 = n137 ^ n34 ;
  assign n618 = n137 & n617 ;
  assign n619 = n618 ^ n613 ;
  assign n620 = n619 ^ n137 ;
  assign n621 = n616 & n620 ;
  assign n622 = n621 ^ n618 ;
  assign n623 = n622 ^ n137 ;
  assign n624 = ~n607 & n623 ;
  assign n625 = n624 ^ n607 ;
  assign n626 = ~n602 & ~n625 ;
  assign n627 = x5 & ~n626 ;
  assign n628 = n186 & n217 ;
  assign n629 = x3 & n628 ;
  assign n630 = ~n627 & ~n629 ;
  assign n631 = ~n597 & n630 ;
  assign n632 = n24 & ~n631 ;
  assign n633 = ~n584 & ~n632 ;
  assign n634 = n548 & n633 ;
  assign n635 = ~n519 & n634 ;
  assign n636 = n266 & ~n635 ;
  assign n637 = n132 & n265 ;
  assign n638 = ~x0 & ~x13 ;
  assign n639 = ~x14 & n638 ;
  assign n640 = x5 & ~x7 ;
  assign n641 = n39 & n640 ;
  assign n642 = ~x5 & x9 ;
  assign n643 = n473 & n642 ;
  assign n644 = ~n641 & ~n643 ;
  assign n645 = n639 & ~n644 ;
  assign n646 = n528 & n640 ;
  assign n647 = x11 & n357 ;
  assign n648 = n646 & n647 ;
  assign n649 = x5 & ~x14 ;
  assign n650 = n89 & n148 ;
  assign n651 = ~n649 & n650 ;
  assign n652 = ~n648 & ~n651 ;
  assign n653 = ~n645 & n652 ;
  assign n654 = ~x12 & ~n653 ;
  assign n655 = x0 & x12 ;
  assign n656 = ~x7 & n655 ;
  assign n657 = ~n35 & ~n282 ;
  assign n658 = n657 ^ n528 ;
  assign n659 = n658 ^ n657 ;
  assign n660 = n657 ^ n34 ;
  assign n661 = n660 ^ n657 ;
  assign n662 = n659 & n661 ;
  assign n663 = n662 ^ n657 ;
  assign n664 = ~x5 & ~n663 ;
  assign n665 = n664 ^ n657 ;
  assign n666 = n656 & ~n665 ;
  assign n667 = ~n654 & ~n666 ;
  assign n668 = ~n637 & n667 ;
  assign n669 = n550 & ~n668 ;
  assign n670 = ~x12 & n265 ;
  assign n671 = ~n486 & ~n670 ;
  assign n672 = n165 & ~n671 ;
  assign n673 = ~n86 & n672 ;
  assign n674 = x9 & x14 ;
  assign n675 = ~x13 & n674 ;
  assign n676 = n215 & n675 ;
  assign n677 = ~n89 & ~n676 ;
  assign n678 = x5 & ~n677 ;
  assign n679 = ~x12 & n528 ;
  assign n680 = n118 & n679 ;
  assign n681 = ~n678 & ~n680 ;
  assign n682 = n429 & ~n681 ;
  assign n683 = n107 & n670 ;
  assign n684 = x0 & n22 ;
  assign n685 = n676 & n684 ;
  assign n686 = ~n683 & ~n685 ;
  assign n687 = ~n682 & n686 ;
  assign n688 = ~n673 & n687 ;
  assign n689 = n313 & ~n688 ;
  assign n690 = n25 & n354 ;
  assign n691 = ~n309 & ~n690 ;
  assign n692 = ~x0 & x9 ;
  assign n693 = n259 & n692 ;
  assign n694 = ~n691 & n693 ;
  assign n695 = n61 & n640 ;
  assign n696 = n39 & n695 ;
  assign n697 = n313 & n696 ;
  assign n698 = ~n694 & ~n697 ;
  assign n699 = ~n87 & ~n698 ;
  assign n700 = n549 & n552 ;
  assign n701 = ~x5 & ~x14 ;
  assign n702 = ~n104 & ~n701 ;
  assign n703 = n35 & n246 ;
  assign n704 = n702 & n703 ;
  assign n705 = n704 ^ x13 ;
  assign n706 = n705 ^ n704 ;
  assign n707 = n704 ^ n332 ;
  assign n708 = n707 ^ n704 ;
  assign n709 = n706 & n708 ;
  assign n710 = n709 ^ n704 ;
  assign n711 = ~x7 & n710 ;
  assign n712 = n711 ^ n704 ;
  assign n713 = ~n700 & ~n712 ;
  assign n714 = n354 & ~n713 ;
  assign n715 = ~n699 & ~n714 ;
  assign n716 = n679 & n684 ;
  assign n717 = ~x12 & n294 ;
  assign n718 = ~x0 & n217 ;
  assign n719 = n717 & n718 ;
  assign n720 = ~n132 & n246 ;
  assign n721 = ~x7 & x13 ;
  assign n722 = ~n649 & n721 ;
  assign n723 = ~n720 & n722 ;
  assign n724 = ~n719 & ~n723 ;
  assign n725 = ~n716 & n724 ;
  assign n726 = n363 & ~n725 ;
  assign n727 = n715 & ~n726 ;
  assign n728 = ~n689 & n727 ;
  assign n729 = ~n669 & n728 ;
  assign n730 = x15 & ~n729 ;
  assign n731 = x5 & ~x12 ;
  assign n732 = n469 & n731 ;
  assign n733 = ~n149 & ~n732 ;
  assign n734 = n148 & ~n733 ;
  assign n735 = ~n131 & ~n734 ;
  assign n736 = ~x1 & ~n735 ;
  assign n737 = n217 & n528 ;
  assign n738 = ~n640 & ~n737 ;
  assign n739 = n117 & n337 ;
  assign n740 = ~n738 & n739 ;
  assign n741 = ~n736 & ~n740 ;
  assign n742 = ~x1 & n436 ;
  assign n743 = ~n217 & ~n721 ;
  assign n744 = n742 & ~n743 ;
  assign n745 = ~n258 & ~n263 ;
  assign n746 = ~x3 & ~n745 ;
  assign n747 = ~n520 & ~n746 ;
  assign n748 = n38 & ~n747 ;
  assign n749 = ~n744 & ~n748 ;
  assign n750 = n749 ^ x0 ;
  assign n751 = n750 ^ n749 ;
  assign n752 = ~n217 & ~n640 ;
  assign n753 = ~x14 & n153 ;
  assign n754 = ~n217 & ~n753 ;
  assign n755 = ~n752 & ~n754 ;
  assign n756 = n550 & n755 ;
  assign n757 = ~n309 & ~n756 ;
  assign n758 = n757 ^ n749 ;
  assign n759 = n751 & n758 ;
  assign n760 = n759 ^ n749 ;
  assign n761 = n741 & n760 ;
  assign n762 = n34 & ~n761 ;
  assign n763 = x12 & n149 ;
  assign n764 = ~x14 & n732 ;
  assign n765 = ~n763 & ~n764 ;
  assign n766 = n450 & ~n765 ;
  assign n767 = n51 & ~n263 ;
  assign n768 = ~x0 & x13 ;
  assign n769 = ~n230 & n337 ;
  assign n770 = n768 & n769 ;
  assign n771 = ~n767 & ~n770 ;
  assign n772 = ~n701 & ~n771 ;
  assign n773 = ~n766 & ~n772 ;
  assign n774 = n468 & ~n773 ;
  assign n775 = x1 & x11 ;
  assign n776 = n50 & n775 ;
  assign n777 = n52 & n776 ;
  assign n778 = n25 & n101 ;
  assign n779 = n308 & n778 ;
  assign n780 = n294 & n608 ;
  assign n781 = n21 & n780 ;
  assign n782 = n39 & n100 ;
  assign n783 = n781 & n782 ;
  assign n784 = ~n779 & ~n783 ;
  assign n785 = ~n777 & n784 ;
  assign n786 = ~n774 & n785 ;
  assign n787 = ~n762 & n786 ;
  assign n788 = ~n730 & n787 ;
  assign n789 = n247 & ~n788 ;
  assign n790 = x13 & n34 ;
  assign n791 = n100 & n790 ;
  assign n792 = x1 & x4 ;
  assign n793 = ~x0 & n792 ;
  assign n794 = x12 & n549 ;
  assign n795 = ~n793 & ~n794 ;
  assign n796 = n795 ^ n608 ;
  assign n797 = n796 ^ n791 ;
  assign n799 = ~x1 & ~x4 ;
  assign n798 = ~x4 & n450 ;
  assign n800 = n799 ^ n798 ;
  assign n801 = n608 & ~n800 ;
  assign n802 = n801 ^ n799 ;
  assign n803 = ~n797 & n802 ;
  assign n804 = n803 ^ n801 ;
  assign n805 = n804 ^ n799 ;
  assign n806 = n805 ^ n608 ;
  assign n807 = n791 & n806 ;
  assign n808 = ~n789 & ~n807 ;
  assign n809 = ~n636 & n808 ;
  assign n810 = n809 ^ x6 ;
  assign n811 = n810 ^ n809 ;
  assign n812 = n357 & n538 ;
  assign n813 = n25 & n812 ;
  assign n814 = x0 & ~n109 ;
  assign n815 = ~n775 & n814 ;
  assign n816 = ~x0 & ~x1 ;
  assign n817 = ~x1 & x13 ;
  assign n818 = ~x11 & n817 ;
  assign n819 = n62 & n818 ;
  assign n820 = n816 & ~n819 ;
  assign n821 = ~n815 & ~n820 ;
  assign n822 = n52 & n821 ;
  assign n823 = ~n813 & ~n822 ;
  assign n824 = ~x7 & n434 ;
  assign n825 = n34 & n817 ;
  assign n826 = n824 & n825 ;
  assign n827 = n823 & ~n826 ;
  assign n828 = x3 & ~n827 ;
  assign n829 = x3 & ~x13 ;
  assign n830 = ~n469 & ~n829 ;
  assign n831 = n812 & ~n830 ;
  assign n832 = x3 & ~x14 ;
  assign n833 = ~n436 & ~n832 ;
  assign n834 = n831 & n833 ;
  assign n835 = n191 & n561 ;
  assign n836 = n195 & n679 ;
  assign n837 = ~n835 & ~n836 ;
  assign n838 = n450 & ~n837 ;
  assign n839 = ~n90 & ~n566 ;
  assign n840 = n308 & ~n839 ;
  assign n841 = ~x0 & n840 ;
  assign n842 = ~n838 & ~n841 ;
  assign n843 = ~n834 & n842 ;
  assign n844 = n22 & ~n843 ;
  assign n845 = n609 ^ n529 ;
  assign n846 = n845 ^ n529 ;
  assign n847 = n529 ^ x12 ;
  assign n848 = n847 ^ n529 ;
  assign n849 = ~n846 & ~n848 ;
  assign n850 = n849 ^ n529 ;
  assign n851 = x0 & n850 ;
  assign n852 = n851 ^ n529 ;
  assign n853 = n371 & n852 ;
  assign n854 = n51 & n370 ;
  assign n855 = ~x14 & n854 ;
  assign n856 = ~n853 & ~n855 ;
  assign n857 = ~n844 & n856 ;
  assign n858 = x15 & ~n857 ;
  assign n859 = n25 & n39 ;
  assign n860 = n739 & n859 ;
  assign n861 = x0 & ~x3 ;
  assign n862 = n258 & n264 ;
  assign n863 = n99 & n294 ;
  assign n864 = n862 & n863 ;
  assign n865 = ~x5 & n49 ;
  assign n866 = ~n25 & ~n865 ;
  assign n867 = x7 & n731 ;
  assign n868 = ~x1 & ~n867 ;
  assign n869 = n34 & ~n868 ;
  assign n870 = ~n866 & n869 ;
  assign n871 = ~n864 & ~n870 ;
  assign n872 = n861 & ~n871 ;
  assign n873 = ~x4 & ~n872 ;
  assign n874 = ~n860 & n873 ;
  assign n875 = ~x1 & n642 ;
  assign n876 = n356 & n875 ;
  assign n877 = n34 & ~n153 ;
  assign n878 = ~n567 & ~n877 ;
  assign n879 = n57 & ~n878 ;
  assign n880 = x1 & x12 ;
  assign n881 = n265 & n880 ;
  assign n882 = ~n879 & ~n881 ;
  assign n883 = ~n876 & n882 ;
  assign n884 = n85 & ~n883 ;
  assign n885 = n874 & ~n884 ;
  assign n886 = ~n858 & n885 ;
  assign n887 = ~n828 & n886 ;
  assign n888 = n454 & n520 ;
  assign n889 = n888 ^ x4 ;
  assign n890 = ~x12 & x14 ;
  assign n891 = ~n38 & ~n890 ;
  assign n892 = ~x7 & n34 ;
  assign n893 = ~n891 & n892 ;
  assign n894 = x7 & ~n62 ;
  assign n895 = n89 & ~n894 ;
  assign n896 = ~n87 & n486 ;
  assign n897 = ~n895 & ~n896 ;
  assign n898 = x15 & ~n897 ;
  assign n899 = ~n893 & ~n898 ;
  assign n900 = n308 & ~n899 ;
  assign n901 = n320 & ~n585 ;
  assign n902 = n39 & ~n901 ;
  assign n903 = ~n34 & ~n902 ;
  assign n904 = n339 & ~n903 ;
  assign n905 = ~x1 & x15 ;
  assign n906 = n522 & ~n677 ;
  assign n907 = x3 & n890 ;
  assign n908 = n486 & n907 ;
  assign n909 = x11 & x13 ;
  assign n910 = ~x7 & n909 ;
  assign n911 = n384 & n910 ;
  assign n912 = ~n908 & ~n911 ;
  assign n913 = ~n906 & n912 ;
  assign n914 = n905 & ~n913 ;
  assign n915 = ~n904 & ~n914 ;
  assign n916 = ~n900 & n915 ;
  assign n917 = ~x5 & ~n916 ;
  assign n918 = ~x1 & n25 ;
  assign n919 = ~x15 & ~n87 ;
  assign n920 = n385 & ~n919 ;
  assign n921 = n918 & n920 ;
  assign n922 = n384 & n909 ;
  assign n923 = ~x12 & n922 ;
  assign n924 = ~n276 & n923 ;
  assign n925 = ~n921 & ~n924 ;
  assign n926 = ~x1 & ~x14 ;
  assign n927 = x1 & x14 ;
  assign n928 = ~n926 & ~n927 ;
  assign n929 = x15 & n928 ;
  assign n930 = n929 ^ n927 ;
  assign n931 = ~x12 & n930 ;
  assign n932 = ~n505 & n931 ;
  assign n933 = ~x11 & n49 ;
  assign n934 = ~x1 & n73 ;
  assign n935 = ~n470 & n934 ;
  assign n936 = n933 & n935 ;
  assign n937 = n186 & n550 ;
  assign n938 = n313 & n877 ;
  assign n939 = ~n937 & ~n938 ;
  assign n940 = ~n936 & n939 ;
  assign n941 = ~n932 & n940 ;
  assign n942 = n640 & ~n941 ;
  assign n943 = x1 & ~x9 ;
  assign n944 = ~n28 & ~n109 ;
  assign n945 = n943 & ~n944 ;
  assign n946 = x12 ^ x3 ;
  assign n947 = n946 ^ x12 ;
  assign n948 = n947 ^ n89 ;
  assign n949 = n905 ^ x12 ;
  assign n950 = ~n948 & n949 ;
  assign n951 = n950 ^ n905 ;
  assign n952 = n89 & n951 ;
  assign n953 = ~n945 & ~n952 ;
  assign n954 = n25 & ~n953 ;
  assign n955 = ~n942 & ~n954 ;
  assign n956 = n925 & n955 ;
  assign n957 = ~n917 & n956 ;
  assign n958 = n957 ^ x0 ;
  assign n959 = n958 ^ n957 ;
  assign n960 = n343 & n675 ;
  assign n961 = n231 & n538 ;
  assign n962 = n960 & n961 ;
  assign n963 = ~x5 & n42 ;
  assign n964 = n385 & n963 ;
  assign n965 = n880 & n964 ;
  assign n966 = n129 & n572 ;
  assign n967 = ~n965 & ~n966 ;
  assign n968 = ~n34 & ~n169 ;
  assign n969 = ~n527 & ~n968 ;
  assign n970 = ~x7 & ~n969 ;
  assign n971 = n967 & n970 ;
  assign n972 = ~n962 & n971 ;
  assign n973 = x7 & ~n578 ;
  assign n974 = ~x1 & n149 ;
  assign n975 = n35 & n974 ;
  assign n976 = ~n554 & ~n975 ;
  assign n977 = ~n43 & ~n976 ;
  assign n978 = x5 ^ x3 ;
  assign n979 = n978 ^ x14 ;
  assign n980 = n979 ^ x1 ;
  assign n981 = n980 ^ n186 ;
  assign n982 = x5 ^ x1 ;
  assign n983 = n982 ^ x1 ;
  assign n984 = x14 ^ x1 ;
  assign n985 = n984 ^ x1 ;
  assign n986 = ~n983 & n985 ;
  assign n987 = n986 ^ x1 ;
  assign n988 = n987 ^ n980 ;
  assign n989 = n981 & ~n988 ;
  assign n990 = n989 ^ n986 ;
  assign n991 = n990 ^ x1 ;
  assign n992 = n991 ^ n186 ;
  assign n993 = n980 & ~n992 ;
  assign n994 = n993 ^ n980 ;
  assign n995 = ~n977 & ~n994 ;
  assign n996 = n995 ^ x12 ;
  assign n997 = n996 ^ n995 ;
  assign n998 = n89 & n525 ;
  assign n999 = ~x5 & n550 ;
  assign n1000 = ~n232 & ~n999 ;
  assign n1001 = x15 & ~n657 ;
  assign n1002 = ~n1000 & n1001 ;
  assign n1003 = ~n998 & ~n1002 ;
  assign n1004 = n1003 ^ n995 ;
  assign n1005 = n997 & n1004 ;
  assign n1006 = n1005 ^ n995 ;
  assign n1007 = n973 & n1006 ;
  assign n1008 = ~n972 & ~n1007 ;
  assign n1009 = n1008 ^ n957 ;
  assign n1010 = n959 & ~n1009 ;
  assign n1011 = n1010 ^ n957 ;
  assign n1012 = n1011 ^ n888 ;
  assign n1013 = ~n889 & ~n1012 ;
  assign n1014 = n1013 ^ n1010 ;
  assign n1015 = n1014 ^ n957 ;
  assign n1016 = n1015 ^ x4 ;
  assign n1017 = ~n888 & n1016 ;
  assign n1018 = n1017 ^ n888 ;
  assign n1019 = ~n887 & n1018 ;
  assign n1020 = x7 & x9 ;
  assign n1021 = ~x0 & n909 ;
  assign n1022 = n1020 & n1021 ;
  assign n1023 = n742 & n1022 ;
  assign n1024 = x2 & ~n1023 ;
  assign n1025 = ~n295 & ~n1024 ;
  assign n1026 = ~n1019 & ~n1025 ;
  assign n1027 = ~x1 & x4 ;
  assign n1028 = ~x14 & n129 ;
  assign n1029 = n892 & n1028 ;
  assign n1030 = ~n246 & n1029 ;
  assign n1031 = n477 & n655 ;
  assign n1032 = n1031 ^ x7 ;
  assign n1033 = n215 & n384 ;
  assign n1034 = ~n540 & ~n1033 ;
  assign n1035 = n1034 ^ x0 ;
  assign n1036 = n1035 ^ n1034 ;
  assign n1037 = ~x12 & n195 ;
  assign n1038 = ~n191 & ~n1037 ;
  assign n1039 = n1038 ^ n1034 ;
  assign n1040 = ~n1036 & n1039 ;
  assign n1041 = n1040 ^ n1034 ;
  assign n1042 = n1041 ^ n1031 ;
  assign n1043 = ~n1032 & n1042 ;
  assign n1044 = n1043 ^ n1040 ;
  assign n1045 = n1044 ^ n1034 ;
  assign n1046 = n1045 ^ x7 ;
  assign n1047 = ~n1031 & ~n1046 ;
  assign n1048 = n1047 ^ n1031 ;
  assign n1049 = n1048 ^ n1031 ;
  assign n1050 = n701 & ~n1049 ;
  assign n1051 = ~n338 & ~n466 ;
  assign n1052 = ~x12 & ~n1051 ;
  assign n1053 = n105 & n1052 ;
  assign n1054 = ~n1050 & ~n1053 ;
  assign n1055 = ~n1030 & n1054 ;
  assign n1056 = n1055 ^ x13 ;
  assign n1057 = n1056 ^ n1055 ;
  assign n1058 = x0 & ~n1051 ;
  assign n1059 = ~x0 & n503 ;
  assign n1060 = n522 & n1059 ;
  assign n1061 = ~n1058 & ~n1060 ;
  assign n1062 = x5 & ~n1061 ;
  assign n1063 = n149 & n794 ;
  assign n1064 = ~n1062 & ~n1063 ;
  assign n1065 = n39 & ~n1064 ;
  assign n1066 = n195 & n684 ;
  assign n1067 = ~n1065 & ~n1066 ;
  assign n1068 = n1067 ^ n1055 ;
  assign n1069 = n1057 & n1068 ;
  assign n1070 = n1069 ^ n1055 ;
  assign n1071 = x15 & ~n1070 ;
  assign n1072 = n1027 & n1071 ;
  assign n1073 = x0 & ~x4 ;
  assign n1074 = n361 & n690 ;
  assign n1075 = n309 & n566 ;
  assign n1076 = ~n1074 & ~n1075 ;
  assign n1077 = n1073 & ~n1076 ;
  assign n1078 = ~x4 & ~x14 ;
  assign n1079 = ~x3 & n1078 ;
  assign n1080 = n21 & n373 ;
  assign n1081 = ~n134 & n1080 ;
  assign n1082 = n426 ^ x0 ;
  assign n1083 = n1082 ^ n426 ;
  assign n1084 = x1 & ~x13 ;
  assign n1085 = ~n817 & ~n1084 ;
  assign n1086 = ~n337 & n1085 ;
  assign n1087 = n1086 ^ n426 ;
  assign n1088 = n1083 & n1087 ;
  assign n1089 = n1088 ^ n426 ;
  assign n1090 = n859 & n1089 ;
  assign n1091 = ~n1081 & ~n1090 ;
  assign n1092 = n1079 & ~n1091 ;
  assign n1093 = x9 ^ x4 ;
  assign n1094 = n259 ^ n88 ;
  assign n1095 = n259 ^ x9 ;
  assign n1096 = n1095 ^ n259 ;
  assign n1097 = n1094 & ~n1096 ;
  assign n1098 = n1097 ^ n259 ;
  assign n1099 = ~n1093 & n1098 ;
  assign n1100 = n309 & n1099 ;
  assign n1101 = n354 & n1020 ;
  assign n1102 = n222 & n259 ;
  assign n1103 = n1101 & n1102 ;
  assign n1104 = ~n1100 & ~n1103 ;
  assign n1105 = x0 & ~n1104 ;
  assign n1106 = n222 & n816 ;
  assign n1107 = n89 & n466 ;
  assign n1108 = n1106 & n1107 ;
  assign n1109 = ~n1105 & ~n1108 ;
  assign n1110 = ~n87 & ~n1109 ;
  assign n1111 = ~x7 & n149 ;
  assign n1112 = ~x4 & n77 ;
  assign n1113 = ~x1 & n34 ;
  assign n1114 = ~n134 & n1113 ;
  assign n1115 = ~n572 & ~n1114 ;
  assign n1116 = n1112 & ~n1115 ;
  assign n1117 = n1111 & n1116 ;
  assign n1118 = ~n1110 & ~n1117 ;
  assign n1119 = ~n1092 & n1118 ;
  assign n1120 = ~n1077 & n1119 ;
  assign n1121 = x15 & ~n1120 ;
  assign n1122 = n216 & n999 ;
  assign n1123 = ~x4 & x5 ;
  assign n1124 = ~x9 & n1123 ;
  assign n1125 = ~x3 & ~x13 ;
  assign n1126 = n99 & ~n1125 ;
  assign n1127 = n927 & n933 ;
  assign n1128 = ~n308 & ~n1127 ;
  assign n1129 = ~n1126 & n1128 ;
  assign n1130 = n1124 & ~n1129 ;
  assign n1131 = ~n1122 & ~n1130 ;
  assign n1132 = n148 & ~n1131 ;
  assign n1133 = ~x2 & ~n1132 ;
  assign n1134 = n701 & n829 ;
  assign n1135 = ~n764 & ~n1134 ;
  assign n1136 = n429 & ~n1135 ;
  assign n1137 = x0 & n466 ;
  assign n1138 = ~x5 & x13 ;
  assign n1139 = ~n717 & ~n1138 ;
  assign n1140 = n1137 & ~n1139 ;
  assign n1141 = ~n61 & ~n639 ;
  assign n1142 = n453 & ~n1141 ;
  assign n1143 = ~n1140 & ~n1142 ;
  assign n1144 = ~n1136 & n1143 ;
  assign n1145 = n610 & ~n1144 ;
  assign n1146 = n29 & n684 ;
  assign n1147 = n38 & n1146 ;
  assign n1148 = ~n1145 & ~n1147 ;
  assign n1149 = n88 & ~n1051 ;
  assign n1150 = x5 & x14 ;
  assign n1151 = ~n640 & ~n1150 ;
  assign n1152 = n307 & n1151 ;
  assign n1153 = n1149 & n1152 ;
  assign n1154 = x14 ^ x7 ;
  assign n1155 = n107 ^ x14 ;
  assign n1156 = n1155 ^ n107 ;
  assign n1157 = n107 ^ n104 ;
  assign n1158 = ~n1156 & n1157 ;
  assign n1159 = n1158 ^ n107 ;
  assign n1160 = ~n1154 & n1159 ;
  assign n1161 = ~n505 & n1160 ;
  assign n1162 = ~n1153 & ~n1161 ;
  assign n1163 = n343 & ~n1162 ;
  assign n1164 = ~x7 & n153 ;
  assign n1165 = n282 & n656 ;
  assign n1166 = ~n647 & ~n1165 ;
  assign n1167 = n100 & ~n1166 ;
  assign n1168 = ~n1164 & n1167 ;
  assign n1169 = n566 & n640 ;
  assign n1170 = n117 & n1169 ;
  assign n1171 = x15 & n1170 ;
  assign n1172 = ~n1168 & ~n1171 ;
  assign n1173 = ~n1163 & n1172 ;
  assign n1174 = n166 & n361 ;
  assign n1175 = n434 & n549 ;
  assign n1176 = n282 & n1175 ;
  assign n1177 = ~x14 & n133 ;
  assign n1178 = n148 & n1177 ;
  assign n1179 = n118 & n1178 ;
  assign n1180 = n399 & n693 ;
  assign n1181 = n434 & n1180 ;
  assign n1182 = ~n1179 & ~n1181 ;
  assign n1183 = ~n1176 & n1182 ;
  assign n1184 = n1183 ^ x3 ;
  assign n1185 = n1184 ^ n1183 ;
  assign n1186 = n1185 ^ n1174 ;
  assign n1187 = n109 & n429 ;
  assign n1188 = x7 & ~n132 ;
  assign n1189 = x7 & n99 ;
  assign n1190 = ~n1188 & ~n1189 ;
  assign n1191 = n701 & n933 ;
  assign n1192 = x0 & ~n110 ;
  assign n1193 = ~n1191 & n1192 ;
  assign n1194 = ~n1190 & ~n1193 ;
  assign n1195 = ~n1187 & ~n1194 ;
  assign n1196 = n1195 ^ x9 ;
  assign n1197 = ~x9 & n1196 ;
  assign n1198 = n1197 ^ n1183 ;
  assign n1199 = n1198 ^ x9 ;
  assign n1200 = ~n1186 & n1199 ;
  assign n1201 = n1200 ^ n1197 ;
  assign n1202 = n1201 ^ x9 ;
  assign n1203 = ~n1174 & ~n1202 ;
  assign n1204 = n1203 ^ n1174 ;
  assign n1205 = n1173 & ~n1204 ;
  assign n1206 = n1148 & n1205 ;
  assign n1207 = x1 & ~n1206 ;
  assign n1208 = n49 & n640 ;
  assign n1209 = n539 & n1208 ;
  assign n1210 = ~n524 & ~n1209 ;
  assign n1211 = ~x3 & n434 ;
  assign n1212 = ~n1052 & ~n1211 ;
  assign n1213 = x13 & ~n1212 ;
  assign n1214 = ~x5 & x12 ;
  assign n1215 = n522 & ~n1214 ;
  assign n1216 = ~n1213 & ~n1215 ;
  assign n1217 = n1113 & ~n1216 ;
  assign n1218 = x0 & n1217 ;
  assign n1219 = n520 & n863 ;
  assign n1220 = n101 & n1219 ;
  assign n1221 = ~n1218 & ~n1220 ;
  assign n1222 = n1210 & n1221 ;
  assign n1223 = ~n1207 & n1222 ;
  assign n1224 = x4 & ~n1223 ;
  assign n1225 = n1133 & ~n1224 ;
  assign n1226 = ~n1121 & n1225 ;
  assign n1227 = ~n1072 & n1226 ;
  assign n1228 = ~n1026 & ~n1227 ;
  assign n1229 = ~n98 & ~n434 ;
  assign n1230 = ~x4 & ~x7 ;
  assign n1231 = ~x5 & ~x12 ;
  assign n1232 = ~n1230 & ~n1231 ;
  assign n1233 = n450 & ~n1232 ;
  assign n1234 = x4 & x12 ;
  assign n1235 = n189 & n1234 ;
  assign n1236 = n104 & n1235 ;
  assign n1237 = ~n1233 & ~n1236 ;
  assign n1238 = n922 & ~n1237 ;
  assign n1239 = ~n1229 & n1238 ;
  assign n1240 = ~n1228 & ~n1239 ;
  assign n1241 = n1240 ^ n809 ;
  assign n1242 = ~n811 & n1241 ;
  assign n1243 = n1242 ^ n809 ;
  assign n1244 = n449 & n1243 ;
  assign n1245 = n19 & ~n1244 ;
  assign n1246 = ~x2 & ~x3 ;
  assign n1247 = n450 & n1246 ;
  assign n1248 = ~x0 & x2 ;
  assign n1249 = x3 & n1248 ;
  assign n1250 = ~x1 & n1249 ;
  assign n1251 = ~n1247 & ~n1250 ;
  assign n1252 = ~x8 & x9 ;
  assign n1253 = ~n88 & ~n259 ;
  assign n1254 = ~x5 & ~x6 ;
  assign n1255 = n1230 & n1254 ;
  assign n1256 = x10 & x12 ;
  assign n1257 = x14 & n1256 ;
  assign n1258 = n1255 & n1257 ;
  assign n1259 = ~x10 & ~n399 ;
  assign n1260 = x6 & ~x12 ;
  assign n1261 = ~x4 & ~x5 ;
  assign n1262 = n1260 & n1261 ;
  assign n1263 = n1259 & n1262 ;
  assign n1264 = x4 & ~x10 ;
  assign n1265 = ~x12 & n1264 ;
  assign n1266 = ~x5 & x14 ;
  assign n1267 = ~x6 & ~x7 ;
  assign n1268 = ~n1266 & n1267 ;
  assign n1269 = n1265 & n1268 ;
  assign n1270 = ~n1263 & ~n1269 ;
  assign n1271 = ~n1258 & n1270 ;
  assign n1272 = ~n1253 & ~n1271 ;
  assign n1273 = x6 & x7 ;
  assign n1274 = n250 & ~n1273 ;
  assign n1275 = ~x10 & n731 ;
  assign n1276 = ~x6 & x7 ;
  assign n1277 = ~n291 & ~n1276 ;
  assign n1278 = n1275 & ~n1277 ;
  assign n1279 = n74 & n1278 ;
  assign n1280 = ~n1274 & n1279 ;
  assign n1281 = ~n1272 & ~n1280 ;
  assign n1282 = x15 & ~n1281 ;
  assign n1283 = ~x6 & x10 ;
  assign n1284 = n222 & n1283 ;
  assign n1285 = x6 & x10 ;
  assign n1286 = ~x4 & n1285 ;
  assign n1287 = x7 & n1286 ;
  assign n1288 = ~n1284 & ~n1287 ;
  assign n1289 = n933 & ~n1288 ;
  assign n1290 = x5 & x6 ;
  assign n1291 = n1230 & n1290 ;
  assign n1292 = n98 & n1254 ;
  assign n1293 = ~n1291 & ~n1292 ;
  assign n1294 = ~x10 & x11 ;
  assign n1295 = ~n109 & ~n1294 ;
  assign n1296 = ~n1293 & ~n1295 ;
  assign n1297 = ~n1289 & ~n1296 ;
  assign n1298 = ~x6 & ~x12 ;
  assign n1299 = n294 & n1298 ;
  assign n1300 = x10 & ~x11 ;
  assign n1301 = ~n1294 & ~n1300 ;
  assign n1302 = n1299 & ~n1301 ;
  assign n1303 = x10 & x13 ;
  assign n1304 = ~n215 & ~n1303 ;
  assign n1305 = x6 & ~n909 ;
  assign n1306 = ~n1304 & n1305 ;
  assign n1307 = ~n1302 & ~n1306 ;
  assign n1308 = n1230 & ~n1307 ;
  assign n1309 = ~x10 & x13 ;
  assign n1310 = x13 & ~n87 ;
  assign n1311 = ~n1309 & ~n1310 ;
  assign n1312 = x6 & ~x7 ;
  assign n1313 = n53 & n1312 ;
  assign n1314 = ~n1311 & n1313 ;
  assign n1315 = ~n1308 & ~n1314 ;
  assign n1316 = ~x10 & ~x11 ;
  assign n1317 = n753 & n1316 ;
  assign n1318 = n1276 & n1317 ;
  assign n1319 = x4 & n1318 ;
  assign n1320 = x4 & ~x7 ;
  assign n1321 = n88 & n1283 ;
  assign n1322 = ~n277 & ~n1260 ;
  assign n1323 = n259 & ~n1322 ;
  assign n1324 = ~n1321 & ~n1323 ;
  assign n1325 = n1320 & ~n1324 ;
  assign n1326 = ~n1319 & ~n1325 ;
  assign n1327 = n1315 & n1326 ;
  assign n1328 = n190 & ~n1327 ;
  assign n1329 = n1297 & ~n1328 ;
  assign n1330 = x4 & ~x12 ;
  assign n1331 = ~n1273 & ~n1330 ;
  assign n1332 = ~x5 & ~x10 ;
  assign n1333 = ~n587 & n909 ;
  assign n1334 = n1332 & n1333 ;
  assign n1335 = ~n1331 & n1334 ;
  assign n1336 = x6 & ~n99 ;
  assign n1337 = ~n88 & ~n1336 ;
  assign n1338 = n98 & ~n1337 ;
  assign n1339 = n394 & n910 ;
  assign n1340 = ~x4 & x7 ;
  assign n1341 = x11 ^ x6 ;
  assign n1342 = n1341 ^ x11 ;
  assign n1343 = n88 ^ x11 ;
  assign n1344 = n1342 & n1343 ;
  assign n1345 = n1344 ^ x11 ;
  assign n1346 = n1340 & n1345 ;
  assign n1347 = ~n1339 & ~n1346 ;
  assign n1348 = ~n1338 & n1347 ;
  assign n1349 = n1348 ^ x10 ;
  assign n1350 = n1349 ^ n1348 ;
  assign n1351 = n1350 ^ x5 ;
  assign n1352 = ~n291 & ~n394 ;
  assign n1353 = n1352 ^ x7 ;
  assign n1354 = n1352 & n1353 ;
  assign n1355 = n1354 ^ n1348 ;
  assign n1356 = n1355 ^ n1352 ;
  assign n1357 = n1351 & ~n1356 ;
  assign n1358 = n1357 ^ n1354 ;
  assign n1359 = n1358 ^ n1352 ;
  assign n1360 = x5 & n1359 ;
  assign n1361 = ~n1335 & ~n1360 ;
  assign n1362 = n1329 & n1361 ;
  assign n1363 = ~n1282 & n1362 ;
  assign n1364 = n1252 & ~n1363 ;
  assign n1365 = x8 & ~x12 ;
  assign n1366 = ~x9 & x13 ;
  assign n1367 = n1365 & n1366 ;
  assign n1368 = ~x13 & n603 ;
  assign n1369 = ~x8 & n1368 ;
  assign n1370 = ~n1367 & ~n1369 ;
  assign n1371 = n33 & ~n1370 ;
  assign n1372 = x11 ^ x10 ;
  assign n1373 = n1293 ^ x11 ;
  assign n1374 = n1373 ^ n1293 ;
  assign n1375 = n1374 ^ n1372 ;
  assign n1376 = ~n249 & ~n252 ;
  assign n1377 = n1376 ^ n22 ;
  assign n1378 = n22 & ~n1377 ;
  assign n1379 = n1378 ^ n1293 ;
  assign n1380 = n1379 ^ n22 ;
  assign n1381 = n1375 & ~n1380 ;
  assign n1382 = n1381 ^ n1378 ;
  assign n1383 = n1382 ^ n22 ;
  assign n1384 = n1372 & n1383 ;
  assign n1385 = n1371 & n1384 ;
  assign n1386 = ~n43 & ~n1370 ;
  assign n1387 = n25 & ~n1352 ;
  assign n1388 = n1300 & n1387 ;
  assign n1389 = n1386 & n1388 ;
  assign n1390 = ~x8 & n1309 ;
  assign n1391 = n222 & n1312 ;
  assign n1392 = n1390 & n1391 ;
  assign n1393 = n215 & n1392 ;
  assign n1394 = x8 & x12 ;
  assign n1395 = x13 & n1394 ;
  assign n1396 = ~x9 & n1395 ;
  assign n1397 = ~x6 & n222 ;
  assign n1398 = ~n1301 & n1397 ;
  assign n1399 = n1396 & n1398 ;
  assign n1400 = ~n1393 & ~n1399 ;
  assign n1401 = ~n1389 & n1400 ;
  assign n1402 = ~n1385 & n1401 ;
  assign n1403 = ~n1364 & n1402 ;
  assign n1404 = x8 & x9 ;
  assign n1405 = x10 & x11 ;
  assign n1406 = n22 & n1405 ;
  assign n1407 = n25 & n1316 ;
  assign n1408 = ~n1406 & ~n1407 ;
  assign n1409 = ~n153 & n1376 ;
  assign n1410 = ~n1408 & n1409 ;
  assign n1411 = n22 & n252 ;
  assign n1412 = n38 & n1294 ;
  assign n1413 = n1411 & n1412 ;
  assign n1414 = n1123 & n1276 ;
  assign n1415 = x10 & ~x13 ;
  assign n1416 = n314 & n1415 ;
  assign n1417 = n1414 & n1416 ;
  assign n1418 = ~n1413 & ~n1417 ;
  assign n1419 = ~n43 & ~n1418 ;
  assign n1433 = x4 & x14 ;
  assign n1434 = n1352 & ~n1433 ;
  assign n1435 = x10 & ~x12 ;
  assign n1436 = ~n284 & n1435 ;
  assign n1437 = ~n1434 & n1436 ;
  assign n1440 = x6 & ~x10 ;
  assign n1438 = ~x4 & ~x12 ;
  assign n1439 = n528 & ~n1438 ;
  assign n1441 = n1440 ^ n1439 ;
  assign n1442 = n1441 ^ n1437 ;
  assign n1443 = x4 & n277 ;
  assign n1444 = n1443 ^ n120 ;
  assign n1445 = ~n1440 & ~n1444 ;
  assign n1446 = n1445 ^ n120 ;
  assign n1447 = ~n1442 & ~n1446 ;
  assign n1448 = n1447 ^ n1445 ;
  assign n1449 = n1448 ^ n120 ;
  assign n1450 = n1449 ^ n1440 ;
  assign n1451 = ~n1437 & n1450 ;
  assign n1452 = n190 & ~n1451 ;
  assign n1427 = n475 & n1123 ;
  assign n1453 = n267 & n1427 ;
  assign n1454 = ~x13 & n42 ;
  assign n1455 = n1261 & n1454 ;
  assign n1456 = x4 & ~x5 ;
  assign n1457 = ~x4 & ~x13 ;
  assign n1458 = ~n1456 & ~n1457 ;
  assign n1459 = ~n1352 & n1458 ;
  assign n1460 = ~n1455 & ~n1459 ;
  assign n1461 = ~n1453 & n1460 ;
  assign n1462 = n1256 & ~n1461 ;
  assign n1463 = ~n1452 & ~n1462 ;
  assign n1464 = ~x11 & ~n1463 ;
  assign n1420 = ~x4 & x12 ;
  assign n1421 = n1321 & n1420 ;
  assign n1422 = ~x5 & ~n314 ;
  assign n1423 = n1286 & ~n1422 ;
  assign n1424 = ~n1421 & ~n1423 ;
  assign n1425 = n53 & n1283 ;
  assign n1426 = n334 & n1425 ;
  assign n1428 = n1298 & n1316 ;
  assign n1429 = n1427 & n1428 ;
  assign n1430 = ~n1426 & ~n1429 ;
  assign n1431 = ~n1284 & n1430 ;
  assign n1432 = n1424 & n1431 ;
  assign n1465 = n1464 ^ n1432 ;
  assign n1466 = n1465 ^ n1432 ;
  assign n1467 = ~x10 & x15 ;
  assign n1468 = ~x12 & n1467 ;
  assign n1469 = ~n1256 & ~n1468 ;
  assign n1470 = n909 & n1254 ;
  assign n1471 = ~x4 & n1470 ;
  assign n1472 = ~n1469 & n1471 ;
  assign n1473 = n1472 ^ n1432 ;
  assign n1474 = n1473 ^ n1432 ;
  assign n1475 = ~n1466 & ~n1474 ;
  assign n1476 = n1475 ^ n1432 ;
  assign n1477 = ~x7 & n1476 ;
  assign n1478 = n1477 ^ n1432 ;
  assign n1479 = ~n1419 & n1478 ;
  assign n1480 = ~n1410 & n1479 ;
  assign n1481 = n1404 & ~n1480 ;
  assign n1482 = ~x7 & ~x9 ;
  assign n1483 = x12 & n17 ;
  assign n1484 = x13 & n291 ;
  assign n1485 = n1275 & n1484 ;
  assign n1486 = ~n1483 & ~n1485 ;
  assign n1487 = x11 & ~n1486 ;
  assign n1488 = n1459 & n1487 ;
  assign n1489 = x10 & x14 ;
  assign n1490 = ~n194 & ~n1138 ;
  assign n1491 = n394 & ~n1490 ;
  assign n1492 = x5 & ~x6 ;
  assign n1493 = x8 & x13 ;
  assign n1494 = ~x4 & n1493 ;
  assign n1495 = ~n1492 & n1494 ;
  assign n1496 = ~n1491 & ~n1495 ;
  assign n1497 = x12 & ~n1496 ;
  assign n1498 = ~x13 & n1365 ;
  assign n1499 = n1397 & n1498 ;
  assign n1500 = ~n1497 & ~n1499 ;
  assign n1501 = n1489 & ~n1500 ;
  assign n1502 = x5 & ~x10 ;
  assign n1503 = x6 & ~x8 ;
  assign n1504 = ~x4 & n1503 ;
  assign n1505 = n717 & n1504 ;
  assign n1506 = x4 & x8 ;
  assign n1507 = x14 & n1506 ;
  assign n1508 = n133 & n1507 ;
  assign n1509 = ~n1505 & ~n1508 ;
  assign n1510 = n1502 & ~n1509 ;
  assign n1511 = ~x12 & n1493 ;
  assign n1512 = n1284 & n1511 ;
  assign n1513 = ~n1510 & ~n1512 ;
  assign n1514 = ~n1501 & n1513 ;
  assign n1515 = n1514 ^ x11 ;
  assign n1516 = n1515 ^ n1514 ;
  assign n1517 = n1516 ^ x15 ;
  assign n1518 = ~x5 & x8 ;
  assign n1519 = n1309 & n1518 ;
  assign n1520 = n17 & ~n284 ;
  assign n1521 = ~x13 & n434 ;
  assign n1522 = ~n1231 & ~n1521 ;
  assign n1523 = n1520 & ~n1522 ;
  assign n1524 = ~n1519 & ~n1523 ;
  assign n1525 = n291 & ~n1524 ;
  assign n1526 = ~x5 & n38 ;
  assign n1527 = ~n194 & ~n1526 ;
  assign n1528 = ~x8 & ~x12 ;
  assign n1529 = ~n1394 & ~n1528 ;
  assign n1530 = ~x10 & ~x14 ;
  assign n1531 = n291 & n1530 ;
  assign n1532 = ~n1529 & n1531 ;
  assign n1533 = ~n1527 & n1532 ;
  assign n1534 = n18 & n38 ;
  assign n1535 = n1397 & n1534 ;
  assign n1536 = ~n1533 & ~n1535 ;
  assign n1537 = ~n1525 & n1536 ;
  assign n1538 = ~n119 & ~n1457 ;
  assign n1539 = ~n1493 & ~n1528 ;
  assign n1540 = ~x6 & n1539 ;
  assign n1541 = n1538 & n1540 ;
  assign n1542 = ~x4 & n133 ;
  assign n1543 = x8 & n1542 ;
  assign n1544 = ~n1541 & ~n1543 ;
  assign n1545 = n1489 & ~n1544 ;
  assign n1546 = ~x8 & ~n86 ;
  assign n1547 = ~x6 & ~n1546 ;
  assign n1548 = ~x10 & n119 ;
  assign n1549 = n1547 & n1548 ;
  assign n1550 = ~x8 & x13 ;
  assign n1551 = ~x10 & ~x12 ;
  assign n1552 = ~x10 & ~x13 ;
  assign n1553 = x14 & ~n1552 ;
  assign n1554 = ~n1551 & n1553 ;
  assign n1555 = ~n1550 & ~n1554 ;
  assign n1556 = n252 & ~n1555 ;
  assign n1557 = ~n1256 & n1556 ;
  assign n1558 = ~n1549 & ~n1557 ;
  assign n1559 = x13 & n1435 ;
  assign n1560 = ~x6 & n1506 ;
  assign n1561 = n1559 & n1560 ;
  assign n1562 = ~x8 & x10 ;
  assign n1563 = n403 & n528 ;
  assign n1564 = n1562 & n1563 ;
  assign n1565 = ~n1561 & ~n1564 ;
  assign n1566 = n1558 & n1565 ;
  assign n1567 = ~n1545 & n1566 ;
  assign n1568 = ~x5 & ~n1567 ;
  assign n1569 = n1568 ^ n1537 ;
  assign n1570 = n1537 & ~n1569 ;
  assign n1571 = n1570 ^ n1514 ;
  assign n1572 = n1571 ^ n1537 ;
  assign n1573 = n1517 & n1572 ;
  assign n1574 = n1573 ^ n1570 ;
  assign n1575 = n1574 ^ n1537 ;
  assign n1576 = x15 & n1575 ;
  assign n1577 = n1576 ^ x15 ;
  assign n1578 = ~n1488 & ~n1577 ;
  assign n1579 = n1482 & ~n1578 ;
  assign n1580 = ~n1481 & ~n1579 ;
  assign n1581 = ~x4 & x8 ;
  assign n1582 = ~x6 & x13 ;
  assign n1583 = ~x5 & x6 ;
  assign n1584 = ~n1582 & ~n1583 ;
  assign n1585 = n215 & ~n1584 ;
  assign n1586 = x6 & ~x11 ;
  assign n1587 = ~x5 & n1586 ;
  assign n1588 = ~x12 & x15 ;
  assign n1589 = ~n284 & n1588 ;
  assign n1590 = n1587 & n1589 ;
  assign n1591 = ~n1585 & ~n1590 ;
  assign n1592 = n1581 & ~n1591 ;
  assign n1593 = n1542 & n1587 ;
  assign n1594 = n42 & n1593 ;
  assign n1595 = ~n1592 & ~n1594 ;
  assign n1596 = x10 & ~n1595 ;
  assign n1597 = x5 & x10 ;
  assign n1598 = ~x8 & x12 ;
  assign n1599 = ~x8 & ~x11 ;
  assign n1600 = ~x6 & ~n1599 ;
  assign n1601 = ~n1598 & ~n1600 ;
  assign n1602 = x8 & ~n503 ;
  assign n1603 = ~x4 & ~n215 ;
  assign n1604 = n475 & n1603 ;
  assign n1605 = ~n1602 & n1604 ;
  assign n1606 = ~n1601 & n1605 ;
  assign n1607 = x15 & n62 ;
  assign n1608 = x8 & ~x13 ;
  assign n1609 = ~x11 & n1608 ;
  assign n1610 = n1607 & n1609 ;
  assign n1611 = ~x8 & x11 ;
  assign n1612 = ~n153 & n1611 ;
  assign n1613 = ~n1610 & ~n1612 ;
  assign n1614 = ~n1352 & ~n1613 ;
  assign n1615 = ~n1606 & ~n1614 ;
  assign n1616 = n1597 & ~n1615 ;
  assign n1617 = ~n1596 & ~n1616 ;
  assign n1618 = ~x6 & x15 ;
  assign n1619 = x4 & ~x8 ;
  assign n1620 = n1551 & n1619 ;
  assign n1621 = x5 & n1620 ;
  assign n1622 = ~n1123 & ~n1456 ;
  assign n1623 = ~x12 & n18 ;
  assign n1624 = ~n1483 & ~n1623 ;
  assign n1625 = ~n87 & ~n1624 ;
  assign n1626 = ~n1622 & n1625 ;
  assign n1627 = ~n1621 & ~n1626 ;
  assign n1628 = n1618 & ~n1627 ;
  assign n1629 = n249 & n1256 ;
  assign n1630 = x5 & x8 ;
  assign n1631 = ~x14 & n1630 ;
  assign n1632 = n1629 & n1631 ;
  assign n1633 = ~x8 & x15 ;
  assign n1634 = ~x4 & n1290 ;
  assign n1635 = n1551 & n1634 ;
  assign n1636 = n1633 & n1635 ;
  assign n1637 = ~n1632 & ~n1636 ;
  assign n1638 = ~n1628 & n1637 ;
  assign n1639 = ~n1253 & ~n1638 ;
  assign n1640 = x15 & n1550 ;
  assign n1641 = n1262 & n1640 ;
  assign n1642 = ~x6 & x8 ;
  assign n1643 = ~x4 & n1642 ;
  assign n1644 = ~x8 & n252 ;
  assign n1645 = ~n153 & n1644 ;
  assign n1646 = ~n476 & n1394 ;
  assign n1647 = ~n1550 & ~n1646 ;
  assign n1648 = ~n1352 & ~n1647 ;
  assign n1649 = ~n1645 & ~n1648 ;
  assign n1650 = ~n1643 & n1649 ;
  assign n1651 = x5 & ~n1650 ;
  assign n1652 = ~x4 & n1394 ;
  assign n1653 = ~n1456 & ~n1652 ;
  assign n1654 = x13 & n1322 ;
  assign n1655 = ~n1653 & n1654 ;
  assign n1656 = n277 & n284 ;
  assign n1657 = x8 & x15 ;
  assign n1658 = n1456 & n1657 ;
  assign n1659 = n1656 & n1658 ;
  assign n1660 = ~n1655 & ~n1659 ;
  assign n1661 = ~n1651 & n1660 ;
  assign n1662 = ~n1641 & n1661 ;
  assign n1663 = n1294 & ~n1662 ;
  assign n1664 = ~n1639 & ~n1663 ;
  assign n1665 = ~x8 & n249 ;
  assign n1666 = n49 & n1665 ;
  assign n1667 = x8 & ~x14 ;
  assign n1668 = n249 & n1667 ;
  assign n1669 = x6 & x8 ;
  assign n1670 = ~x4 & n1669 ;
  assign n1671 = ~x6 & ~x8 ;
  assign n1672 = ~n1669 & ~n1671 ;
  assign n1673 = x4 & n1672 ;
  assign n1674 = ~n1670 & ~n1673 ;
  assign n1675 = x14 & ~n1674 ;
  assign n1676 = ~n1668 & ~n1675 ;
  assign n1677 = n153 & ~n1676 ;
  assign n1678 = ~n1666 & ~n1677 ;
  assign n1679 = x15 & ~n1678 ;
  assign n1680 = n252 & n1511 ;
  assign n1681 = ~n1679 & ~n1680 ;
  assign n1682 = n1681 ^ n42 ;
  assign n1683 = n1682 ^ n1681 ;
  assign n1684 = n133 & n1669 ;
  assign n1685 = n1684 ^ n1681 ;
  assign n1686 = n1685 ^ n1681 ;
  assign n1687 = n1683 & n1686 ;
  assign n1688 = n1687 ^ n1681 ;
  assign n1689 = ~x5 & ~n1688 ;
  assign n1690 = n1689 ^ n1681 ;
  assign n1691 = n1316 & ~n1690 ;
  assign n1692 = n1664 & ~n1691 ;
  assign n1693 = n1617 & n1692 ;
  assign n1694 = n264 & ~n1693 ;
  assign n1695 = n1580 & ~n1694 ;
  assign n1696 = n1403 & n1695 ;
  assign n1697 = ~n1251 & ~n1696 ;
  assign n1698 = ~n1365 & ~n1598 ;
  assign n1699 = ~x9 & n259 ;
  assign n1700 = ~n1489 & ~n1530 ;
  assign n1701 = n354 & ~n1700 ;
  assign n1702 = x0 & x2 ;
  assign n1703 = ~x10 & n1702 ;
  assign n1704 = ~n210 & ~n1703 ;
  assign n1705 = n1701 & ~n1704 ;
  assign n1706 = ~x10 & x14 ;
  assign n1707 = n1702 & n1706 ;
  assign n1708 = x10 & ~x14 ;
  assign n1709 = n210 & n1708 ;
  assign n1710 = ~n1707 & ~n1709 ;
  assign n1711 = ~n558 & ~n1710 ;
  assign n1712 = ~n1705 & ~n1711 ;
  assign n1713 = n1699 & ~n1712 ;
  assign n1714 = n214 & n354 ;
  assign n1715 = x0 & ~x2 ;
  assign n1716 = ~n1248 & ~n1715 ;
  assign n1717 = ~n1700 & ~n1716 ;
  assign n1719 = x2 & x10 ;
  assign n1718 = ~x2 & ~x10 ;
  assign n1720 = n1719 ^ n1718 ;
  assign n1721 = ~x0 & n1720 ;
  assign n1722 = n1721 ^ n1719 ;
  assign n1723 = ~n1717 & ~n1722 ;
  assign n1724 = n1714 & ~n1723 ;
  assign n1725 = ~x11 & n1724 ;
  assign n1726 = ~n1713 & ~n1725 ;
  assign n1727 = n25 & ~n1726 ;
  assign n1728 = ~x9 & x11 ;
  assign n1729 = n1084 & n1728 ;
  assign n1730 = ~n1722 & n1729 ;
  assign n1731 = ~x11 & n214 ;
  assign n1733 = ~x0 & ~x10 ;
  assign n1732 = x0 & x10 ;
  assign n1734 = n1733 ^ n1732 ;
  assign n1735 = x14 ^ x2 ;
  assign n1736 = n1732 ^ x14 ;
  assign n1737 = n1735 & n1736 ;
  assign n1738 = n1737 ^ x14 ;
  assign n1739 = n1734 & ~n1738 ;
  assign n1740 = n1739 ^ n1733 ;
  assign n1741 = n1740 ^ n1717 ;
  assign n1742 = ~x1 & n1741 ;
  assign n1743 = n1742 ^ n1717 ;
  assign n1744 = n1731 & n1743 ;
  assign n1745 = ~n1730 & ~n1744 ;
  assign n1746 = x3 & ~n1745 ;
  assign n1747 = x0 & ~x10 ;
  assign n1748 = n292 & n1747 ;
  assign n1749 = n1248 & n1708 ;
  assign n1750 = ~n1748 & ~n1749 ;
  assign n1751 = n550 & n1731 ;
  assign n1752 = ~n1750 & n1751 ;
  assign n1753 = ~n1746 & ~n1752 ;
  assign n1754 = n22 & ~n1753 ;
  assign n1755 = ~n1727 & ~n1754 ;
  assign n1756 = ~n1352 & ~n1755 ;
  assign n1757 = x3 & ~n1716 ;
  assign n1758 = x9 & x10 ;
  assign n1759 = n88 & n1758 ;
  assign n1760 = ~x9 & ~x10 ;
  assign n1761 = n285 & n1760 ;
  assign n1762 = ~n1759 & ~n1761 ;
  assign n1763 = n252 & ~n1762 ;
  assign n1764 = n1699 & ~n1700 ;
  assign n1765 = ~x10 & n88 ;
  assign n1766 = x9 & n1765 ;
  assign n1767 = ~n1764 & ~n1766 ;
  assign n1768 = n249 & ~n1767 ;
  assign n1769 = ~n1763 & ~n1768 ;
  assign n1770 = n1757 & ~n1769 ;
  assign n1771 = n57 & n1770 ;
  assign n1772 = x4 & x10 ;
  assign n1773 = n217 & n1772 ;
  assign n1774 = n1246 & n1773 ;
  assign n1775 = x2 & ~x3 ;
  assign n1776 = n252 & n1706 ;
  assign n1777 = n25 & n1776 ;
  assign n1778 = n640 & n1283 ;
  assign n1779 = x7 & x10 ;
  assign n1780 = n1261 & n1779 ;
  assign n1781 = ~n1778 & ~n1780 ;
  assign n1782 = ~n1777 & n1781 ;
  assign n1783 = n1775 & ~n1782 ;
  assign n1784 = n249 & n1708 ;
  assign n1785 = ~n1776 & ~n1784 ;
  assign n1786 = ~x2 & x3 ;
  assign n1787 = ~x7 & n1786 ;
  assign n1788 = ~x5 & n1787 ;
  assign n1789 = ~n1785 & n1788 ;
  assign n1790 = ~x3 & x10 ;
  assign n1791 = n280 & n1790 ;
  assign n1792 = n1312 & n1791 ;
  assign n1793 = ~n1789 & ~n1792 ;
  assign n1794 = ~n1783 & n1793 ;
  assign n1795 = ~n1774 & n1794 ;
  assign n1796 = n21 & ~n1795 ;
  assign n1797 = ~x10 & n252 ;
  assign n1798 = n78 & n1797 ;
  assign n1799 = ~n1775 & ~n1786 ;
  assign n1800 = n918 & ~n1799 ;
  assign n1801 = x2 & ~x5 ;
  assign n1802 = n199 & n1801 ;
  assign n1803 = ~n1800 & ~n1802 ;
  assign n1804 = n1798 & ~n1803 ;
  assign n1805 = n1312 ^ n1276 ;
  assign n1806 = n1805 ^ n1312 ;
  assign n1807 = n1312 ^ n1078 ;
  assign n1808 = n1807 ^ n1312 ;
  assign n1809 = n1806 & n1808 ;
  assign n1810 = n1809 ^ n1312 ;
  assign n1811 = ~x3 & n1810 ;
  assign n1812 = n1811 ^ n1312 ;
  assign n1813 = n280 & n1812 ;
  assign n1814 = x2 & x7 ;
  assign n1815 = n249 & n1814 ;
  assign n1816 = n1028 & n1815 ;
  assign n1817 = ~n219 & ~n1816 ;
  assign n1818 = ~n1813 & n1817 ;
  assign n1819 = n816 & ~n1818 ;
  assign n1820 = x10 & n1819 ;
  assign n1821 = ~n1804 & ~n1820 ;
  assign n1822 = ~n22 & ~n1246 ;
  assign n1823 = x2 & x3 ;
  assign n1824 = ~n25 & ~n1823 ;
  assign n1825 = ~n1822 & ~n1824 ;
  assign n1826 = ~x14 & n249 ;
  assign n1827 = x1 & n1826 ;
  assign n1828 = n1825 & n1827 ;
  assign n1829 = n408 & n1775 ;
  assign n1830 = x4 & n1829 ;
  assign n1831 = ~n1787 & ~n1830 ;
  assign n1832 = ~x1 & n1492 ;
  assign n1833 = ~n1831 & n1832 ;
  assign n1834 = ~x2 & ~x5 ;
  assign n1835 = n1340 ^ n252 ;
  assign n1836 = n1835 ^ n1340 ;
  assign n1837 = n1340 ^ n399 ;
  assign n1838 = n1837 ^ n1340 ;
  assign n1839 = n1836 & n1838 ;
  assign n1840 = n1839 ^ n1340 ;
  assign n1841 = x1 & n1840 ;
  assign n1842 = n1841 ^ n1340 ;
  assign n1843 = n1834 & n1842 ;
  assign n1844 = x3 & n1843 ;
  assign n1845 = ~n1833 & ~n1844 ;
  assign n1846 = ~n1828 & n1845 ;
  assign n1847 = n1732 & ~n1846 ;
  assign n1848 = n1821 & ~n1847 ;
  assign n1849 = ~n1796 & n1848 ;
  assign n1850 = n1699 & ~n1849 ;
  assign n1851 = ~x14 & n1316 ;
  assign n1852 = n1714 & n1851 ;
  assign n1853 = ~n1759 & ~n1764 ;
  assign n1854 = n355 & ~n1853 ;
  assign n1855 = ~n1852 & ~n1854 ;
  assign n1856 = n1702 & ~n1855 ;
  assign n1857 = ~x0 & n396 ;
  assign n1858 = n829 & n1728 ;
  assign n1859 = ~x3 & n1758 ;
  assign n1860 = n88 & n1859 ;
  assign n1861 = ~x14 & n1860 ;
  assign n1862 = ~n1858 & ~n1861 ;
  assign n1863 = n1857 & ~n1862 ;
  assign n1864 = n88 & n384 ;
  assign n1865 = ~n1858 & ~n1864 ;
  assign n1866 = x10 & n926 ;
  assign n1867 = ~n1865 & n1866 ;
  assign n1868 = n550 & n1699 ;
  assign n1869 = ~n1867 & ~n1868 ;
  assign n1870 = n1715 & ~n1869 ;
  assign n1871 = ~x3 & n1729 ;
  assign n1872 = n1749 & n1871 ;
  assign n1873 = ~n1870 & ~n1872 ;
  assign n1874 = ~n1863 & n1873 ;
  assign n1875 = ~n1856 & n1874 ;
  assign n1876 = ~n1293 & ~n1875 ;
  assign n1877 = n210 & n253 ;
  assign n1878 = n1285 & n1877 ;
  assign n1879 = n249 & n1707 ;
  assign n1880 = ~n1878 & ~n1879 ;
  assign n1886 = ~x5 & n721 ;
  assign n1881 = n1111 & n1731 ;
  assign n1882 = n316 & n1699 ;
  assign n1883 = ~n1881 & ~n1882 ;
  assign n1887 = n1886 ^ n1883 ;
  assign n1888 = n1887 ^ n1883 ;
  assign n1884 = n1883 ^ n384 ;
  assign n1885 = n1884 ^ n1883 ;
  assign n1889 = n1888 ^ n1885 ;
  assign n1890 = n1883 ^ x11 ;
  assign n1891 = n1890 ^ n1883 ;
  assign n1892 = n1891 ^ n1888 ;
  assign n1893 = n1888 & ~n1892 ;
  assign n1894 = n1893 ^ n1888 ;
  assign n1895 = n1889 & n1894 ;
  assign n1896 = n1895 ^ n1893 ;
  assign n1897 = n1896 ^ n1883 ;
  assign n1898 = n1897 ^ n1888 ;
  assign n1899 = x1 & ~n1898 ;
  assign n1900 = n1899 ^ n1883 ;
  assign n1901 = ~n1880 & ~n1900 ;
  assign n1902 = ~x9 & ~x13 ;
  assign n1903 = n473 & n1902 ;
  assign n1904 = x5 & ~n1716 ;
  assign n1905 = n252 ^ n249 ;
  assign n1906 = x10 & n1905 ;
  assign n1907 = n1906 ^ n249 ;
  assign n1908 = n1904 & ~n1907 ;
  assign n1909 = n1903 & n1908 ;
  assign n1910 = n354 & n1909 ;
  assign n1911 = ~n1901 & ~n1910 ;
  assign n1912 = ~n1876 & n1911 ;
  assign n1913 = ~n1850 & n1912 ;
  assign n1914 = ~n1771 & n1913 ;
  assign n1915 = ~n1756 & n1914 ;
  assign n1916 = x15 & ~n1915 ;
  assign n1917 = n396 & n861 ;
  assign n1918 = n1414 & n1917 ;
  assign n1919 = n21 & n1786 ;
  assign n1920 = n1411 & n1919 ;
  assign n1921 = ~n1918 & ~n1920 ;
  assign n1922 = ~n528 & ~n1921 ;
  assign n1923 = n1294 & n1922 ;
  assign n1924 = n450 & n1823 ;
  assign n1925 = n1255 & n1924 ;
  assign n1926 = n222 & n1246 ;
  assign n1927 = n816 & n1273 ;
  assign n1928 = n1926 & n1927 ;
  assign n1929 = ~n1925 & ~n1928 ;
  assign n1930 = ~n284 & ~n1929 ;
  assign n1931 = ~x1 & n1823 ;
  assign n1932 = x0 & ~x13 ;
  assign n1933 = ~n284 & ~n1932 ;
  assign n1934 = n1931 & n1933 ;
  assign n1935 = n292 & n1125 ;
  assign n1936 = n450 & n1935 ;
  assign n1937 = ~n1934 & ~n1936 ;
  assign n1938 = n1414 & ~n1937 ;
  assign n1939 = ~n1930 & ~n1938 ;
  assign n1940 = n1405 & ~n1939 ;
  assign n1941 = n313 & n1715 ;
  assign n1942 = n21 & n1775 ;
  assign n1943 = ~n1941 & ~n1942 ;
  assign n1944 = n1294 & ~n1943 ;
  assign n1945 = x7 & n1290 ;
  assign n1946 = x4 & n284 ;
  assign n1947 = n1945 & n1946 ;
  assign n1948 = n1944 & n1947 ;
  assign n1949 = ~n1940 & ~n1948 ;
  assign n1950 = ~n1923 & n1949 ;
  assign n1951 = ~x9 & ~n1950 ;
  assign n1952 = x2 & ~x10 ;
  assign n1953 = ~x2 & x10 ;
  assign n1954 = ~n1952 & ~n1953 ;
  assign n1955 = x0 & ~n1954 ;
  assign n1956 = ~n1865 & n1955 ;
  assign n1957 = ~x9 & n1775 ;
  assign n1958 = n638 & n1294 ;
  assign n1959 = n1957 & n1958 ;
  assign n1960 = n73 & n1248 ;
  assign n1961 = n1415 & n1960 ;
  assign n1962 = x11 & n1961 ;
  assign n1963 = ~n1959 & ~n1962 ;
  assign n1964 = ~n1956 & n1963 ;
  assign n1965 = x1 & ~n1964 ;
  assign n1966 = n1699 & n1718 ;
  assign n1967 = n88 & n286 ;
  assign n1968 = ~n1966 & ~n1967 ;
  assign n1969 = ~x0 & x10 ;
  assign n1970 = ~n1747 & ~n1969 ;
  assign n1971 = n313 & ~n1970 ;
  assign n1972 = ~n1968 & n1971 ;
  assign n1973 = ~n1965 & ~n1972 ;
  assign n1974 = ~n43 & ~n1973 ;
  assign n1975 = n1366 & n1944 ;
  assign n1976 = ~n1974 & ~n1975 ;
  assign n1977 = ~n1293 & ~n1976 ;
  assign n1978 = n223 & n1765 ;
  assign n1979 = x9 & n221 ;
  assign n1980 = n1273 & n1979 ;
  assign n1981 = n1978 & n1980 ;
  assign n1982 = ~n1977 & ~n1981 ;
  assign n1983 = ~n1951 & n1982 ;
  assign n1984 = x7 ^ x6 ;
  assign n1985 = n1261 ^ n222 ;
  assign n1986 = n1261 ^ x7 ;
  assign n1987 = n1986 ^ n1261 ;
  assign n1988 = n1985 & ~n1987 ;
  assign n1989 = n1988 ^ n1261 ;
  assign n1990 = ~n1984 & n1989 ;
  assign n1991 = ~x9 & x10 ;
  assign n1992 = x11 & n1991 ;
  assign n1993 = n1247 & n1992 ;
  assign n1994 = ~x1 & ~x9 ;
  assign n1995 = n1405 & n1994 ;
  assign n1996 = n364 & n1316 ;
  assign n1997 = ~n1995 & ~n1996 ;
  assign n1998 = n1249 & ~n1997 ;
  assign n1999 = ~n1993 & ~n1998 ;
  assign n2000 = x13 & ~n1999 ;
  assign n2001 = ~x0 & n221 ;
  assign n2002 = ~n1767 & n2001 ;
  assign n2003 = n63 & n2002 ;
  assign n2004 = ~n2000 & ~n2003 ;
  assign n2005 = ~x2 & ~x9 ;
  assign n2006 = ~n286 & ~n2005 ;
  assign n2007 = ~n1699 & ~n1731 ;
  assign n2008 = n2006 & ~n2007 ;
  assign n2009 = n1969 & n2008 ;
  assign n2010 = n313 & n2009 ;
  assign n2011 = n1864 & n1969 ;
  assign n2012 = n1732 ^ x3 ;
  assign n2013 = n2012 ^ n1732 ;
  assign n2014 = n1970 ^ n1732 ;
  assign n2015 = n2013 & ~n2014 ;
  assign n2016 = n2015 ^ n1732 ;
  assign n2017 = n1699 & n2016 ;
  assign n2018 = ~n2011 & ~n2017 ;
  assign n2019 = n221 & ~n2018 ;
  assign n2020 = n1766 & n1941 ;
  assign n2021 = ~x10 & n21 ;
  assign n2022 = ~n1865 & n2021 ;
  assign n2023 = x2 & n2022 ;
  assign n2024 = ~n2020 & ~n2023 ;
  assign n2025 = ~n2019 & n2024 ;
  assign n2026 = ~n2010 & n2025 ;
  assign n2027 = n2026 ^ x15 ;
  assign n2028 = n2027 ^ n2004 ;
  assign n2029 = ~x9 & n285 ;
  assign n2030 = ~n1731 & ~n2029 ;
  assign n2031 = x3 & n1718 ;
  assign n2032 = ~n2030 & n2031 ;
  assign n2033 = x14 & ~n1865 ;
  assign n2034 = ~n1954 & n2033 ;
  assign n2035 = ~n2032 & ~n2034 ;
  assign n2036 = n816 & ~n2035 ;
  assign n2037 = ~x1 & n85 ;
  assign n2038 = x1 & x2 ;
  assign n2039 = ~x3 & n2038 ;
  assign n2040 = ~n2037 & ~n2039 ;
  assign n2045 = n2040 ^ n1699 ;
  assign n2053 = n2045 ^ n2040 ;
  assign n2041 = ~x1 & x9 ;
  assign n2042 = ~n943 & ~n2041 ;
  assign n2043 = n292 & ~n2042 ;
  assign n2044 = n2043 ^ n2040 ;
  assign n2046 = n2045 ^ n2044 ;
  assign n2047 = n2046 ^ n2045 ;
  assign n2048 = n2047 ^ n2040 ;
  assign n2049 = n2046 ^ n861 ;
  assign n2050 = n2049 ^ n2046 ;
  assign n2051 = n2050 ^ n2048 ;
  assign n2052 = n2048 & n2051 ;
  assign n2054 = n2053 ^ n2052 ;
  assign n2055 = n2054 ^ n2048 ;
  assign n2056 = n2040 ^ n1731 ;
  assign n2057 = n2052 ^ n2048 ;
  assign n2058 = n2056 & n2057 ;
  assign n2059 = n2058 ^ n2040 ;
  assign n2060 = n2055 & n2059 ;
  assign n2061 = n2060 ^ n2040 ;
  assign n2062 = n2061 ^ n1699 ;
  assign n2063 = n2062 ^ n2040 ;
  assign n2064 = ~x10 & n2063 ;
  assign n2065 = ~n2036 & ~n2064 ;
  assign n2066 = n2065 ^ x14 ;
  assign n2067 = ~x15 & n2066 ;
  assign n2068 = n2067 ^ n2065 ;
  assign n2069 = ~n2028 & n2068 ;
  assign n2070 = n2069 ^ n2067 ;
  assign n2071 = n2070 ^ n2065 ;
  assign n2072 = n2071 ^ x15 ;
  assign n2073 = n2004 & ~n2072 ;
  assign n2074 = n1990 & ~n2073 ;
  assign n2075 = ~x1 & ~x2 ;
  assign n2076 = n1728 & n2075 ;
  assign n2077 = n522 & n1597 ;
  assign n2078 = n2076 & n2077 ;
  assign n2079 = x9 & ~x11 ;
  assign n2080 = ~n1716 & n2079 ;
  assign n2081 = ~n691 & n2080 ;
  assign n2082 = n1700 & n2081 ;
  assign n2083 = ~n2078 & ~n2082 ;
  assign n2084 = x13 & ~n2083 ;
  assign n2085 = n25 & n1699 ;
  assign n2086 = x14 ^ x10 ;
  assign n2087 = n1702 ^ n210 ;
  assign n2088 = n1702 ^ x14 ;
  assign n2089 = n2088 ^ n1702 ;
  assign n2090 = n2087 & n2089 ;
  assign n2091 = n2090 ^ n1702 ;
  assign n2092 = ~n2086 & n2091 ;
  assign n2093 = n2085 & n2092 ;
  assign n2094 = n355 & n2093 ;
  assign n2095 = ~n2084 & ~n2094 ;
  assign n2096 = n1376 & ~n2095 ;
  assign n2097 = ~n2074 & ~n2096 ;
  assign n2098 = n1983 & n2097 ;
  assign n2099 = ~n1916 & n2098 ;
  assign n2100 = ~n1698 & ~n2099 ;
  assign n2101 = ~n1697 & ~n2100 ;
  assign n2102 = n1456 & n1747 ;
  assign n2103 = x13 & n1503 ;
  assign n2104 = n308 & n2103 ;
  assign n2105 = x6 & x9 ;
  assign n2106 = n308 & n2105 ;
  assign n2107 = ~x15 & n528 ;
  assign n2108 = n2106 & ~n2107 ;
  assign n2109 = ~x1 & n66 ;
  assign n2110 = x1 & ~n457 ;
  assign n2111 = ~n2109 & ~n2110 ;
  assign n2112 = x13 & ~n2111 ;
  assign n2113 = ~n267 & n2112 ;
  assign n2114 = ~n2108 & ~n2113 ;
  assign n2115 = x8 & ~n2114 ;
  assign n2116 = ~n2104 & ~n2115 ;
  assign n2117 = n586 & ~n2116 ;
  assign n2118 = ~n1267 & ~n1273 ;
  assign n2119 = x3 & x8 ;
  assign n2120 = ~n586 & n2119 ;
  assign n2121 = n2118 & n2120 ;
  assign n2122 = n364 & n2121 ;
  assign n2123 = x1 & x7 ;
  assign n2124 = x13 & n1598 ;
  assign n2125 = n2123 & n2124 ;
  assign n2126 = ~x6 & x9 ;
  assign n2127 = x6 ^ x3 ;
  assign n2128 = n2126 & n2127 ;
  assign n2129 = n2128 ^ n2127 ;
  assign n2130 = n2125 & n2129 ;
  assign n2131 = ~n2122 & ~n2130 ;
  assign n2132 = ~n2117 & n2131 ;
  assign n2135 = n2132 ^ n308 ;
  assign n2136 = n2135 ^ n2132 ;
  assign n2133 = n2132 ^ n2126 ;
  assign n2134 = n2133 ^ n2132 ;
  assign n2137 = n2136 ^ n2134 ;
  assign n2138 = x7 & ~x8 ;
  assign n2139 = n721 & n1394 ;
  assign n2140 = ~n2138 & ~n2139 ;
  assign n2141 = n2140 ^ n2132 ;
  assign n2142 = n2141 ^ n2132 ;
  assign n2143 = n2142 ^ n2136 ;
  assign n2144 = n2136 & ~n2143 ;
  assign n2145 = n2144 ^ n2136 ;
  assign n2146 = n2137 & n2145 ;
  assign n2147 = n2146 ^ n2144 ;
  assign n2148 = n2147 ^ n2132 ;
  assign n2149 = n2148 ^ n2136 ;
  assign n2150 = ~x2 & ~n2149 ;
  assign n2151 = n2150 ^ n2132 ;
  assign n2152 = n2102 & ~n2151 ;
  assign n2153 = ~n99 & ~n1552 ;
  assign n2154 = ~n1304 & ~n2153 ;
  assign n2155 = n1252 & n2154 ;
  assign n2156 = x8 & ~x9 ;
  assign n2157 = ~x10 & n2156 ;
  assign n2158 = n38 & n2157 ;
  assign n2159 = x11 & n2158 ;
  assign n2160 = ~n2155 & ~n2159 ;
  assign n2161 = n1990 & ~n2160 ;
  assign n2162 = x13 & ~n1352 ;
  assign n2163 = ~n373 & ~n859 ;
  assign n2164 = n2162 & ~n2163 ;
  assign n2165 = n1397 & n1903 ;
  assign n2166 = ~n2164 & ~n2165 ;
  assign n2167 = n1365 & ~n2166 ;
  assign n2168 = x9 & ~x13 ;
  assign n2169 = ~n1366 & ~n2168 ;
  assign n2170 = n99 & ~n2169 ;
  assign n2171 = ~x8 & n222 ;
  assign n2172 = n1273 & n2171 ;
  assign n2173 = n2170 & n2172 ;
  assign n2174 = ~x5 & n257 ;
  assign n2175 = n314 & n1493 ;
  assign n2176 = n2174 & n2175 ;
  assign n2177 = n1376 & n2176 ;
  assign n2178 = ~n2173 & ~n2177 ;
  assign n2179 = ~n2167 & n2178 ;
  assign n2180 = ~x10 & ~n2179 ;
  assign n2181 = x6 & ~x9 ;
  assign n2182 = ~n2126 & ~n2181 ;
  assign n2183 = n1506 & n1551 ;
  assign n2184 = n25 & n74 ;
  assign n2185 = n2183 & n2184 ;
  assign n2186 = ~x7 & ~x8 ;
  assign n2187 = n49 & n2186 ;
  assign n2188 = n1261 & n1405 ;
  assign n2189 = n2187 & n2188 ;
  assign n2190 = ~n2185 & ~n2189 ;
  assign n2191 = ~n2182 & ~n2190 ;
  assign n2192 = n1254 & n1256 ;
  assign n2193 = n721 & n2192 ;
  assign n2194 = n153 & n1273 ;
  assign n2195 = n1502 & n2194 ;
  assign n2196 = ~n2193 & ~n2195 ;
  assign n2197 = ~n1581 & ~n1619 ;
  assign n2198 = n1404 ^ x9 ;
  assign n2199 = n1404 ^ x11 ;
  assign n2200 = n2199 ^ n1404 ;
  assign n2201 = ~n2198 & n2200 ;
  assign n2202 = n2201 ^ n1404 ;
  assign n2203 = ~n2197 & n2202 ;
  assign n2204 = ~n2196 & n2203 ;
  assign n2205 = ~n2191 & ~n2204 ;
  assign n2206 = ~x4 & ~n1322 ;
  assign n2207 = ~n395 & ~n2206 ;
  assign n2208 = ~x7 & x10 ;
  assign n2209 = n118 & n2208 ;
  assign n2210 = ~n2207 & n2209 ;
  assign n2211 = n1608 & n2210 ;
  assign n2212 = n2205 & ~n2211 ;
  assign n2213 = ~n2180 & n2212 ;
  assign n2214 = ~n2161 & n2213 ;
  assign n2215 = ~n470 & ~n1251 ;
  assign n2216 = ~n2214 & n2215 ;
  assign n2217 = ~n2152 & ~n2216 ;
  assign n2218 = ~n1492 & ~n1583 ;
  assign n2219 = x9 & n2218 ;
  assign n2220 = x7 & ~n1518 ;
  assign n2221 = n1919 & n2220 ;
  assign n2222 = n2219 & n2221 ;
  assign n2223 = x3 & x6 ;
  assign n2224 = n17 & n2223 ;
  assign n2225 = x8 & ~x10 ;
  assign n2226 = ~x3 & n2225 ;
  assign n2227 = n403 & n1138 ;
  assign n2228 = ~n1492 & ~n2227 ;
  assign n2229 = n2226 & ~n2228 ;
  assign n2230 = ~n129 & ~n2229 ;
  assign n2231 = ~n2224 & n2230 ;
  assign n2232 = n1814 & ~n2231 ;
  assign n2233 = ~x13 & ~x15 ;
  assign n2234 = ~x14 & n2233 ;
  assign n2235 = n608 & n2234 ;
  assign n2236 = n149 & n1953 ;
  assign n2237 = ~n2118 & n2236 ;
  assign n2238 = ~n2235 & n2237 ;
  assign n2239 = x6 & n1952 ;
  assign n2240 = ~x3 & x6 ;
  assign n2241 = ~n1823 & ~n2240 ;
  assign n2242 = ~n2239 & ~n2241 ;
  assign n2243 = x5 & ~n1051 ;
  assign n2244 = ~n2242 & n2243 ;
  assign n2245 = ~n2238 & ~n2244 ;
  assign n2246 = ~x8 & ~n2245 ;
  assign n2247 = ~x2 & n2225 ;
  assign n2248 = n129 & n2247 ;
  assign n2249 = n1312 & n2248 ;
  assign n2250 = ~n2246 & ~n2249 ;
  assign n2251 = ~n2232 & n2250 ;
  assign n2252 = n21 & ~n2251 ;
  assign n2253 = ~x1 & n1786 ;
  assign n2254 = n1671 & n2253 ;
  assign n2255 = n25 & n2254 ;
  assign n2256 = x0 & x8 ;
  assign n2257 = x2 & x6 ;
  assign n2258 = ~x10 & n49 ;
  assign n2259 = n217 & n354 ;
  assign n2260 = n2258 & n2259 ;
  assign n2261 = n2257 & n2260 ;
  assign n2262 = n2256 & n2261 ;
  assign n2263 = ~n2255 & ~n2262 ;
  assign n2264 = n194 & ~n470 ;
  assign n2265 = ~n434 & ~n2264 ;
  assign n2266 = n1276 & ~n2265 ;
  assign n2267 = ~x5 & ~n135 ;
  assign n2268 = n38 & n2118 ;
  assign n2269 = ~n2267 & n2268 ;
  assign n2270 = ~n2266 & ~n2269 ;
  assign n2271 = ~x0 & n1953 ;
  assign n2272 = ~x3 & ~x8 ;
  assign n2273 = n2271 & n2272 ;
  assign n2274 = ~x1 & n2273 ;
  assign n2275 = ~n2270 & n2274 ;
  assign n2276 = ~x2 & x8 ;
  assign n2277 = x2 & ~x8 ;
  assign n2278 = ~n2276 & ~n2277 ;
  assign n2279 = ~x7 & ~n2278 ;
  assign n2280 = x1 & n2223 ;
  assign n2281 = ~x5 & ~n17 ;
  assign n2282 = x2 & x8 ;
  assign n2283 = ~n1719 & ~n2282 ;
  assign n2284 = n2281 & n2283 ;
  assign n2285 = n2280 & ~n2284 ;
  assign n2286 = ~n2279 & n2285 ;
  assign n2287 = x3 & n25 ;
  assign n2288 = ~n2286 & ~n2287 ;
  assign n2289 = ~n1503 & ~n1642 ;
  assign n2290 = n1718 & ~n2289 ;
  assign n2291 = ~x1 & ~n2290 ;
  assign n2292 = ~n22 & ~n2208 ;
  assign n2293 = ~n2291 & n2292 ;
  assign n2294 = ~n2288 & n2293 ;
  assign n2295 = x0 & n2294 ;
  assign n2296 = ~n2275 & ~n2295 ;
  assign n2297 = n2263 & n2296 ;
  assign n2298 = ~n2252 & n2297 ;
  assign n2299 = x9 & ~n2298 ;
  assign n2300 = n1276 & n2001 ;
  assign n2301 = n129 & n2300 ;
  assign n2302 = ~x3 & ~x6 ;
  assign n2303 = ~n2186 & ~n2302 ;
  assign n2304 = x7 & x8 ;
  assign n2305 = ~n2223 & ~n2304 ;
  assign n2306 = n165 & ~n2305 ;
  assign n2307 = ~n2303 & n2306 ;
  assign n2308 = ~x7 & n1254 ;
  assign n2309 = ~x8 & ~x14 ;
  assign n2310 = n50 & ~n2309 ;
  assign n2311 = n2308 & n2310 ;
  assign n2312 = ~n2307 & ~n2311 ;
  assign n2313 = x1 & ~n2312 ;
  assign n2314 = n117 & n1492 ;
  assign n2315 = n189 & n2314 ;
  assign n2316 = ~n2309 & n2315 ;
  assign n2317 = ~n2313 & ~n2316 ;
  assign n2318 = n1435 & ~n2317 ;
  assign n2319 = n149 & n450 ;
  assign n2320 = ~x10 & n1394 ;
  assign n2321 = n1273 & n2320 ;
  assign n2322 = n2319 & n2321 ;
  assign n2323 = ~n2318 & ~n2322 ;
  assign n2324 = ~x2 & ~n2323 ;
  assign n2325 = n2038 & n2119 ;
  assign n2326 = n129 & n2038 ;
  assign n2327 = ~n2325 & ~n2326 ;
  assign n2328 = ~x6 & ~n1630 ;
  assign n2329 = ~n1188 & ~n2328 ;
  assign n2331 = ~x10 & x12 ;
  assign n2330 = ~x12 & n1562 ;
  assign n2332 = n2331 ^ n2330 ;
  assign n2333 = n429 & n2332 ;
  assign n2334 = n2333 ^ n2331 ;
  assign n2335 = n2329 & n2334 ;
  assign n2336 = ~n2327 & n2335 ;
  assign n2337 = ~n2324 & ~n2336 ;
  assign n2338 = n1366 & ~n2337 ;
  assign n2339 = n1669 & n1702 ;
  assign n2340 = n49 & n1760 ;
  assign n2341 = n2339 & n2340 ;
  assign n2342 = x5 & x9 ;
  assign n2343 = n2271 ^ n1703 ;
  assign n2344 = n2289 ^ n2271 ;
  assign n2345 = n2344 ^ n2271 ;
  assign n2346 = n2343 & n2345 ;
  assign n2347 = n2346 ^ n2271 ;
  assign n2348 = n2342 & n2347 ;
  assign n2349 = ~n2341 & ~n2348 ;
  assign n2350 = x7 & ~n2349 ;
  assign n2351 = x0 & x6 ;
  assign n2352 = x2 & n2351 ;
  assign n2353 = n2258 & n2352 ;
  assign n2354 = ~x6 & n2271 ;
  assign n2355 = ~n2353 & ~n2354 ;
  assign n2356 = n153 & n470 ;
  assign n2357 = n551 & ~n2356 ;
  assign n2358 = n2138 & n2357 ;
  assign n2359 = ~n2355 & n2358 ;
  assign n2360 = n1394 & n2351 ;
  assign n2361 = n1952 & n2360 ;
  assign n2362 = ~x8 & n210 ;
  assign n2363 = ~n269 & n1435 ;
  assign n2364 = n2362 & n2363 ;
  assign n2365 = ~n2361 & ~n2364 ;
  assign n2366 = n2365 ^ x10 ;
  assign n2367 = n2366 ^ n2365 ;
  assign n2368 = n210 & n1642 ;
  assign n2369 = ~x12 & n33 ;
  assign n2370 = n2368 & n2369 ;
  assign n2371 = n2370 ^ n2365 ;
  assign n2372 = n2371 ^ n2365 ;
  assign n2373 = n2367 & n2372 ;
  assign n2374 = n2373 ^ n2365 ;
  assign n2375 = ~x9 & ~n2374 ;
  assign n2376 = n2375 ^ n2365 ;
  assign n2377 = n1886 & ~n2376 ;
  assign n2378 = ~n2359 & ~n2377 ;
  assign n2379 = ~n2350 & n2378 ;
  assign n2380 = ~n558 & ~n2379 ;
  assign n2381 = ~n2338 & ~n2380 ;
  assign n2382 = ~n2301 & n2381 ;
  assign n2383 = ~n2299 & n2382 ;
  assign n2384 = n2383 ^ x4 ;
  assign n2385 = n2384 ^ n2383 ;
  assign n2386 = ~x7 & x8 ;
  assign n2387 = ~x2 & x13 ;
  assign n2388 = ~x9 & n1435 ;
  assign n2389 = n2387 & n2388 ;
  assign n2390 = n2386 & n2389 ;
  assign n2391 = ~x7 & n2282 ;
  assign n2392 = ~n1758 & ~n2340 ;
  assign n2393 = n2391 & ~n2392 ;
  assign n2394 = ~n1020 & ~n2393 ;
  assign n2395 = ~n2390 & n2394 ;
  assign n2396 = ~x6 & ~n2395 ;
  assign n2397 = ~x2 & ~x8 ;
  assign n2398 = ~x7 & n2397 ;
  assign n2399 = n1260 & n1366 ;
  assign n2400 = ~n2126 & ~n2399 ;
  assign n2401 = n2398 & ~n2400 ;
  assign n2402 = x10 & n2401 ;
  assign n2403 = ~n2396 & ~n2402 ;
  assign n2404 = n308 & ~n2403 ;
  assign n2415 = x1 & ~x8 ;
  assign n2416 = n2257 & n2415 ;
  assign n2417 = n1669 & ~n1718 ;
  assign n2418 = ~n221 & n2417 ;
  assign n2419 = ~n2416 & ~n2418 ;
  assign n2420 = n1020 & ~n2419 ;
  assign n2421 = n1779 & n2075 ;
  assign n2422 = ~x6 & n1252 ;
  assign n2423 = n2421 & n2422 ;
  assign n2424 = ~x1 & x6 ;
  assign n2425 = n2391 & n2424 ;
  assign n2426 = n2340 & n2425 ;
  assign n2427 = ~n2423 & ~n2426 ;
  assign n2428 = ~n2420 & n2427 ;
  assign n2405 = ~n2282 & ~n2397 ;
  assign n2406 = n1273 & n2340 ;
  assign n2407 = n2405 & n2406 ;
  assign n2408 = n1020 & ~n1954 ;
  assign n2409 = n2289 & n2408 ;
  assign n2410 = ~x6 & ~x10 ;
  assign n2411 = n286 & n2410 ;
  assign n2412 = n2139 & n2411 ;
  assign n2413 = ~n2409 & ~n2412 ;
  assign n2414 = ~n2407 & n2413 ;
  assign n2429 = n2428 ^ n2414 ;
  assign n2430 = n2429 ^ n2428 ;
  assign n2431 = n2428 ^ x1 ;
  assign n2432 = n2431 ^ n2428 ;
  assign n2433 = ~n2430 & n2432 ;
  assign n2434 = n2433 ^ n2428 ;
  assign n2435 = ~x3 & ~n2434 ;
  assign n2436 = n2435 ^ n2428 ;
  assign n2437 = ~n2404 & n2436 ;
  assign n2438 = n104 & ~n2437 ;
  assign n2439 = n528 & n598 ;
  assign n2440 = n1669 & ~n2439 ;
  assign n2441 = n264 & n2440 ;
  assign n2442 = ~x6 & n2156 ;
  assign n2443 = n49 & n2442 ;
  assign n2444 = ~n49 & ~n1404 ;
  assign n2445 = ~x8 & ~x9 ;
  assign n2446 = ~n1404 & ~n2445 ;
  assign n2447 = ~n2444 & ~n2446 ;
  assign n2448 = n1276 & n2447 ;
  assign n2449 = ~n2443 & ~n2448 ;
  assign n2450 = ~n2441 & n2449 ;
  assign n2451 = n313 & ~n2450 ;
  assign n2452 = ~n1276 & ~n1312 ;
  assign n2453 = n460 & ~n2452 ;
  assign n2454 = x6 & n1020 ;
  assign n2455 = ~n2453 & ~n2454 ;
  assign n2456 = x1 & n2272 ;
  assign n2457 = ~n2455 & n2456 ;
  assign n2458 = ~x3 & x8 ;
  assign n2459 = n1273 ^ n49 ;
  assign n2460 = n1273 ^ n1267 ;
  assign n2461 = n2460 ^ n1267 ;
  assign n2462 = x12 & n476 ;
  assign n2463 = n2462 ^ n1267 ;
  assign n2464 = n2461 & n2463 ;
  assign n2465 = n2464 ^ n1267 ;
  assign n2466 = n2459 & ~n2465 ;
  assign n2467 = n2466 ^ n49 ;
  assign n2468 = ~n2042 & n2467 ;
  assign n2469 = x13 & n403 ;
  assign n2470 = n397 & n1994 ;
  assign n2471 = n2469 & n2470 ;
  assign n2472 = x7 & n364 ;
  assign n2473 = ~x6 & n2472 ;
  assign n2474 = ~n2471 & ~n2473 ;
  assign n2475 = ~n2468 & n2474 ;
  assign n2476 = n2458 & ~n2475 ;
  assign n2477 = ~n2457 & ~n2476 ;
  assign n2478 = ~n2451 & n2477 ;
  assign n2479 = n1952 & ~n2478 ;
  assign n2480 = n1020 & ~n2424 ;
  assign n2481 = n460 & ~n2123 ;
  assign n2482 = ~n2480 & ~n2481 ;
  assign n2483 = ~x6 & ~x9 ;
  assign n2484 = n18 & ~n2483 ;
  assign n2485 = ~x1 & ~n2484 ;
  assign n2486 = ~n2208 & ~n2272 ;
  assign n2487 = ~x2 & n2486 ;
  assign n2488 = n2303 & n2487 ;
  assign n2489 = ~n2485 & n2488 ;
  assign n2490 = ~n2482 & n2489 ;
  assign n2491 = n257 & n1283 ;
  assign n2492 = n308 & n2491 ;
  assign n2493 = ~n121 & ~n522 ;
  assign n2494 = n2424 & ~n2493 ;
  assign n2495 = n457 & n2494 ;
  assign n2496 = ~x10 & n2495 ;
  assign n2497 = ~n2492 & ~n2496 ;
  assign n2498 = ~n2278 & ~n2497 ;
  assign n2499 = ~n2490 & ~n2498 ;
  assign n2500 = x9 & n2304 ;
  assign n2501 = ~x1 & n2223 ;
  assign n2502 = n2500 & n2501 ;
  assign n2503 = ~x6 & n1404 ;
  assign n2504 = n308 & n2503 ;
  assign n2505 = ~x8 & n66 ;
  assign n2506 = x9 & n1669 ;
  assign n2507 = ~n2223 & ~n2506 ;
  assign n2508 = ~n2505 & n2507 ;
  assign n2509 = n2123 & ~n2508 ;
  assign n2510 = ~n2504 & ~n2509 ;
  assign n2511 = ~n2502 & n2510 ;
  assign n2512 = x2 & ~n2511 ;
  assign n2513 = n2499 & ~n2512 ;
  assign n2514 = ~n2479 & n2513 ;
  assign n2515 = n165 & ~n2514 ;
  assign n2516 = n692 & n1254 ;
  assign n2517 = n1952 & ~n2140 ;
  assign n2518 = n1718 & n2304 ;
  assign n2519 = ~n2517 & ~n2518 ;
  assign n2520 = n308 & ~n2519 ;
  assign n2521 = n1779 & n2272 ;
  assign n2522 = n532 & n2387 ;
  assign n2523 = n2521 & n2522 ;
  assign n2524 = ~n2520 & ~n2523 ;
  assign n2525 = n2516 & ~n2524 ;
  assign n2526 = ~n2515 & ~n2525 ;
  assign n2527 = ~n2438 & n2526 ;
  assign n2528 = n2527 ^ n2383 ;
  assign n2529 = n2385 & n2528 ;
  assign n2530 = n2529 ^ n2383 ;
  assign n2531 = ~n2222 & n2530 ;
  assign n2532 = n2217 & n2531 ;
  assign n2533 = n2101 & n2532 ;
  assign n2534 = ~n1245 & n2533 ;
  assign n2598 = x2 & ~x6 ;
  assign n2599 = n250 & n2598 ;
  assign n2600 = x2 & ~n1352 ;
  assign n2601 = ~x2 & n252 ;
  assign n2602 = ~n2600 & ~n2601 ;
  assign n2603 = ~x14 & ~n2602 ;
  assign n2604 = ~n2599 & ~n2603 ;
  assign n2605 = ~x8 & ~n2604 ;
  assign n2606 = ~x6 & n247 ;
  assign n2607 = n1667 & n2606 ;
  assign n2608 = ~n2605 & ~n2607 ;
  assign n2609 = n384 & ~n2608 ;
  assign n2558 = x8 & x14 ;
  assign n2610 = n249 & n2558 ;
  assign n2535 = ~n252 & ~n267 ;
  assign n2536 = ~n1433 & n2535 ;
  assign n2611 = ~x8 & ~n2536 ;
  assign n2612 = ~n2610 & ~n2611 ;
  assign n2613 = x2 & n66 ;
  assign n2614 = ~n2612 & n2613 ;
  assign n2537 = n2536 ^ x14 ;
  assign n2538 = n2537 ^ n2536 ;
  assign n2539 = n2536 ^ n249 ;
  assign n2540 = n2539 ^ n2536 ;
  assign n2541 = n2538 & n2540 ;
  assign n2542 = n2541 ^ n2536 ;
  assign n2543 = ~x9 & ~n2542 ;
  assign n2544 = n2543 ^ n2536 ;
  assign n2615 = ~x2 & n2119 ;
  assign n2616 = ~n2544 & n2615 ;
  assign n2586 = ~x2 & ~x14 ;
  assign n2617 = n41 & n2181 ;
  assign n2618 = n2586 & n2617 ;
  assign n2619 = ~x8 & n2618 ;
  assign n2620 = ~n2616 & ~n2619 ;
  assign n2621 = ~n2614 & n2620 ;
  assign n2622 = ~n2609 & n2621 ;
  assign n2545 = n1248 & ~n2544 ;
  assign n2546 = n249 & n1702 ;
  assign n2547 = n674 & n2546 ;
  assign n2548 = ~x2 & x9 ;
  assign n2549 = ~x0 & x14 ;
  assign n2550 = n252 & n2549 ;
  assign n2551 = n2548 & n2550 ;
  assign n2552 = ~n2547 & ~n2551 ;
  assign n2553 = ~n2545 & n2552 ;
  assign n2554 = n2458 & ~n2553 ;
  assign n2555 = x0 & ~x6 ;
  assign n2556 = n2282 & n2555 ;
  assign n2557 = n250 & n2556 ;
  assign n2559 = ~n252 & ~n2558 ;
  assign n2560 = ~n249 & ~n2309 ;
  assign n2561 = ~n1716 & n2560 ;
  assign n2562 = ~n2559 & n2561 ;
  assign n2563 = ~n2557 & ~n2562 ;
  assign n2564 = n73 & ~n2563 ;
  assign n2565 = ~x9 & ~x14 ;
  assign n2566 = n249 & n1715 ;
  assign n2567 = n278 & n2257 ;
  assign n2568 = ~n2566 & ~n2567 ;
  assign n2569 = n2565 & ~n2568 ;
  assign n2570 = x14 & n252 ;
  assign n2571 = n2570 ^ n2536 ;
  assign n2572 = n2536 ^ x2 ;
  assign n2573 = n2572 ^ n2536 ;
  assign n2574 = n2573 ^ n357 ;
  assign n2575 = ~n2571 & ~n2574 ;
  assign n2576 = n2575 ^ n2570 ;
  assign n2577 = n357 & n2576 ;
  assign n2578 = ~n2569 & ~n2577 ;
  assign n2579 = n2272 & ~n2578 ;
  assign n2580 = ~n2564 & ~n2579 ;
  assign n2581 = ~n2554 & n2580 ;
  assign n2623 = n2622 ^ n2581 ;
  assign n2582 = ~x4 & n1823 ;
  assign n2583 = n269 & n2582 ;
  assign n2584 = n2445 & n2583 ;
  assign n2585 = x9 & n252 ;
  assign n2587 = ~x3 & x14 ;
  assign n2588 = ~n832 & ~n2587 ;
  assign n2589 = n2405 & n2588 ;
  assign n2590 = ~n2586 & n2589 ;
  assign n2591 = n2585 & n2590 ;
  assign n2592 = ~x3 & n2586 ;
  assign n2593 = n249 & n1404 ;
  assign n2594 = n2592 & n2593 ;
  assign n2595 = ~n2591 & ~n2594 ;
  assign n2596 = ~n2584 & n2595 ;
  assign n2597 = n2596 ^ n2581 ;
  assign n2624 = n2623 ^ n2597 ;
  assign n2625 = n2597 ^ x0 ;
  assign n2626 = n2625 ^ n2597 ;
  assign n2627 = n2624 & n2626 ;
  assign n2628 = n2627 ^ n2597 ;
  assign n2629 = ~x1 & n2628 ;
  assign n2630 = n2629 ^ n2581 ;
  assign n2631 = x15 & ~n2630 ;
  assign n2632 = ~x2 & n450 ;
  assign n2633 = n2272 & n2585 ;
  assign n2634 = n2632 & n2633 ;
  assign n2635 = n798 & n2442 ;
  assign n2636 = n1503 & ~n2042 ;
  assign n2637 = n278 & n2636 ;
  assign n2638 = ~n2635 & ~n2637 ;
  assign n2639 = n21 & n2156 ;
  assign n2640 = ~x1 & ~x8 ;
  assign n2641 = n357 & n2640 ;
  assign n2642 = ~n2639 & ~n2641 ;
  assign n2643 = ~n1352 & ~n2642 ;
  assign n2644 = n2638 & ~n2643 ;
  assign n2645 = n1823 & ~n2644 ;
  assign n2646 = x1 & ~n1674 ;
  assign n2647 = ~x6 & n799 ;
  assign n2648 = x8 & n2647 ;
  assign n2649 = ~n2646 & ~n2648 ;
  assign n2650 = ~x2 & n101 ;
  assign n2651 = ~n2649 & n2650 ;
  assign n2652 = n2651 ^ x3 ;
  assign n2653 = n2652 ^ n2651 ;
  assign n2654 = n2653 ^ n2645 ;
  assign n2655 = ~x8 & n357 ;
  assign n2656 = x1 & ~n1352 ;
  assign n2657 = ~n2647 & ~n2656 ;
  assign n2658 = n2655 & ~n2657 ;
  assign n2659 = ~x0 & n2156 ;
  assign n2660 = x1 & ~x4 ;
  assign n2661 = ~x6 & n2660 ;
  assign n2662 = n2659 & n2661 ;
  assign n2663 = ~n2658 & ~n2662 ;
  assign n2664 = n2663 ^ x2 ;
  assign n2665 = x2 & ~n2664 ;
  assign n2666 = n2665 ^ n2651 ;
  assign n2667 = n2666 ^ x2 ;
  assign n2668 = n2654 & n2667 ;
  assign n2669 = n2668 ^ n2665 ;
  assign n2670 = n2669 ^ x2 ;
  assign n2671 = ~n2645 & n2670 ;
  assign n2672 = n2671 ^ n2645 ;
  assign n2673 = ~n2634 & ~n2672 ;
  assign n2674 = ~x14 & ~n2673 ;
  assign n2675 = ~n2631 & ~n2674 ;
  assign n2676 = n2154 & ~n2675 ;
  assign n2677 = ~n1256 & ~n1551 ;
  assign n2704 = ~x0 & x8 ;
  assign n2705 = x9 & n2704 ;
  assign n2706 = n817 & n2705 ;
  assign n2707 = ~x8 & n1366 ;
  assign n2708 = ~n2168 & ~n2707 ;
  assign n2709 = x0 & ~x8 ;
  assign n2710 = ~n2704 & ~n2709 ;
  assign n2711 = x1 & ~n2710 ;
  assign n2712 = ~n2708 & n2711 ;
  assign n2713 = ~n2706 & ~n2712 ;
  assign n2714 = n1823 & ~n2713 ;
  assign n2715 = n1493 & n1715 ;
  assign n2716 = n365 & n2715 ;
  assign n2717 = n829 & n2632 ;
  assign n2718 = n1404 & n2717 ;
  assign n2719 = ~n2716 & ~n2718 ;
  assign n2720 = ~n2714 & n2719 ;
  assign n2721 = n249 & ~n2720 ;
  assign n2678 = x3 & ~x8 ;
  assign n2679 = ~x9 & n2678 ;
  assign n2680 = ~x2 & n1404 ;
  assign n2681 = ~n2679 & ~n2680 ;
  assign n2682 = ~n1786 & ~n2681 ;
  assign n2683 = ~n1085 & n2555 ;
  assign n2684 = n425 & n816 ;
  assign n2685 = ~n2683 & ~n2684 ;
  assign n2686 = ~x4 & ~n2685 ;
  assign n2687 = ~x0 & n394 ;
  assign n2688 = n817 & n2687 ;
  assign n2689 = ~n2686 & ~n2688 ;
  assign n2690 = n2682 & ~n2689 ;
  assign n2691 = ~n228 & ~n266 ;
  assign n2692 = ~n1672 & ~n2691 ;
  assign n2693 = n61 & ~n2692 ;
  assign n2694 = ~n266 & ~n1671 ;
  assign n2695 = ~x9 & n550 ;
  assign n2696 = ~n2694 & n2695 ;
  assign n2697 = n2693 & n2696 ;
  assign n2698 = ~x0 & n550 ;
  assign n2699 = n1550 & n2181 ;
  assign n2700 = n207 & n2699 ;
  assign n2701 = n2698 & n2700 ;
  assign n2702 = ~n2697 & ~n2701 ;
  assign n2703 = ~n2690 & n2702 ;
  assign n2722 = n2721 ^ n2703 ;
  assign n2723 = n2722 ^ n2721 ;
  assign n2724 = n207 & n1503 ;
  assign n2725 = n1581 & n2598 ;
  assign n2726 = ~n2724 & ~n2725 ;
  assign n2727 = x13 & ~n2726 ;
  assign n2728 = ~n457 & n2727 ;
  assign n2729 = n1642 & n2168 ;
  assign n2730 = n2582 & n2729 ;
  assign n2731 = ~n2728 & ~n2730 ;
  assign n2732 = n816 & ~n2731 ;
  assign n2733 = n2732 ^ n2721 ;
  assign n2734 = n2733 ^ n2721 ;
  assign n2735 = n2723 & ~n2734 ;
  assign n2736 = n2735 ^ n2721 ;
  assign n2737 = x11 & ~n2736 ;
  assign n2738 = n2737 ^ n2721 ;
  assign n2739 = ~x8 & x14 ;
  assign n2740 = x4 & ~n2739 ;
  assign n2741 = n1352 & ~n2740 ;
  assign n2742 = n1702 & n2741 ;
  assign n2743 = ~n2309 & ~n2558 ;
  assign n2744 = ~n2568 & ~n2743 ;
  assign n2745 = n266 & n1642 ;
  assign n2746 = n77 & n2745 ;
  assign n2747 = ~n2744 & ~n2746 ;
  assign n2748 = ~n2742 & n2747 ;
  assign n2749 = ~n2724 & n2748 ;
  assign n2750 = n74 & ~n2749 ;
  assign n2751 = n384 & n2750 ;
  assign n2752 = ~x8 & n266 ;
  assign n2753 = ~n306 & ~n2752 ;
  assign n2754 = ~n1716 & ~n2753 ;
  assign n2755 = ~n1503 & n2754 ;
  assign n2756 = n507 & n909 ;
  assign n2757 = n2755 & n2756 ;
  assign n2758 = ~x0 & n252 ;
  assign n2759 = x8 & ~n2586 ;
  assign n2760 = n2758 & ~n2759 ;
  assign n2761 = x8 & n252 ;
  assign n2762 = ~n1826 & ~n2761 ;
  assign n2763 = ~n1667 & ~n1716 ;
  assign n2764 = ~n2762 & n2763 ;
  assign n2765 = ~x8 & ~n78 ;
  assign n2766 = n2606 & ~n2765 ;
  assign n2767 = ~n2764 & ~n2766 ;
  assign n2768 = ~n2760 & n2767 ;
  assign n2769 = n75 & ~n2768 ;
  assign n2770 = ~n2757 & ~n2769 ;
  assign n2771 = ~n2751 & n2770 ;
  assign n2772 = n2771 ^ x1 ;
  assign n2773 = n2772 ^ n2771 ;
  assign n2774 = n2773 ^ x15 ;
  assign n2775 = x11 & n469 ;
  assign n2776 = n252 & n2445 ;
  assign n2777 = ~n2593 & ~n2776 ;
  assign n2778 = ~x14 & ~n2593 ;
  assign n2779 = ~n2777 & ~n2778 ;
  assign n2780 = n2775 & n2779 ;
  assign n2781 = n235 & n269 ;
  assign n2782 = n74 & n1404 ;
  assign n2783 = n2781 & n2782 ;
  assign n2784 = ~n2780 & ~n2783 ;
  assign n2785 = n210 & ~n2784 ;
  assign n2786 = x3 & n74 ;
  assign n2787 = n2741 & n2786 ;
  assign n2788 = n1644 & n2775 ;
  assign n2789 = ~n2787 & ~n2788 ;
  assign n2792 = n2789 ^ x8 ;
  assign n2793 = n2792 ^ n2789 ;
  assign n2790 = n2789 ^ n1078 ;
  assign n2791 = n2790 ^ n2789 ;
  assign n2794 = n2793 ^ n2791 ;
  assign n2795 = n909 & n2302 ;
  assign n2796 = n2795 ^ n2789 ;
  assign n2797 = n2796 ^ n2789 ;
  assign n2798 = n2797 ^ n2793 ;
  assign n2799 = n2793 & n2798 ;
  assign n2800 = n2799 ^ n2793 ;
  assign n2801 = n2794 & n2800 ;
  assign n2802 = n2801 ^ n2799 ;
  assign n2803 = n2802 ^ n2789 ;
  assign n2804 = n2803 ^ n2793 ;
  assign n2805 = ~x9 & ~n2804 ;
  assign n2806 = n2805 ^ n2789 ;
  assign n2807 = n1702 & ~n2806 ;
  assign n2808 = ~n2785 & ~n2807 ;
  assign n2809 = ~x13 & n2079 ;
  assign n2810 = n2809 ^ n2606 ;
  assign n2811 = n2810 ^ n1644 ;
  assign n2812 = n2811 ^ n2809 ;
  assign n2813 = n2812 ^ n2811 ;
  assign n2814 = ~x14 & n74 ;
  assign n2815 = n2814 ^ n909 ;
  assign n2816 = x9 & n2815 ;
  assign n2817 = n2816 ^ n909 ;
  assign n2818 = ~x8 & n2817 ;
  assign n2819 = n2818 ^ n2811 ;
  assign n2820 = n2819 ^ n2810 ;
  assign n2821 = n2813 & ~n2820 ;
  assign n2822 = n2821 ^ n2818 ;
  assign n2823 = ~n2558 & ~n2818 ;
  assign n2824 = n2823 ^ n2810 ;
  assign n2825 = ~n2822 & ~n2824 ;
  assign n2826 = n2825 ^ n2823 ;
  assign n2827 = ~n2810 & n2826 ;
  assign n2828 = n2827 ^ n2821 ;
  assign n2829 = n2828 ^ n2606 ;
  assign n2830 = n2829 ^ n2818 ;
  assign n2831 = n50 & ~n2830 ;
  assign n2832 = ~x9 & n909 ;
  assign n2833 = n528 & n2079 ;
  assign n2834 = ~n2832 & ~n2833 ;
  assign n2835 = n2834 ^ x14 ;
  assign n2836 = n2835 ^ n2834 ;
  assign n2837 = n2834 ^ n2809 ;
  assign n2838 = n2837 ^ n2834 ;
  assign n2839 = ~n2836 & n2838 ;
  assign n2840 = n2839 ^ n2834 ;
  assign n2841 = ~x8 & ~n2840 ;
  assign n2842 = n2841 ^ n2834 ;
  assign n2843 = n218 & ~n2842 ;
  assign n2844 = n2351 & n2843 ;
  assign n2845 = ~n2831 & ~n2844 ;
  assign n2846 = n2845 ^ n2808 ;
  assign n2847 = n2808 & n2846 ;
  assign n2848 = n2847 ^ n2771 ;
  assign n2849 = n2848 ^ n2808 ;
  assign n2850 = ~n2774 & n2849 ;
  assign n2851 = n2850 ^ n2847 ;
  assign n2852 = n2851 ^ n2808 ;
  assign n2853 = x15 & n2852 ;
  assign n2854 = n2853 ^ x15 ;
  assign n2855 = ~n2738 & ~n2854 ;
  assign n2856 = ~n470 & ~n2855 ;
  assign n2857 = ~x8 & ~x13 ;
  assign n2858 = x6 & n41 ;
  assign n2859 = n2548 & n2858 ;
  assign n2860 = n2857 & n2859 ;
  assign n2861 = ~n2728 & ~n2860 ;
  assign n2862 = n24 & ~n2861 ;
  assign n2863 = n384 & n2277 ;
  assign n2864 = ~x9 & n2615 ;
  assign n2865 = ~n2863 & ~n2864 ;
  assign n2866 = ~n1085 & n2758 ;
  assign n2867 = x0 & ~n1352 ;
  assign n2868 = n817 & n2867 ;
  assign n2869 = ~n2866 & ~n2868 ;
  assign n2870 = ~n2865 & ~n2869 ;
  assign n2871 = x1 & n1366 ;
  assign n2872 = ~n228 & ~n1669 ;
  assign n2873 = n2871 & ~n2872 ;
  assign n2874 = n117 & n2873 ;
  assign n2875 = ~n2692 & n2874 ;
  assign n2876 = ~x3 & n2156 ;
  assign n2877 = ~x4 & x13 ;
  assign n2878 = n2598 & n2877 ;
  assign n2879 = n2876 & n2878 ;
  assign n2880 = n450 & n2879 ;
  assign n2881 = ~n2875 & ~n2880 ;
  assign n2882 = ~n2870 & n2881 ;
  assign n2883 = ~n2862 & n2882 ;
  assign n2884 = n2883 ^ x11 ;
  assign n2885 = n2884 ^ n2883 ;
  assign n2886 = ~x9 & n1493 ;
  assign n2887 = n2001 & n2886 ;
  assign n2888 = n21 & n1608 ;
  assign n2889 = ~n1085 & n2709 ;
  assign n2890 = ~n2888 & ~n2889 ;
  assign n2891 = n2548 & ~n2890 ;
  assign n2892 = ~n2887 & ~n2891 ;
  assign n2893 = x3 & ~n2892 ;
  assign n2894 = n234 & n1252 ;
  assign n2895 = ~n830 & n2894 ;
  assign n2896 = ~n2893 & ~n2895 ;
  assign n2897 = n252 & ~n2896 ;
  assign n2898 = n2897 ^ n2883 ;
  assign n2899 = ~n2885 & ~n2898 ;
  assign n2900 = n2899 ^ n2883 ;
  assign n2901 = ~n43 & ~n2900 ;
  assign n2902 = ~n2856 & ~n2901 ;
  assign n2903 = n2677 & ~n2902 ;
  assign n2904 = ~x9 & x15 ;
  assign n2905 = ~x9 & ~n2904 ;
  assign n2906 = x1 & ~x6 ;
  assign n2907 = n1416 & n2906 ;
  assign n2908 = n235 & n2907 ;
  assign n2909 = n1330 & n1440 ;
  assign n2910 = n538 & n2909 ;
  assign n2911 = n469 & n2910 ;
  assign n2912 = ~n2908 & ~n2911 ;
  assign n2913 = ~n1716 & ~n2912 ;
  assign n2914 = ~n1352 & ~n1943 ;
  assign n2915 = n210 & n252 ;
  assign n2916 = ~n2546 & ~n2915 ;
  assign n2917 = ~n558 & ~n2916 ;
  assign n2918 = ~n2914 & ~n2917 ;
  assign n2919 = n2154 & ~n2918 ;
  assign n2920 = ~n249 & ~n1551 ;
  assign n2921 = ~n252 & ~n1256 ;
  assign n2922 = ~n2920 & ~n2921 ;
  assign n2923 = ~n1943 & n2922 ;
  assign n2924 = ~n1253 & n2923 ;
  assign n2925 = ~n2919 & ~n2924 ;
  assign n2926 = ~n2913 & n2925 ;
  assign n2927 = n1667 & ~n2926 ;
  assign n2928 = n1256 & n1671 ;
  assign n2929 = ~x4 & n1715 ;
  assign n2930 = n2928 & n2929 ;
  assign n2931 = n1551 & n1669 ;
  assign n2932 = x4 & n2931 ;
  assign n2933 = n1248 & n2932 ;
  assign n2934 = ~n2930 & ~n2933 ;
  assign n2935 = n818 & ~n2934 ;
  assign n2936 = ~n469 & ~n2935 ;
  assign n2937 = x8 & ~x11 ;
  assign n2938 = ~x2 & n792 ;
  assign n2939 = n1551 & n2351 ;
  assign n2940 = n2938 & n2939 ;
  assign n2941 = n2937 & n2940 ;
  assign n2942 = ~x4 & n277 ;
  assign n2943 = n1599 & n2038 ;
  assign n2944 = n2942 & n2943 ;
  assign n2945 = ~x12 & n1669 ;
  assign n2946 = n207 & n538 ;
  assign n2947 = n2945 & n2946 ;
  assign n2948 = ~n2944 & ~n2947 ;
  assign n2949 = n1969 & ~n2948 ;
  assign n2950 = ~x4 & x11 ;
  assign n2951 = n24 & n2950 ;
  assign n2952 = x12 & n1952 ;
  assign n2953 = n1671 & n2952 ;
  assign n2954 = n2951 & n2953 ;
  assign n2955 = ~x3 & ~n2954 ;
  assign n2956 = ~n2949 & n2955 ;
  assign n2957 = ~n2941 & n2956 ;
  assign n2958 = ~n2936 & ~n2957 ;
  assign n2959 = n1412 & n1917 ;
  assign n2960 = n1416 & n1919 ;
  assign n2961 = ~n2959 & ~n2960 ;
  assign n2962 = ~n1674 & ~n2961 ;
  assign n2963 = ~x14 & n2962 ;
  assign n2964 = ~n2958 & ~n2963 ;
  assign n2965 = ~n2927 & n2964 ;
  assign n2966 = n2965 ^ x14 ;
  assign n2967 = n1405 & n2917 ;
  assign n2968 = x0 & ~n2602 ;
  assign n2969 = ~n2567 & ~n2968 ;
  assign n2970 = n1316 & ~n2969 ;
  assign n2971 = n308 & n2970 ;
  assign n2972 = ~n2967 & ~n2971 ;
  assign n2973 = n2857 & ~n2972 ;
  assign n2974 = n816 & n1246 ;
  assign n2975 = n252 & n2974 ;
  assign n2976 = n1405 & n2975 ;
  assign n2977 = ~x4 & ~x10 ;
  assign n2978 = ~x6 & ~x11 ;
  assign n2979 = n2977 & n2978 ;
  assign n2980 = n1924 & n2979 ;
  assign n2981 = ~n2976 & ~n2980 ;
  assign n2982 = n1608 & ~n2981 ;
  assign n2983 = n1644 & n1765 ;
  assign n2984 = x11 ^ x8 ;
  assign n2985 = n2984 ^ x13 ;
  assign n2986 = n1797 ^ x8 ;
  assign n2987 = n2986 ^ n1797 ;
  assign n2988 = ~n1285 & ~n2410 ;
  assign n2989 = n2988 ^ n1285 ;
  assign n2990 = x4 & n2989 ;
  assign n2991 = n2990 ^ n1285 ;
  assign n2992 = n2991 ^ n1797 ;
  assign n2993 = ~n2987 & n2992 ;
  assign n2994 = n2993 ^ n1797 ;
  assign n2995 = n2994 ^ n2984 ;
  assign n2996 = ~n2985 & n2995 ;
  assign n2997 = n2996 ^ n2993 ;
  assign n2998 = n2997 ^ n1797 ;
  assign n2999 = n2998 ^ x13 ;
  assign n3000 = n2984 & ~n2999 ;
  assign n3001 = n3000 ^ n2984 ;
  assign n3002 = ~n2983 & ~n3001 ;
  assign n3003 = ~n1251 & ~n3002 ;
  assign n3004 = ~n2982 & ~n3003 ;
  assign n3005 = ~n2973 & n3004 ;
  assign n3006 = n3005 ^ x12 ;
  assign n3007 = n3006 ^ n3005 ;
  assign n3008 = n1316 & n2917 ;
  assign n3009 = ~x2 & ~n1352 ;
  assign n3010 = ~n2606 & ~n3009 ;
  assign n3011 = ~x0 & ~n3010 ;
  assign n3012 = ~n2566 & ~n3011 ;
  assign n3013 = n538 & n1790 ;
  assign n3014 = ~n3012 & n3013 ;
  assign n3015 = ~n3008 & ~n3014 ;
  assign n3016 = n1550 & ~n3015 ;
  assign n3017 = n31 & n2075 ;
  assign n3018 = ~x6 & n17 ;
  assign n3019 = n1021 & n3018 ;
  assign n3020 = n3017 & n3019 ;
  assign n3021 = ~x4 & n1283 ;
  assign n3022 = n1316 & n1376 ;
  assign n3023 = ~n3021 & ~n3022 ;
  assign n3024 = ~n1251 & ~n3023 ;
  assign n3025 = ~n1253 & n3024 ;
  assign n3026 = ~x8 & n3025 ;
  assign n3027 = ~n3020 & ~n3026 ;
  assign n3028 = ~n3016 & n3027 ;
  assign n3029 = n3028 ^ n3005 ;
  assign n3030 = n3007 & n3029 ;
  assign n3031 = n3030 ^ n3005 ;
  assign n3032 = n3031 ^ n2965 ;
  assign n3033 = n2966 & ~n3032 ;
  assign n3034 = n3033 ^ n3030 ;
  assign n3035 = n3034 ^ n3005 ;
  assign n3036 = n3035 ^ x14 ;
  assign n3037 = n2965 & ~n3036 ;
  assign n3038 = n3037 ^ n2965 ;
  assign n3039 = n3038 ^ n2965 ;
  assign n3040 = ~n2905 & ~n3039 ;
  assign n3041 = ~n2903 & ~n3040 ;
  assign n3042 = ~n2676 & n3041 ;
  assign n3043 = n210 & n249 ;
  assign n3044 = n1493 & n3043 ;
  assign n3045 = n2388 & n3044 ;
  assign n3046 = n161 & n1991 ;
  assign n3047 = n1715 & n3046 ;
  assign n3048 = x2 & x12 ;
  assign n3049 = x14 & n3048 ;
  assign n3050 = n768 & n1991 ;
  assign n3051 = n3049 & n3050 ;
  assign n3052 = x9 & n1703 ;
  assign n3053 = ~n3051 & ~n3052 ;
  assign n3054 = ~n3047 & n3053 ;
  assign n3055 = n1665 & ~n3054 ;
  assign n3056 = ~x12 & n252 ;
  assign n3057 = n1562 & n1702 ;
  assign n3058 = n294 & n1760 ;
  assign n3059 = x0 & n2405 ;
  assign n3060 = ~x0 & n2282 ;
  assign n3061 = ~n3059 & ~n3060 ;
  assign n3062 = n3058 & ~n3061 ;
  assign n3063 = ~n3057 & ~n3062 ;
  assign n3064 = n3056 & ~n3063 ;
  assign n3065 = n38 & n1760 ;
  assign n3066 = ~n2320 & ~n3065 ;
  assign n3067 = n3043 & ~n3066 ;
  assign n3068 = x9 & ~x12 ;
  assign n3069 = ~x9 & x14 ;
  assign n3070 = n1256 & n3069 ;
  assign n3071 = ~n3068 & ~n3070 ;
  assign n3072 = n3044 & ~n3071 ;
  assign n3073 = ~n3067 & ~n3072 ;
  assign n3074 = ~n3064 & n3073 ;
  assign n3075 = ~n3055 & n3074 ;
  assign n3076 = x11 & ~n3075 ;
  assign n3077 = ~n3045 & ~n3076 ;
  assign n3078 = ~n558 & ~n3077 ;
  assign n3079 = n3042 & ~n3078 ;
  assign n3080 = n1294 & n2156 ;
  assign n3081 = n2280 & n3080 ;
  assign n3082 = n3081 ^ x6 ;
  assign n3083 = ~n153 & n1758 ;
  assign n3084 = n2678 & n3083 ;
  assign n3085 = ~x12 & n909 ;
  assign n3086 = n2226 & n3085 ;
  assign n3087 = ~n153 & ~n1316 ;
  assign n3088 = ~n1551 & n2505 ;
  assign n3089 = ~n3087 & n3088 ;
  assign n3090 = ~n3086 & ~n3089 ;
  assign n3091 = x14 & ~n3090 ;
  assign n3092 = ~n3084 & ~n3091 ;
  assign n3093 = n3092 ^ x1 ;
  assign n3094 = n3093 ^ n3092 ;
  assign n3095 = ~x12 & n17 ;
  assign n3096 = ~x10 & n38 ;
  assign n3097 = ~x11 & n528 ;
  assign n3098 = n17 & ~n3097 ;
  assign n3099 = ~n3096 & ~n3098 ;
  assign n3100 = ~n3095 & n3099 ;
  assign n3101 = ~n1294 & n3100 ;
  assign n3102 = n73 & ~n3101 ;
  assign n3103 = ~n314 & ~n3097 ;
  assign n3104 = ~x10 & n3103 ;
  assign n3105 = ~n1991 & ~n3104 ;
  assign n3106 = n2119 & n3105 ;
  assign n3107 = ~x10 & n62 ;
  assign n3108 = n1611 & n3107 ;
  assign n3109 = n281 & n2330 ;
  assign n3110 = ~n3108 & ~n3109 ;
  assign n3111 = n507 & ~n3110 ;
  assign n3112 = ~n3106 & ~n3111 ;
  assign n3113 = ~n3102 & n3112 ;
  assign n3114 = n3113 ^ n3092 ;
  assign n3115 = n3094 & n3114 ;
  assign n3116 = n3115 ^ n3092 ;
  assign n3117 = n3116 ^ n3081 ;
  assign n3118 = n3082 & n3117 ;
  assign n3119 = n3118 ^ n3115 ;
  assign n3120 = n3119 ^ n3092 ;
  assign n3121 = n3120 ^ x6 ;
  assign n3122 = ~n3081 & n3121 ;
  assign n3123 = n3122 ^ n3081 ;
  assign n3124 = n3123 ^ n3081 ;
  assign n3125 = n266 & ~n3124 ;
  assign n3126 = n308 & n3080 ;
  assign n3127 = n208 & n3126 ;
  assign n3128 = n17 & n1113 ;
  assign n3129 = n1252 & n1300 ;
  assign n3130 = ~n3080 & ~n3129 ;
  assign n3131 = n880 & ~n3130 ;
  assign n3132 = x13 & n3131 ;
  assign n3133 = ~n3128 & ~n3132 ;
  assign n3134 = n2858 & ~n3133 ;
  assign n3135 = ~n1404 & ~n1405 ;
  assign n3136 = ~n1316 & ~n2445 ;
  assign n3137 = x3 & ~n318 ;
  assign n3138 = n134 & n3137 ;
  assign n3139 = ~n284 & n3138 ;
  assign n3140 = n161 & n354 ;
  assign n3141 = ~n3139 & ~n3140 ;
  assign n3142 = ~n3136 & ~n3141 ;
  assign n3143 = x13 & n426 ;
  assign n3144 = n1301 & ~n2446 ;
  assign n3145 = n3143 & ~n3144 ;
  assign n3146 = ~n3142 & ~n3145 ;
  assign n3147 = ~n3135 & ~n3146 ;
  assign n3148 = n39 & n1706 ;
  assign n3149 = n2678 & n3148 ;
  assign n3150 = ~x3 & ~n34 ;
  assign n3151 = ~n3135 & n3150 ;
  assign n3152 = ~n3149 & ~n3151 ;
  assign n3153 = n880 & ~n3152 ;
  assign n3154 = ~x10 & n890 ;
  assign n3155 = n1113 & n2458 ;
  assign n3156 = n3154 & n3155 ;
  assign n3157 = ~n3153 & ~n3156 ;
  assign n3158 = x13 & ~n3157 ;
  assign n3159 = ~n369 & ~n2937 ;
  assign n3160 = ~x3 & ~n1405 ;
  assign n3161 = ~x1 & x8 ;
  assign n3162 = ~x3 & x12 ;
  assign n3163 = n3161 & ~n3162 ;
  assign n3164 = ~n3160 & ~n3163 ;
  assign n3165 = ~n314 & ~n1611 ;
  assign n3166 = x10 & ~n3165 ;
  assign n3167 = n3164 & ~n3166 ;
  assign n3168 = n3159 & n3167 ;
  assign n3169 = n3168 ^ x9 ;
  assign n3170 = n3169 ^ n3168 ;
  assign n3171 = n3170 ^ n3158 ;
  assign n3172 = x1 & ~x10 ;
  assign n3173 = ~x12 & n3172 ;
  assign n3174 = n2119 & n3173 ;
  assign n3175 = n3174 ^ x11 ;
  assign n3176 = x11 & n3175 ;
  assign n3177 = n3176 ^ n3168 ;
  assign n3178 = n3177 ^ x11 ;
  assign n3179 = n3171 & n3178 ;
  assign n3180 = n3179 ^ n3176 ;
  assign n3181 = n3180 ^ x11 ;
  assign n3182 = ~n3158 & n3181 ;
  assign n3183 = n3182 ^ n3158 ;
  assign n3184 = ~n3147 & ~n3183 ;
  assign n3185 = n2601 & ~n3184 ;
  assign n3186 = ~n3134 & ~n3185 ;
  assign n3187 = ~n3127 & n3186 ;
  assign n3188 = ~n3125 & n3187 ;
  assign n3189 = ~x0 & ~n3188 ;
  assign n3190 = n3079 & ~n3189 ;
  assign n3194 = ~x9 & n2038 ;
  assign n3195 = n3154 & n3194 ;
  assign n3196 = ~x14 & n1256 ;
  assign n3197 = ~x1 & n2548 ;
  assign n3198 = n3196 & n3197 ;
  assign n3199 = ~n3195 & ~n3198 ;
  assign n3200 = n2709 & ~n3199 ;
  assign n3201 = ~x9 & n221 ;
  assign n3202 = n3196 & n3201 ;
  assign n3203 = ~x1 & n286 ;
  assign n3204 = n3154 & n3203 ;
  assign n3205 = ~n3202 & ~n3204 ;
  assign n3206 = n2704 & ~n3205 ;
  assign n3207 = ~n3200 & ~n3206 ;
  assign n3191 = n1365 & n1748 ;
  assign n3192 = n1598 & n1749 ;
  assign n3193 = ~n3191 & ~n3192 ;
  assign n3208 = n3207 ^ n3193 ;
  assign n3209 = n3208 ^ n3207 ;
  assign n3210 = n3207 ^ n364 ;
  assign n3211 = n3210 ^ n3207 ;
  assign n3212 = ~n3209 & n3211 ;
  assign n3213 = n3212 ^ n3207 ;
  assign n3214 = ~x3 & ~n3213 ;
  assign n3215 = n3214 ^ n3207 ;
  assign n3216 = n1376 & ~n3215 ;
  assign n3217 = ~x14 & n1551 ;
  assign n3218 = n2682 & n3217 ;
  assign n3219 = n2867 & n3218 ;
  assign n3220 = ~x6 & n1073 ;
  assign n3221 = n3217 & n3220 ;
  assign n3222 = n1256 & n2570 ;
  assign n3223 = ~n3221 & ~n3222 ;
  assign n3224 = n507 & n2405 ;
  assign n3225 = ~n3223 & n3224 ;
  assign n3226 = ~x12 & n1747 ;
  assign n3227 = n247 & n1671 ;
  assign n3228 = ~x2 & n1433 ;
  assign n3229 = n1669 & n3228 ;
  assign n3230 = ~n3227 & ~n3229 ;
  assign n3231 = n3226 & ~n3230 ;
  assign n3232 = ~x0 & n1256 ;
  assign n3233 = n252 & n2276 ;
  assign n3234 = ~x14 & n1671 ;
  assign n3235 = n247 & n3234 ;
  assign n3236 = ~n3233 & ~n3235 ;
  assign n3237 = n3232 & ~n3236 ;
  assign n3238 = ~n3231 & ~n3237 ;
  assign n3239 = n73 & ~n3238 ;
  assign n3240 = ~x0 & ~n1352 ;
  assign n3241 = ~n2865 & n3240 ;
  assign n3242 = n1257 & n3241 ;
  assign n3243 = ~n3239 & ~n3242 ;
  assign n3244 = ~n3225 & n3243 ;
  assign n3245 = n228 & n1503 ;
  assign n3246 = x14 & n3245 ;
  assign n3247 = ~n2745 & ~n3246 ;
  assign n3248 = x0 & ~n3247 ;
  assign n3249 = x6 & ~x14 ;
  assign n3250 = n278 & n3249 ;
  assign n3251 = n2276 & n3250 ;
  assign n3252 = ~n3248 & ~n3251 ;
  assign n3253 = n1551 & ~n3252 ;
  assign n3254 = ~x6 & n1667 ;
  assign n3255 = n266 & n3254 ;
  assign n3256 = ~n3245 & ~n3255 ;
  assign n3257 = n3232 & ~n3256 ;
  assign n3258 = ~n3253 & ~n3257 ;
  assign n3259 = n384 & ~n3258 ;
  assign n3260 = n86 & n1248 ;
  assign n3261 = n18 & n3260 ;
  assign n3262 = n73 & n3261 ;
  assign n3263 = n655 & n1562 ;
  assign n3264 = x2 & x14 ;
  assign n3265 = n384 & n3264 ;
  assign n3266 = n3263 & n3265 ;
  assign n3267 = n17 & n62 ;
  assign n3268 = n101 & n3267 ;
  assign n3269 = ~n1799 & n3268 ;
  assign n3270 = ~n3266 & ~n3269 ;
  assign n3271 = ~n3262 & n3270 ;
  assign n3272 = ~n1376 & ~n3271 ;
  assign n3273 = ~n3259 & ~n3272 ;
  assign n3274 = n3244 & n3273 ;
  assign n3275 = ~n3219 & n3274 ;
  assign n3276 = x1 & ~n3275 ;
  assign n3277 = x3 & n78 ;
  assign n3278 = ~x0 & ~n2588 ;
  assign n3279 = ~n3277 & ~n3278 ;
  assign n3280 = n3056 & ~n3279 ;
  assign n3281 = n2680 & n3280 ;
  assign n3282 = x2 & ~x12 ;
  assign n3283 = x0 & ~x14 ;
  assign n3284 = n2446 ^ n2156 ;
  assign n3285 = x3 & ~n3284 ;
  assign n3286 = n3285 ^ n2156 ;
  assign n3287 = n249 & n3286 ;
  assign n3288 = ~n2633 & ~n3287 ;
  assign n3289 = n3283 & ~n3288 ;
  assign n3290 = ~x4 & n2289 ;
  assign n3291 = ~n1673 & ~n3290 ;
  assign n3292 = n77 & ~n3291 ;
  assign n3293 = n66 & ~n3292 ;
  assign n3296 = x0 & x4 ;
  assign n3297 = n267 & n3296 ;
  assign n3294 = ~x0 & ~x4 ;
  assign n3295 = ~x6 & n3294 ;
  assign n3298 = n3297 ^ n3295 ;
  assign n3299 = n3297 ^ x8 ;
  assign n3300 = n3299 ^ n3297 ;
  assign n3301 = n3300 ^ n3293 ;
  assign n3302 = n3301 ^ n3292 ;
  assign n3303 = n3298 & ~n3302 ;
  assign n3304 = n3303 ^ n3297 ;
  assign n3305 = n3293 & n3304 ;
  assign n3306 = n3305 ^ n3293 ;
  assign n3307 = n3306 ^ n66 ;
  assign n3308 = ~n3289 & ~n3307 ;
  assign n3309 = n3282 & ~n3308 ;
  assign n3310 = ~n3281 & ~n3309 ;
  assign n3311 = n3310 ^ x10 ;
  assign n3312 = n3311 ^ n3310 ;
  assign n3313 = n3312 ^ x1 ;
  assign n3314 = x2 & ~x14 ;
  assign n3315 = ~n252 & ~n3314 ;
  assign n3316 = ~n249 & ~n292 ;
  assign n3317 = ~n3315 & ~n3316 ;
  assign n3318 = n2709 & n3317 ;
  assign n3319 = ~x0 & n3246 ;
  assign n3320 = n1642 & n3294 ;
  assign n3321 = n292 & n3320 ;
  assign n3322 = ~n3319 & ~n3321 ;
  assign n3323 = ~n3318 & n3322 ;
  assign n3324 = n384 & ~n3323 ;
  assign n3325 = ~x0 & ~n2570 ;
  assign n3326 = n2397 & ~n2536 ;
  assign n3327 = ~n3325 & n3326 ;
  assign n3328 = n78 & n1352 ;
  assign n3329 = n269 & n3294 ;
  assign n3330 = ~n3328 & ~n3329 ;
  assign n3331 = ~n2278 & ~n3330 ;
  assign n3332 = ~n3327 & ~n3331 ;
  assign n3333 = n66 & ~n3332 ;
  assign n3334 = x8 ^ x3 ;
  assign n3335 = n3334 ^ x0 ;
  assign n3336 = n3335 ^ x8 ;
  assign n3337 = n3336 ^ x0 ;
  assign n3338 = n3337 ^ n3336 ;
  assign n3341 = n3336 ^ n2725 ;
  assign n3342 = ~n3336 & n3341 ;
  assign n3339 = n252 & ~n3335 ;
  assign n3345 = n3342 ^ n3339 ;
  assign n3340 = n3339 ^ n3338 ;
  assign n3343 = n3342 ^ n3336 ;
  assign n3344 = ~n3340 & ~n3343 ;
  assign n3346 = n3345 ^ n3344 ;
  assign n3347 = ~n3338 & n3346 ;
  assign n3348 = n3347 ^ n3342 ;
  assign n3349 = n3348 ^ n3344 ;
  assign n3350 = n3069 & n3349 ;
  assign n3351 = ~n3333 & ~n3350 ;
  assign n3352 = ~n3324 & n3351 ;
  assign n3353 = n3352 ^ x12 ;
  assign n3354 = x12 & ~n3353 ;
  assign n3355 = n3354 ^ n3310 ;
  assign n3356 = n3355 ^ x12 ;
  assign n3357 = ~n3313 & ~n3356 ;
  assign n3358 = n3357 ^ n3354 ;
  assign n3359 = n3358 ^ x12 ;
  assign n3360 = ~x1 & n3359 ;
  assign n3361 = ~n3276 & ~n3360 ;
  assign n3362 = x15 & ~n3361 ;
  assign n3366 = x9 & n2922 ;
  assign n3364 = n1702 & n2309 ;
  assign n3363 = n210 & n2558 ;
  assign n3365 = n3364 ^ n3363 ;
  assign n3367 = n3366 ^ n3365 ;
  assign n3368 = n3367 ^ n3363 ;
  assign n3374 = n3368 ^ n3365 ;
  assign n3375 = n3374 ^ n3363 ;
  assign n3376 = n3375 ^ n3363 ;
  assign n3377 = n249 & n1551 ;
  assign n3378 = n3377 ^ n3365 ;
  assign n3379 = n3378 ^ n3365 ;
  assign n3380 = n3379 ^ n3363 ;
  assign n3381 = n3376 & n3380 ;
  assign n3369 = n252 & n1256 ;
  assign n3370 = n3369 ^ n3365 ;
  assign n3371 = n3370 ^ n3368 ;
  assign n3372 = n3371 ^ n3363 ;
  assign n3373 = n3368 & n3372 ;
  assign n3382 = n3381 ^ n3373 ;
  assign n3383 = n3382 ^ n3368 ;
  assign n3384 = n3373 ^ n3363 ;
  assign n3385 = n3384 ^ n3375 ;
  assign n3386 = ~n3363 & n3385 ;
  assign n3387 = n3386 ^ n3373 ;
  assign n3388 = n3383 & n3387 ;
  assign n3389 = n3388 ^ n3381 ;
  assign n3390 = n3389 ^ n3386 ;
  assign n3391 = n3390 ^ n3368 ;
  assign n3392 = n3391 ^ n3363 ;
  assign n3393 = n3392 ^ n3375 ;
  assign n3394 = n3393 ^ n3364 ;
  assign n3395 = n355 & n3394 ;
  assign n3396 = n2606 & n3154 ;
  assign n3397 = n503 & n1285 ;
  assign n3398 = n218 & n3397 ;
  assign n3399 = ~n3396 & ~n3398 ;
  assign n3400 = x9 & n2640 ;
  assign n3401 = ~n3399 & n3400 ;
  assign n3402 = n2325 & n2565 ;
  assign n3403 = n2922 & n3402 ;
  assign n3404 = x3 & n2922 ;
  assign n3405 = ~n3377 & ~n3404 ;
  assign n3406 = x14 & n2445 ;
  assign n3407 = n2038 & n3406 ;
  assign n3408 = ~n3405 & n3407 ;
  assign n3409 = ~n3403 & ~n3408 ;
  assign n3410 = ~n3401 & n3409 ;
  assign n3411 = n3410 ^ x0 ;
  assign n3412 = n3411 ^ n3410 ;
  assign n3413 = n292 & n943 ;
  assign n3414 = n2922 & n3413 ;
  assign n3415 = n2678 & n3414 ;
  assign n3416 = ~n3369 & ~n3404 ;
  assign n3417 = n943 & n2276 ;
  assign n3418 = ~x14 & n3417 ;
  assign n3419 = ~n3416 & n3418 ;
  assign n3420 = n2601 & n3196 ;
  assign n3421 = x3 & ~x6 ;
  assign n3422 = ~x4 & n3421 ;
  assign n3423 = n1952 & n3422 ;
  assign n3424 = n890 & n3423 ;
  assign n3425 = ~n3420 & ~n3424 ;
  assign n3426 = ~x1 & n1404 ;
  assign n3427 = ~n3425 & n3426 ;
  assign n3428 = ~n3419 & ~n3427 ;
  assign n3429 = ~n3415 & n3428 ;
  assign n3430 = n3429 ^ n3410 ;
  assign n3431 = n3412 & n3430 ;
  assign n3432 = n3431 ^ n3410 ;
  assign n3433 = ~n3395 & n3432 ;
  assign n3434 = ~n3362 & n3433 ;
  assign n3435 = ~n3216 & n3434 ;
  assign n3436 = ~n1253 & ~n3435 ;
  assign n3437 = n18 & n890 ;
  assign n3438 = n2566 & n3437 ;
  assign n3439 = n17 & n503 ;
  assign n3440 = n2567 & n3439 ;
  assign n3441 = ~n3438 & ~n3440 ;
  assign n3442 = n2330 & n2978 ;
  assign n3443 = n2929 & n3442 ;
  assign n3444 = n3441 & ~n3443 ;
  assign n3445 = ~n1253 & ~n3444 ;
  assign n3446 = x1 & n252 ;
  assign n3447 = n1732 & ~n2405 ;
  assign n3448 = ~n49 & ~n86 ;
  assign n3449 = ~x11 & n3448 ;
  assign n3450 = ~n1599 & ~n3449 ;
  assign n3451 = n3447 & n3450 ;
  assign n3452 = x8 & n1702 ;
  assign n3453 = x14 & n133 ;
  assign n3454 = ~x10 & ~n3453 ;
  assign n3455 = n3452 & n3454 ;
  assign n3456 = ~n1253 & n3196 ;
  assign n3457 = ~n1294 & ~n3456 ;
  assign n3458 = n2362 & ~n3457 ;
  assign n3459 = ~n3455 & ~n3458 ;
  assign n3460 = ~n3451 & n3459 ;
  assign n3461 = n3446 & ~n3460 ;
  assign n3462 = ~n205 & ~n2555 ;
  assign n3463 = ~n49 & ~n1405 ;
  assign n3464 = ~n3087 & ~n3463 ;
  assign n3465 = ~n3462 & n3464 ;
  assign n3466 = ~n1253 & n2939 ;
  assign n3467 = ~n3465 & ~n3466 ;
  assign n3470 = n3467 ^ x6 ;
  assign n3471 = n3470 ^ n3467 ;
  assign n3468 = n3467 ^ n1256 ;
  assign n3469 = n3468 ^ n3467 ;
  assign n3472 = n3471 ^ n3469 ;
  assign n3473 = ~x0 & ~n1253 ;
  assign n3474 = x0 & n74 ;
  assign n3475 = ~n3473 & ~n3474 ;
  assign n3476 = n3475 ^ n3467 ;
  assign n3477 = n3476 ^ n3467 ;
  assign n3478 = n3477 ^ n3471 ;
  assign n3479 = n3471 & ~n3478 ;
  assign n3480 = n3479 ^ n3471 ;
  assign n3481 = n3472 & n3480 ;
  assign n3482 = n3481 ^ n3479 ;
  assign n3483 = n3482 ^ n3467 ;
  assign n3484 = n3483 ^ n3471 ;
  assign n3485 = x14 & ~n3484 ;
  assign n3486 = n3485 ^ n3467 ;
  assign n3487 = n2397 & ~n3486 ;
  assign n3488 = n2257 & n2558 ;
  assign n3489 = ~n2677 & n3473 ;
  assign n3490 = x0 & n3463 ;
  assign n3491 = ~n1551 & n3490 ;
  assign n3492 = ~n3489 & ~n3491 ;
  assign n3493 = n3488 & ~n3492 ;
  assign n3494 = ~n3487 & ~n3493 ;
  assign n3495 = n71 & ~n3494 ;
  assign n3496 = x1 & ~n3495 ;
  assign n3497 = ~x12 & n267 ;
  assign n3498 = ~n2877 & ~n3497 ;
  assign n3499 = ~n291 & ~n3498 ;
  assign n3500 = n2282 & n3499 ;
  assign n3501 = ~x6 & n503 ;
  assign n3502 = ~n119 & ~n3501 ;
  assign n3503 = ~n394 & n2397 ;
  assign n3504 = ~n3502 & n3503 ;
  assign n3505 = ~n3500 & ~n3504 ;
  assign n3506 = ~n1970 & ~n3505 ;
  assign n3507 = ~x0 & n2877 ;
  assign n3508 = ~x2 & ~x12 ;
  assign n3509 = ~x14 & n3508 ;
  assign n3510 = n3509 ^ x2 ;
  assign n3511 = n3510 ^ n3509 ;
  assign n3512 = n3509 ^ n3107 ;
  assign n3513 = n3512 ^ n3509 ;
  assign n3514 = n3511 & n3513 ;
  assign n3515 = n3514 ^ n3509 ;
  assign n3516 = x8 & n3515 ;
  assign n3517 = n3516 ^ n3509 ;
  assign n3518 = n3507 & n3517 ;
  assign n3519 = n3518 ^ n1732 ;
  assign n3520 = n3519 ^ x6 ;
  assign n3529 = n3520 ^ n3519 ;
  assign n3521 = n249 & n2586 ;
  assign n3522 = n2857 & n3521 ;
  assign n3523 = n3522 ^ n3520 ;
  assign n3524 = n3523 ^ n3519 ;
  assign n3525 = n3520 ^ n3518 ;
  assign n3526 = n3525 ^ n3522 ;
  assign n3527 = n3526 ^ n3524 ;
  assign n3528 = n3524 & ~n3527 ;
  assign n3530 = n3529 ^ n3528 ;
  assign n3531 = n3530 ^ n3524 ;
  assign n3532 = n228 & n1394 ;
  assign n3533 = n281 & n3532 ;
  assign n3534 = n3533 ^ n3519 ;
  assign n3535 = n3528 ^ n3524 ;
  assign n3536 = ~n3534 & n3535 ;
  assign n3537 = n3536 ^ n3519 ;
  assign n3538 = ~n3531 & n3537 ;
  assign n3539 = n3538 ^ n3519 ;
  assign n3540 = n3539 ^ n1732 ;
  assign n3541 = n3540 ^ n3519 ;
  assign n3542 = n369 & ~n3541 ;
  assign n3543 = ~n3506 & n3542 ;
  assign n3544 = x15 & ~n3543 ;
  assign n3545 = ~x0 & n1303 ;
  assign n3546 = ~n2558 & n3545 ;
  assign n3547 = ~n1932 & n2309 ;
  assign n3548 = ~n1747 & n3547 ;
  assign n3549 = ~n3546 & ~n3548 ;
  assign n3550 = n2942 & ~n3549 ;
  assign n3551 = ~n1797 & ~n3021 ;
  assign n3552 = ~n1309 & ~n1415 ;
  assign n3553 = n77 & n1528 ;
  assign n3554 = n3552 & n3553 ;
  assign n3555 = ~n3551 & n3554 ;
  assign n3556 = n1826 & n2857 ;
  assign n3557 = n425 & n1433 ;
  assign n3558 = n2225 & n3557 ;
  assign n3559 = ~n3556 & ~n3558 ;
  assign n3560 = n244 & ~n3559 ;
  assign n3561 = ~n3555 & ~n3560 ;
  assign n3562 = ~n3550 & n3561 ;
  assign n3563 = n3562 ^ x2 ;
  assign n3564 = n3563 ^ n3562 ;
  assign n3565 = n284 & n1551 ;
  assign n3566 = n3295 & n3565 ;
  assign n3573 = ~n58 & n528 ;
  assign n3567 = n528 & n3295 ;
  assign n3568 = ~n3297 & ~n3567 ;
  assign n3574 = n3573 ^ n3568 ;
  assign n3575 = n3574 ^ n3568 ;
  assign n3569 = x12 & ~n1732 ;
  assign n3570 = ~n1733 & n3569 ;
  assign n3571 = n3570 ^ n3568 ;
  assign n3572 = n3571 ^ n3568 ;
  assign n3576 = n3575 ^ n3572 ;
  assign n3577 = n3568 ^ n252 ;
  assign n3578 = n3577 ^ n3568 ;
  assign n3579 = n3578 ^ n3575 ;
  assign n3580 = n3575 & n3579 ;
  assign n3581 = n3580 ^ n3575 ;
  assign n3582 = ~n3576 & n3581 ;
  assign n3583 = n3582 ^ n3580 ;
  assign n3584 = n3583 ^ n3568 ;
  assign n3585 = n3584 ^ n3575 ;
  assign n3586 = ~n1435 & ~n3585 ;
  assign n3587 = n3586 ^ n3568 ;
  assign n3588 = ~n3566 & n3587 ;
  assign n3589 = x8 & ~n3588 ;
  assign n3590 = n2761 & n3154 ;
  assign n3591 = n1629 & n2309 ;
  assign n3592 = ~n3590 & ~n3591 ;
  assign n3593 = n768 & ~n3592 ;
  assign n3594 = ~n890 & ~n1602 ;
  assign n3595 = x6 & n3296 ;
  assign n3596 = n1309 & n3595 ;
  assign n3597 = ~n3594 & n3596 ;
  assign n3598 = ~n3593 & ~n3597 ;
  assign n3599 = ~n3589 & n3598 ;
  assign n3600 = n3599 ^ n3562 ;
  assign n3601 = n3564 & n3600 ;
  assign n3602 = n3601 ^ n3562 ;
  assign n3603 = n538 & n3602 ;
  assign n3604 = n3544 & ~n3603 ;
  assign n3605 = n3043 & ~n3110 ;
  assign n3606 = n561 ^ x11 ;
  assign n3607 = n3606 ^ n561 ;
  assign n3608 = n3448 ^ n561 ;
  assign n3609 = n3608 ^ n561 ;
  assign n3610 = n3607 & ~n3609 ;
  assign n3611 = n3610 ^ n561 ;
  assign n3612 = x10 & n3611 ;
  assign n3613 = n3612 ^ n561 ;
  assign n3614 = n2339 & n3613 ;
  assign n3615 = x4 & n3614 ;
  assign n3616 = ~n3605 & ~n3615 ;
  assign n3617 = ~n3604 & n3616 ;
  assign n3618 = ~n3496 & ~n3617 ;
  assign n3619 = ~n2356 & n2362 ;
  assign n3620 = ~x11 & ~n334 ;
  assign n3621 = ~x8 & ~n3085 ;
  assign n3622 = n1702 & ~n3621 ;
  assign n3623 = ~n3620 & n3622 ;
  assign n3624 = ~n3619 & ~n3623 ;
  assign n3625 = x10 & ~n3624 ;
  assign n3627 = ~n470 & n1551 ;
  assign n3628 = n2278 & n3627 ;
  assign n3629 = ~n2739 & n3628 ;
  assign n3630 = n1708 & n2397 ;
  assign n3631 = n343 & n3630 ;
  assign n3632 = ~n3629 & ~n3631 ;
  assign n3626 = n42 & n1256 ;
  assign n3633 = n3632 ^ n3626 ;
  assign n3634 = n3633 ^ n3632 ;
  assign n3635 = n3632 ^ n2282 ;
  assign n3636 = n3635 ^ n3632 ;
  assign n3637 = n3634 & n3636 ;
  assign n3638 = n3637 ^ n3632 ;
  assign n3639 = ~x0 & ~n3638 ;
  assign n3640 = n3639 ^ n3632 ;
  assign n3641 = ~n1253 & ~n3640 ;
  assign n3642 = n314 & ~n470 ;
  assign n3643 = ~x0 & ~x8 ;
  assign n3644 = n1718 & n3643 ;
  assign n3645 = n3642 & n3644 ;
  assign n3646 = ~n3641 & ~n3645 ;
  assign n3647 = ~n3625 & n3646 ;
  assign n3648 = n2661 & ~n3647 ;
  assign n3649 = ~x0 & ~x6 ;
  assign n3650 = ~n470 & n2282 ;
  assign n3651 = n3649 & n3650 ;
  assign n3652 = x0 & x15 ;
  assign n3653 = n2397 & n3652 ;
  assign n3654 = ~n267 & n3653 ;
  assign n3655 = ~n3651 & ~n3654 ;
  assign n3656 = n2660 & ~n3655 ;
  assign n3657 = n3464 & n3656 ;
  assign n3658 = ~x8 & ~n153 ;
  assign n3659 = ~n1256 & n3658 ;
  assign n3660 = n2566 & n3659 ;
  assign n3661 = n17 & ~n133 ;
  assign n3662 = n2567 & n3661 ;
  assign n3663 = ~n3660 & ~n3662 ;
  assign n3664 = x11 & ~n3663 ;
  assign n3665 = ~n3657 & ~n3664 ;
  assign n3666 = ~n3648 & n3665 ;
  assign n3667 = ~n3618 & n3666 ;
  assign n3668 = ~n3461 & n3667 ;
  assign n3669 = ~n3445 & n3668 ;
  assign n3670 = ~n457 & ~n3669 ;
  assign n3671 = ~x0 & n2548 ;
  assign n3672 = n3642 & n3671 ;
  assign n3673 = ~n86 & ~n1588 ;
  assign n3674 = n1702 & n1728 ;
  assign n3675 = ~n3673 & n3674 ;
  assign n3676 = ~n3672 & ~n3675 ;
  assign n3677 = n1309 & ~n3676 ;
  assign n3678 = ~n470 & n1415 ;
  assign n3679 = n67 & n3671 ;
  assign n3680 = n3678 & n3679 ;
  assign n3681 = ~n3677 & ~n3680 ;
  assign n3684 = n3681 ^ n1992 ;
  assign n3685 = n3684 ^ n3681 ;
  assign n3682 = n3681 ^ n162 ;
  assign n3683 = n3682 ^ n3681 ;
  assign n3686 = n3685 ^ n3683 ;
  assign n3687 = n3681 ^ n210 ;
  assign n3688 = n3687 ^ n3681 ;
  assign n3689 = n3688 ^ n3685 ;
  assign n3690 = n3685 & n3689 ;
  assign n3691 = n3690 ^ n3685 ;
  assign n3692 = ~n3686 & n3691 ;
  assign n3693 = n3692 ^ n3690 ;
  assign n3694 = n3693 ^ n3681 ;
  assign n3695 = n3694 ^ n3685 ;
  assign n3696 = ~x8 & ~n3695 ;
  assign n3697 = n3696 ^ n3681 ;
  assign n3698 = n355 & ~n3697 ;
  assign n3699 = n1376 & n3698 ;
  assign n3700 = n2254 & n2950 ;
  assign n3701 = n41 & n1669 ;
  assign n3702 = n32 & n2978 ;
  assign n3703 = n1550 & n3702 ;
  assign n3704 = ~n3701 & ~n3703 ;
  assign n3705 = n2038 & ~n3704 ;
  assign n3706 = ~n3700 & ~n3705 ;
  assign n3707 = n357 & ~n3706 ;
  assign n3708 = x3 & x10 ;
  assign n3709 = ~x11 & ~n460 ;
  assign n3710 = n792 & n1503 ;
  assign n3711 = n2006 & n3710 ;
  assign n3712 = ~n3709 & n3711 ;
  assign n3713 = n356 & n2075 ;
  assign n3714 = n2593 & n3713 ;
  assign n3715 = ~n3712 & ~n3714 ;
  assign n3716 = n3708 & ~n3715 ;
  assign n3717 = n18 & n249 ;
  assign n3718 = n29 & n2038 ;
  assign n3719 = n3717 & n3718 ;
  assign n3720 = ~n3716 & ~n3719 ;
  assign n3721 = ~n3707 & n3720 ;
  assign n3722 = ~n3699 & n3721 ;
  assign n3723 = ~n3670 & n3722 ;
  assign n3724 = ~n3436 & n3723 ;
  assign n3725 = ~n2282 & ~n3264 ;
  assign n3726 = n550 & n3725 ;
  assign n3727 = n249 & n3726 ;
  assign n3728 = ~x2 & ~x6 ;
  assign n3729 = n2309 & n3728 ;
  assign n3730 = ~n3488 & ~n3729 ;
  assign n3731 = n3730 ^ n2257 ;
  assign n3732 = n3731 ^ n3730 ;
  assign n3733 = n3730 ^ n2739 ;
  assign n3734 = n3733 ^ n3730 ;
  assign n3735 = n3732 & n3734 ;
  assign n3736 = n3735 ^ n3730 ;
  assign n3737 = x1 & ~n3736 ;
  assign n3738 = n3737 ^ n3730 ;
  assign n3739 = n41 & ~n3738 ;
  assign n3740 = ~x8 & n2038 ;
  assign n3741 = ~x1 & ~n2405 ;
  assign n3742 = ~n3740 & ~n3741 ;
  assign n3743 = x14 & ~n3742 ;
  assign n3744 = n3422 & n3743 ;
  assign n3745 = ~x14 & n1503 ;
  assign n3746 = n235 & n3745 ;
  assign n3747 = n2075 & n3746 ;
  assign n3748 = ~n3744 & ~n3747 ;
  assign n3749 = ~n3739 & n3748 ;
  assign n3750 = ~n3727 & n3749 ;
  assign n3751 = n357 & ~n3750 ;
  assign n3752 = n1823 & n2661 ;
  assign n3753 = n2445 & n3752 ;
  assign n3754 = ~n3751 & ~n3753 ;
  assign n3755 = n133 & ~n3754 ;
  assign n3756 = ~x6 & n926 ;
  assign n3757 = n1457 & n3756 ;
  assign n3758 = ~n2865 & n3757 ;
  assign n3759 = n31 & n234 ;
  assign n3760 = ~x14 & n1902 ;
  assign n3761 = n1642 & n3760 ;
  assign n3762 = n3759 & n3761 ;
  assign n3763 = n2109 & n2282 ;
  assign n3764 = n221 & n1125 ;
  assign n3765 = n2445 & n3764 ;
  assign n3766 = ~n3763 & ~n3765 ;
  assign n3767 = n3297 & ~n3766 ;
  assign n3768 = ~n3762 & ~n3767 ;
  assign n3769 = ~x12 & ~n3768 ;
  assign n3770 = n550 & n2700 ;
  assign n3771 = ~n3769 & ~n3770 ;
  assign n3772 = ~n3758 & n3771 ;
  assign n3773 = ~n655 & ~n3772 ;
  assign n3774 = n532 & n2758 ;
  assign n3775 = ~n284 & n3774 ;
  assign n3776 = n3446 & n3453 ;
  assign n3777 = n24 & n3499 ;
  assign n3778 = ~n3776 & ~n3777 ;
  assign n3779 = ~n3775 & n3778 ;
  assign n3780 = n2682 & ~n3779 ;
  assign n3781 = n2698 & n3760 ;
  assign n3782 = ~x9 & n469 ;
  assign n3783 = n450 & n3782 ;
  assign n3784 = ~n3781 & ~n3783 ;
  assign n3785 = n249 & ~n3784 ;
  assign n3786 = n861 & n1330 ;
  assign n3787 = n267 & n943 ;
  assign n3788 = n3786 & n3787 ;
  assign n3789 = n269 & n1457 ;
  assign n3790 = n655 & n2109 ;
  assign n3791 = n3789 & n3790 ;
  assign n3792 = ~n3788 & ~n3791 ;
  assign n3793 = ~n3785 & n3792 ;
  assign n3794 = n2405 & ~n3793 ;
  assign n3795 = ~n3780 & ~n3794 ;
  assign n3796 = ~x4 & n603 ;
  assign n3797 = ~x1 & n469 ;
  assign n3798 = n1671 & n3797 ;
  assign n3799 = n308 & n528 ;
  assign n3800 = ~n2289 & n3799 ;
  assign n3801 = ~n3798 & ~n3800 ;
  assign n3802 = n3796 & ~n3801 ;
  assign n3803 = x8 & ~n267 ;
  assign n3804 = ~n269 & ~n3803 ;
  assign n3805 = x1 & n41 ;
  assign n3806 = n1368 & n3805 ;
  assign n3807 = n3804 & n3806 ;
  assign n3808 = n38 & n2565 ;
  assign n3809 = ~x1 & ~x6 ;
  assign n3810 = n31 & n3809 ;
  assign n3811 = n3808 & n3810 ;
  assign n3812 = ~n3807 & ~n3811 ;
  assign n3813 = ~n3802 & n3812 ;
  assign n3814 = ~n1716 & ~n3813 ;
  assign n3815 = n3795 & ~n3814 ;
  assign n3816 = ~n3773 & n3815 ;
  assign n3817 = ~n3755 & n3816 ;
  assign n3818 = n1300 & ~n3817 ;
  assign n3819 = ~x10 & n1404 ;
  assign n3820 = n3453 & n3819 ;
  assign n3821 = x4 & n1702 ;
  assign n3822 = n2223 & n3821 ;
  assign n3823 = n3820 & n3822 ;
  assign n3824 = ~x6 & n1438 ;
  assign n3825 = x9 ^ x3 ;
  assign n3826 = n2857 ^ n1493 ;
  assign n3827 = n1493 ^ x9 ;
  assign n3828 = n3827 ^ n1493 ;
  assign n3829 = n3826 & n3828 ;
  assign n3830 = n3829 ^ n1493 ;
  assign n3831 = ~n3825 & n3830 ;
  assign n3832 = n3824 & n3831 ;
  assign n3833 = n210 & n3832 ;
  assign n3834 = n1708 & n3833 ;
  assign n3835 = ~n3823 & ~n3834 ;
  assign n3836 = ~x1 & ~n3835 ;
  assign n3837 = n2570 & n3095 ;
  assign n3844 = n249 & n1598 ;
  assign n3845 = n1530 & n3844 ;
  assign n3846 = ~n3837 & ~n3845 ;
  assign n3847 = ~n1716 & ~n3846 ;
  assign n3848 = n252 & n1702 ;
  assign n3849 = n890 & n1562 ;
  assign n3850 = n3848 & n3849 ;
  assign n3851 = n1667 & n2331 ;
  assign n3852 = n3043 & n3851 ;
  assign n3853 = ~n3850 & ~n3852 ;
  assign n3854 = ~n3847 & n3853 ;
  assign n3838 = n1702 & n3837 ;
  assign n3839 = ~x4 & n245 ;
  assign n3840 = n3728 & n3839 ;
  assign n3841 = ~x10 & n2309 ;
  assign n3842 = n3840 & n3841 ;
  assign n3843 = ~n3838 & ~n3842 ;
  assign n3855 = n3854 ^ n3843 ;
  assign n3856 = n3854 ^ x1 ;
  assign n3857 = n3856 ^ n3854 ;
  assign n3858 = n3857 ^ n507 ;
  assign n3859 = n3858 ^ x9 ;
  assign n3860 = n3855 & ~n3859 ;
  assign n3861 = n3860 ^ n3854 ;
  assign n3862 = n507 & n3861 ;
  assign n3863 = n3862 ^ n507 ;
  assign n3864 = n1733 & n3509 ;
  assign n3865 = ~x10 & n1365 ;
  assign n3866 = ~n1716 & ~n3865 ;
  assign n3867 = ~n1546 & n3866 ;
  assign n3868 = n1702 & n2558 ;
  assign n3869 = n1551 & n3868 ;
  assign n3870 = ~n3057 & ~n3869 ;
  assign n3871 = ~n3867 & n3870 ;
  assign n3872 = ~n3864 & n3871 ;
  assign n3873 = n249 & ~n3872 ;
  assign n3877 = ~n1256 & ~n1716 ;
  assign n3878 = x12 & ~n1710 ;
  assign n3879 = ~n3877 & ~n3878 ;
  assign n3880 = ~n3864 & n3879 ;
  assign n3874 = n62 & ~n1955 ;
  assign n3875 = ~n210 & ~n3874 ;
  assign n3876 = ~n1969 & ~n3875 ;
  assign n3881 = n3880 ^ n3876 ;
  assign n3882 = n3880 ^ x8 ;
  assign n3883 = n3882 ^ n3880 ;
  assign n3884 = n3883 ^ n252 ;
  assign n3885 = ~n3881 & n3884 ;
  assign n3886 = n3885 ^ n3876 ;
  assign n3887 = n252 & n3886 ;
  assign n3888 = ~n3873 & ~n3887 ;
  assign n3889 = n1994 & ~n3888 ;
  assign n3890 = n2931 & n3821 ;
  assign n3891 = n249 & n1709 ;
  assign n3892 = n1706 & n3848 ;
  assign n3893 = ~n3891 & ~n3892 ;
  assign n3894 = ~n1529 & ~n3893 ;
  assign n3895 = ~n1716 & ~n3592 ;
  assign n3896 = ~x2 & n3294 ;
  assign n3897 = n2928 & n3896 ;
  assign n3898 = ~n3895 & ~n3897 ;
  assign n3899 = ~n3894 & n3898 ;
  assign n3900 = ~n3890 & n3899 ;
  assign n3901 = n943 & ~n3900 ;
  assign n3902 = n3154 & n3452 ;
  assign n3903 = n210 & n1256 ;
  assign n3904 = n2309 & n3903 ;
  assign n3905 = ~n3902 & ~n3904 ;
  assign n3906 = n1376 & ~n3905 ;
  assign n3907 = n2041 & n3906 ;
  assign n3908 = ~n3901 & ~n3907 ;
  assign n3909 = ~n3889 & n3908 ;
  assign n3910 = n469 & ~n3909 ;
  assign n3911 = n3910 ^ n3863 ;
  assign n3912 = n77 & n1643 ;
  assign n3913 = x0 & ~n2560 ;
  assign n3914 = ~n2559 & n3913 ;
  assign n3915 = ~n3912 & ~n3914 ;
  assign n3916 = n1991 & ~n3915 ;
  assign n3917 = ~n1706 & n3294 ;
  assign n3918 = n2503 & n3917 ;
  assign n3919 = ~n77 & ~n1669 ;
  assign n3920 = n1760 & ~n3919 ;
  assign n3921 = ~n1376 & n3920 ;
  assign n3922 = ~n3918 & ~n3921 ;
  assign n3923 = ~n3916 & n3922 ;
  assign n3924 = n3508 & ~n3923 ;
  assign n3925 = ~n1798 & ~n3220 ;
  assign n3926 = x10 & n252 ;
  assign n3927 = n2549 & n3926 ;
  assign n3928 = n3925 & ~n3927 ;
  assign n3929 = n2156 & ~n3928 ;
  assign n3930 = ~n1797 & ~n3329 ;
  assign n3931 = n2445 & ~n3930 ;
  assign n3932 = n1784 & n2655 ;
  assign n3933 = ~n3931 & ~n3932 ;
  assign n3934 = ~n3929 & n3933 ;
  assign n3935 = n3282 & ~n3934 ;
  assign n3936 = n77 & n3021 ;
  assign n3937 = ~n1797 & ~n3936 ;
  assign n3938 = n3937 ^ n2282 ;
  assign n3939 = n3938 ^ n3937 ;
  assign n3940 = n3937 ^ n3925 ;
  assign n3941 = n3940 ^ n3937 ;
  assign n3942 = ~n3939 & ~n3941 ;
  assign n3943 = n3942 ^ n3937 ;
  assign n3944 = ~n2397 & ~n3943 ;
  assign n3945 = n3944 ^ n3937 ;
  assign n3946 = n570 & ~n3945 ;
  assign n3947 = ~n3935 & ~n3946 ;
  assign n3948 = ~n3924 & n3947 ;
  assign n3949 = n550 & ~n3948 ;
  assign n3950 = ~n1700 & n3824 ;
  assign n3951 = n62 & n1797 ;
  assign n3952 = ~n3950 & ~n3951 ;
  assign n3953 = x8 & ~n3952 ;
  assign n3954 = n252 & n1528 ;
  assign n3955 = ~n1629 & ~n3954 ;
  assign n3956 = ~n3953 & n3955 ;
  assign n3957 = n3956 ^ n252 ;
  assign n3958 = n3957 ^ n3956 ;
  assign n3959 = ~n1598 & ~n3849 ;
  assign n3960 = n3959 ^ n3956 ;
  assign n3961 = n3960 ^ n3956 ;
  assign n3962 = n3958 & ~n3961 ;
  assign n3963 = n3962 ^ n3956 ;
  assign n3964 = ~x0 & ~n3963 ;
  assign n3965 = n3964 ^ n3956 ;
  assign n3966 = n2548 & ~n3965 ;
  assign n3967 = x2 & ~x9 ;
  assign n3968 = n3220 & n3841 ;
  assign n3969 = ~x12 & n3643 ;
  assign n3970 = n267 & n1772 ;
  assign n3971 = n3969 & n3970 ;
  assign n3972 = ~x10 & n1668 ;
  assign n3973 = ~x0 & n3972 ;
  assign n3974 = ~n3971 & ~n3973 ;
  assign n3975 = ~n3968 & n3974 ;
  assign n3976 = n3967 & ~n3975 ;
  assign n3977 = ~x8 & n3970 ;
  assign n3978 = ~n3972 & ~n3977 ;
  assign n3979 = n2650 & ~n3978 ;
  assign n3980 = ~x4 & n267 ;
  assign n3981 = ~x6 & x14 ;
  assign n3982 = ~n3249 & ~n3981 ;
  assign n3983 = x4 & ~n3982 ;
  assign n3984 = ~n3980 & ~n3983 ;
  assign n3985 = n3095 & n3671 ;
  assign n3986 = ~n3984 & n3985 ;
  assign n3987 = ~n3979 & ~n3986 ;
  assign n3988 = n245 & n3021 ;
  assign n3989 = ~x12 & n1732 ;
  assign n3990 = n2741 & n3989 ;
  assign n3991 = ~n250 & ~n1376 ;
  assign n3992 = n3969 & n3991 ;
  assign n3993 = ~n3990 & ~n3992 ;
  assign n3994 = ~n3988 & n3993 ;
  assign n3995 = n286 & ~n3994 ;
  assign n3996 = n3987 & ~n3995 ;
  assign n3997 = ~n3976 & n3996 ;
  assign n3998 = ~n3966 & n3997 ;
  assign n3999 = n354 & ~n3998 ;
  assign n4000 = ~n1562 & n3509 ;
  assign n4001 = n4000 ^ x2 ;
  assign n4002 = n4001 ^ x0 ;
  assign n4010 = n4002 ^ n4001 ;
  assign n4003 = ~x0 & n1394 ;
  assign n4004 = n4003 ^ n4002 ;
  assign n4005 = n4004 ^ n4001 ;
  assign n4006 = n4002 ^ n4000 ;
  assign n4007 = n4006 ^ n4003 ;
  assign n4008 = n4007 ^ n4005 ;
  assign n4009 = n4005 & ~n4008 ;
  assign n4011 = n4010 ^ n4009 ;
  assign n4012 = n4011 ^ n4005 ;
  assign n4013 = n4001 ^ n1698 ;
  assign n4014 = n4009 ^ n4005 ;
  assign n4015 = n4013 & n4014 ;
  assign n4016 = n4015 ^ n4001 ;
  assign n4017 = ~n4012 & n4016 ;
  assign n4018 = n4017 ^ n4001 ;
  assign n4019 = n4018 ^ x2 ;
  assign n4020 = n4019 ^ n4001 ;
  assign n4021 = n249 & n4020 ;
  assign n4022 = n62 & n1702 ;
  assign n4023 = n246 & ~n4022 ;
  assign n4024 = n18 & ~n4023 ;
  assign n4025 = n4024 ^ x12 ;
  assign n4026 = n1749 ^ x8 ;
  assign n4027 = n4026 ^ n1749 ;
  assign n4028 = n1489 & n1715 ;
  assign n4029 = ~n1733 & ~n4028 ;
  assign n4030 = n4029 ^ n1749 ;
  assign n4031 = n4027 & ~n4030 ;
  assign n4032 = n4031 ^ n1749 ;
  assign n4033 = n4032 ^ n4024 ;
  assign n4034 = n4025 & ~n4033 ;
  assign n4035 = n4034 ^ n4031 ;
  assign n4036 = n4035 ^ n1749 ;
  assign n4037 = n4036 ^ x12 ;
  assign n4038 = ~n4024 & ~n4037 ;
  assign n4039 = n4038 ^ n4024 ;
  assign n4040 = n4039 ^ n4024 ;
  assign n4041 = n252 & ~n4040 ;
  assign n4042 = ~n4021 & ~n4041 ;
  assign n4043 = n934 & ~n4042 ;
  assign n4044 = ~n3999 & ~n4043 ;
  assign n4045 = ~n2278 & n3021 ;
  assign n4046 = ~n78 & n4045 ;
  assign n4047 = ~n20 & ~n2598 ;
  assign n4048 = n278 & n2309 ;
  assign n4049 = ~n4047 & n4048 ;
  assign n4050 = n4049 ^ n2746 ;
  assign n4051 = n4050 ^ n2746 ;
  assign n4052 = ~x4 & ~x8 ;
  assign n4053 = n1248 & n3249 ;
  assign n4054 = n4052 & n4053 ;
  assign n4055 = n4054 ^ n2746 ;
  assign n4056 = n4055 ^ n2746 ;
  assign n4057 = ~n4051 & ~n4056 ;
  assign n4058 = n4057 ^ n2746 ;
  assign n4059 = x10 & ~n4058 ;
  assign n4060 = n4059 ^ n2746 ;
  assign n4061 = ~n4046 & ~n4060 ;
  assign n4062 = n3068 & ~n4061 ;
  assign n4063 = n313 & n4062 ;
  assign n4064 = ~x0 & n2277 ;
  assign n4065 = n2536 & n4064 ;
  assign n4066 = n1667 & n2566 ;
  assign n4067 = ~n4065 & ~n4066 ;
  assign n4068 = n2388 & ~n4067 ;
  assign n4069 = n308 & n4068 ;
  assign n4070 = ~n4063 & ~n4069 ;
  assign n4071 = n4044 & n4070 ;
  assign n4072 = ~n3949 & n4071 ;
  assign n4073 = n4072 ^ x13 ;
  assign n4074 = n4073 ^ n4072 ;
  assign n4075 = n1257 & n3203 ;
  assign n4076 = n3201 & n3217 ;
  assign n4077 = ~n4075 & ~n4076 ;
  assign n4078 = n2709 & ~n4077 ;
  assign n4079 = n1257 & n3194 ;
  assign n4080 = n3197 & n3217 ;
  assign n4081 = ~n4079 & ~n4080 ;
  assign n4082 = n2704 & ~n4081 ;
  assign n4083 = ~n4078 & ~n4082 ;
  assign n4084 = ~x3 & ~n4083 ;
  assign n4085 = n1394 & n4028 ;
  assign n4086 = n3217 & n4064 ;
  assign n4087 = ~n4085 & ~n4086 ;
  assign n4088 = n934 & ~n4087 ;
  assign n4089 = ~n4084 & ~n4088 ;
  assign n4090 = n1352 & ~n4089 ;
  assign n4091 = n4090 ^ n4072 ;
  assign n4092 = n4074 & ~n4091 ;
  assign n4093 = n4092 ^ n4072 ;
  assign n4094 = n4093 ^ n3863 ;
  assign n4095 = n3911 & ~n4094 ;
  assign n4096 = n4095 ^ n4092 ;
  assign n4097 = n4096 ^ n4072 ;
  assign n4098 = n4097 ^ n3910 ;
  assign n4099 = ~n3863 & ~n4098 ;
  assign n4100 = n4099 ^ n3863 ;
  assign n4101 = n4100 ^ x11 ;
  assign n4102 = n4101 ^ n4100 ;
  assign n4103 = n294 & ~n2602 ;
  assign n4104 = ~n2878 & ~n4103 ;
  assign n4105 = ~n3521 & n4104 ;
  assign n4106 = n3643 & ~n4105 ;
  assign n4107 = n1493 & n3649 ;
  assign n4108 = n266 & n4107 ;
  assign n4109 = n1826 & n2715 ;
  assign n4110 = ~n4108 & ~n4109 ;
  assign n4111 = ~n4106 & n4110 ;
  assign n4112 = n436 & ~n4111 ;
  assign n4113 = ~x3 & n252 ;
  assign n4114 = ~x13 & n2558 ;
  assign n4115 = n1715 & n4114 ;
  assign n4116 = n768 & n2277 ;
  assign n4117 = x14 & n1394 ;
  assign n4118 = n638 & n4117 ;
  assign n4119 = ~n4116 & ~n4118 ;
  assign n4120 = ~n4115 & n4119 ;
  assign n4121 = n4113 & ~n4120 ;
  assign n4122 = ~n58 & ~n2549 ;
  assign n4123 = n529 & n4122 ;
  assign n4124 = ~x6 & n31 ;
  assign n4125 = n4123 & n4124 ;
  assign n4126 = n2277 & n4125 ;
  assign n4127 = ~n4121 & ~n4126 ;
  assign n4128 = ~n4112 & n4127 ;
  assign n4129 = n2041 & ~n4128 ;
  assign n4130 = n86 & n355 ;
  assign n4131 = n3044 & n4130 ;
  assign n4132 = n86 & n3294 ;
  assign n4133 = n2598 & n4132 ;
  assign n4134 = ~x6 & n266 ;
  assign n4135 = ~n2570 & ~n4134 ;
  assign n4136 = n655 & ~n4135 ;
  assign n4137 = ~n4133 & ~n4136 ;
  assign n4138 = ~n2915 & n4137 ;
  assign n4139 = n1493 & ~n4138 ;
  assign n4140 = x12 & n2746 ;
  assign n4141 = ~n62 & n1550 ;
  assign n4142 = ~n246 & n306 ;
  assign n4143 = n4141 & n4142 ;
  assign n4144 = ~n3246 & ~n3255 ;
  assign n4145 = n1932 & ~n4144 ;
  assign n4146 = ~n4143 & ~n4145 ;
  assign n4147 = ~n4140 & n4146 ;
  assign n4148 = ~n4139 & n4147 ;
  assign n4149 = n934 & ~n4148 ;
  assign n4150 = ~n4131 & ~n4149 ;
  assign n4151 = n1581 & n2906 ;
  assign n4152 = x2 & ~n58 ;
  assign n4153 = x0 & n62 ;
  assign n4154 = ~n4152 & ~n4153 ;
  assign n4155 = n4151 & ~n4154 ;
  assign n4156 = n2038 ^ n880 ;
  assign n4157 = n4156 ^ n2038 ;
  assign n4158 = n2038 ^ x2 ;
  assign n4159 = n4158 ^ n2038 ;
  assign n4160 = n4157 & n4159 ;
  assign n4161 = n4160 ^ n2038 ;
  assign n4162 = ~x8 & ~n4161 ;
  assign n4163 = n4162 ^ n2038 ;
  assign n4164 = x0 & ~n4163 ;
  assign n4165 = ~n221 & ~n2415 ;
  assign n4166 = ~n62 & n4165 ;
  assign n4167 = n252 & ~n4166 ;
  assign n4168 = ~x14 & n655 ;
  assign n4169 = n2397 & ~n4168 ;
  assign n4170 = n4167 & ~n4169 ;
  assign n4171 = ~n4164 & n4170 ;
  assign n4172 = ~n4155 & ~n4171 ;
  assign n4173 = x13 & ~n4172 ;
  assign n4174 = x1 & n4140 ;
  assign n4175 = ~n1365 & ~n2857 ;
  assign n4176 = n3297 & ~n4175 ;
  assign n4177 = n1112 & n1540 ;
  assign n4178 = ~n4176 & ~n4177 ;
  assign n4179 = n2038 & ~n4178 ;
  assign n4180 = ~n4174 & ~n4179 ;
  assign n4181 = ~n4173 & n4180 ;
  assign n4182 = n4181 ^ x1 ;
  assign n4183 = n4182 ^ n4181 ;
  assign n4184 = n1498 & n3295 ;
  assign n4185 = x6 & n153 ;
  assign n4186 = ~x8 & n3296 ;
  assign n4187 = n4185 & n4186 ;
  assign n4188 = n2124 & n3240 ;
  assign n4189 = ~n4187 & ~n4188 ;
  assign n4190 = ~n4184 & n4189 ;
  assign n4191 = n3314 & ~n4190 ;
  assign n4192 = n1248 & n1666 ;
  assign n4193 = n58 & n252 ;
  assign n4194 = n1608 & n4193 ;
  assign n4195 = ~n4192 & ~n4194 ;
  assign n4196 = ~x6 & n134 ;
  assign n4197 = n2586 & ~n2709 ;
  assign n4198 = ~x4 & ~n245 ;
  assign n4199 = n4197 & n4198 ;
  assign n4200 = n4196 & n4199 ;
  assign n4201 = n4195 & ~n4200 ;
  assign n4202 = ~n4191 & n4201 ;
  assign n4203 = n4202 ^ n4181 ;
  assign n4204 = n4203 ^ n4181 ;
  assign n4205 = n4183 & ~n4204 ;
  assign n4206 = n4205 ^ n4181 ;
  assign n4207 = x3 & ~n4206 ;
  assign n4208 = n4207 ^ n4181 ;
  assign n4209 = n4208 ^ x9 ;
  assign n4210 = n4209 ^ n4208 ;
  assign n4211 = n205 & ~n3314 ;
  assign n4212 = ~n2743 & n4211 ;
  assign n4213 = ~n1799 & n4212 ;
  assign n4214 = x6 & n2709 ;
  assign n4215 = x3 & n4214 ;
  assign n4216 = ~n4213 & ~n4215 ;
  assign n4217 = n1027 & ~n4216 ;
  assign n4218 = n85 & n799 ;
  assign n4219 = n269 & n4218 ;
  assign n4220 = ~n2282 & n4219 ;
  assign n4221 = n4220 ^ x1 ;
  assign n4222 = x3 & ~n2709 ;
  assign n4223 = ~n3283 & n4222 ;
  assign n4224 = ~n2309 & n4223 ;
  assign n4225 = ~n2549 & n2598 ;
  assign n4226 = n861 & n2743 ;
  assign n4227 = n4225 & ~n4226 ;
  assign n4228 = ~n4224 & n4227 ;
  assign n4229 = n1715 & ~n2223 ;
  assign n4230 = x8 & n4229 ;
  assign n4231 = n4230 ^ x3 ;
  assign n4232 = n4230 ^ n267 ;
  assign n4233 = n4232 ^ n267 ;
  assign n4234 = n4233 ^ n4231 ;
  assign n4235 = n3745 ^ n1702 ;
  assign n4236 = n3745 & n4235 ;
  assign n4237 = n4236 ^ n267 ;
  assign n4238 = n4237 ^ n3745 ;
  assign n4239 = ~n4234 & ~n4238 ;
  assign n4240 = n4239 ^ n4236 ;
  assign n4241 = n4240 ^ n3745 ;
  assign n4242 = n4231 & n4241 ;
  assign n4243 = n4242 ^ n4230 ;
  assign n4244 = ~n4228 & ~n4243 ;
  assign n4245 = n4244 ^ x4 ;
  assign n4246 = n4245 ^ n4244 ;
  assign n4247 = ~n267 & ~n269 ;
  assign n4248 = ~n2549 & n4247 ;
  assign n4249 = n1246 & n4248 ;
  assign n4250 = n2710 & n4249 ;
  assign n4251 = ~x0 & n1786 ;
  assign n4252 = ~x14 & n1669 ;
  assign n4253 = n4251 & n4252 ;
  assign n4254 = n85 & n269 ;
  assign n4255 = ~n2240 & ~n4254 ;
  assign n4256 = n2277 & ~n4255 ;
  assign n4257 = ~n4253 & ~n4256 ;
  assign n4258 = ~n4250 & n4257 ;
  assign n4259 = n4258 ^ n4244 ;
  assign n4260 = n4246 & n4259 ;
  assign n4261 = n4260 ^ n4244 ;
  assign n4262 = n4261 ^ n4220 ;
  assign n4263 = ~n4221 & n4262 ;
  assign n4264 = n4263 ^ n4260 ;
  assign n4265 = n4264 ^ n4244 ;
  assign n4266 = n4265 ^ x1 ;
  assign n4267 = ~n4220 & ~n4266 ;
  assign n4268 = n4267 ^ n4220 ;
  assign n4269 = n4268 ^ n4220 ;
  assign n4270 = ~n4217 & n4269 ;
  assign n4271 = n153 & ~n4270 ;
  assign n4272 = n252 & n2587 ;
  assign n4273 = ~n2781 & ~n4272 ;
  assign n4274 = n3508 ^ n2709 ;
  assign n4275 = n817 & n3048 ;
  assign n4276 = n4275 ^ n4274 ;
  assign n4277 = n4276 ^ n2709 ;
  assign n4278 = n4277 ^ n4276 ;
  assign n4279 = n4276 ^ n2888 ;
  assign n4280 = n4279 ^ n4274 ;
  assign n4281 = n4278 & ~n4280 ;
  assign n4282 = n4281 ^ n2888 ;
  assign n4283 = ~n1084 & ~n2888 ;
  assign n4284 = n4283 ^ n4274 ;
  assign n4285 = ~n4282 & ~n4284 ;
  assign n4286 = n4285 ^ n4283 ;
  assign n4287 = ~n4274 & n4286 ;
  assign n4288 = n4287 ^ n4281 ;
  assign n4289 = n4288 ^ n3508 ;
  assign n4290 = n4289 ^ n2888 ;
  assign n4291 = ~n4273 & ~n4290 ;
  assign n4292 = n24 & n2610 ;
  assign n4293 = n3161 & ~n3984 ;
  assign n4294 = ~x1 & n252 ;
  assign n4295 = n2739 & n4294 ;
  assign n4296 = ~n4151 & ~n4295 ;
  assign n4297 = ~n4293 & n4296 ;
  assign n4298 = ~x0 & ~n4297 ;
  assign n4299 = ~n4292 & ~n4298 ;
  assign n4300 = n49 & n1246 ;
  assign n4301 = n153 & n1823 ;
  assign n4302 = ~n4300 & ~n4301 ;
  assign n4303 = ~n4299 & ~n4302 ;
  assign n4304 = ~x12 & ~n1716 ;
  assign n4305 = ~n2762 & n3797 ;
  assign n4306 = n832 & ~n1674 ;
  assign n4307 = n1084 & n4306 ;
  assign n4308 = ~n4305 & ~n4307 ;
  assign n4309 = n4304 & ~n4308 ;
  assign n4310 = n861 & n2309 ;
  assign n4311 = n249 & n4310 ;
  assign n4312 = x2 & x13 ;
  assign n4313 = n880 & n4312 ;
  assign n4314 = n4311 & n4313 ;
  assign n4315 = ~n4309 & ~n4314 ;
  assign n4316 = ~n4303 & n4315 ;
  assign n4317 = ~n4291 & n4316 ;
  assign n4318 = ~n4271 & n4317 ;
  assign n4319 = n4318 ^ n4208 ;
  assign n4320 = n4210 & n4319 ;
  assign n4321 = n4320 ^ n4208 ;
  assign n4322 = n4150 & n4321 ;
  assign n4323 = ~n4129 & n4322 ;
  assign n4324 = ~x10 & ~n4323 ;
  assign n4325 = ~x14 & n2168 ;
  assign n4326 = n1644 & n4325 ;
  assign n4327 = ~x9 & n249 ;
  assign n4328 = n1493 & n4327 ;
  assign n4329 = ~n4326 & ~n4328 ;
  assign n4330 = ~n558 & ~n4329 ;
  assign n4331 = n675 & n2858 ;
  assign n4332 = n1079 & n2483 ;
  assign n4333 = ~n4331 & ~n4332 ;
  assign n4334 = n2415 & ~n4333 ;
  assign n4335 = n1084 & n2119 ;
  assign n4336 = ~n2544 & n4335 ;
  assign n4337 = ~n4334 & ~n4336 ;
  assign n4338 = ~n4330 & n4337 ;
  assign n4339 = n3903 & ~n4338 ;
  assign n4340 = n3314 & n3824 ;
  assign n4341 = x6 & n1234 ;
  assign n4342 = n292 & n4341 ;
  assign n4343 = ~n4340 & ~n4342 ;
  assign n4344 = n817 & ~n4343 ;
  assign n4345 = n1563 & n2938 ;
  assign n4346 = ~n4344 & ~n4345 ;
  assign n4347 = n861 & ~n4346 ;
  assign n4348 = ~x3 & n210 ;
  assign n4349 = n717 & n2661 ;
  assign n4350 = n4348 & n4349 ;
  assign n4351 = n1249 & n1563 ;
  assign n4352 = n1027 & n4351 ;
  assign n4353 = ~n4350 & ~n4352 ;
  assign n4354 = ~n4347 & n4353 ;
  assign n4355 = n2445 & ~n4354 ;
  assign n4356 = n1507 & n2501 ;
  assign n4357 = n1931 & n2741 ;
  assign n4358 = n1668 & n2039 ;
  assign n4359 = n1775 & n2415 ;
  assign n4360 = ~n1826 & n4359 ;
  assign n4361 = n2536 & n4360 ;
  assign n4362 = ~n4358 & ~n4361 ;
  assign n4363 = ~n4357 & n4362 ;
  assign n4364 = ~n4356 & n4363 ;
  assign n4365 = n2168 & ~n4364 ;
  assign n4366 = n3232 & n4365 ;
  assign n4367 = ~n4355 & ~n4366 ;
  assign n4368 = ~n4339 & n4367 ;
  assign n4369 = ~n4324 & n4368 ;
  assign n4370 = n4369 ^ n4100 ;
  assign n4371 = ~n4102 & ~n4370 ;
  assign n4372 = n4371 ^ n4100 ;
  assign n4373 = ~n3836 & ~n4372 ;
  assign n4374 = ~n3818 & n4373 ;
  assign n4375 = x15 & ~n4374 ;
  assign n4376 = ~n2038 & ~n2075 ;
  assign n4377 = n425 & n570 ;
  assign n4378 = n4376 & n4377 ;
  assign n4379 = n775 & ~n2483 ;
  assign n4380 = n4379 ^ n2105 ;
  assign n4381 = n4379 ^ x2 ;
  assign n4382 = n4381 ^ x2 ;
  assign n4383 = ~n133 & n538 ;
  assign n4384 = ~n3282 & n4383 ;
  assign n4385 = ~n2038 & ~n4384 ;
  assign n4386 = n4385 ^ x2 ;
  assign n4387 = ~n4382 & n4386 ;
  assign n4388 = n4387 ^ x2 ;
  assign n4389 = n4380 & n4388 ;
  assign n4390 = n4389 ^ n2105 ;
  assign n4391 = ~n4378 & ~n4390 ;
  assign n4392 = x4 & ~n4391 ;
  assign n4393 = n306 & n943 ;
  assign n4394 = ~x4 & n2126 ;
  assign n4395 = ~x2 & n4394 ;
  assign n4396 = ~n4393 & ~n4395 ;
  assign n4397 = ~n3103 & ~n4396 ;
  assign n4398 = ~x9 & n3056 ;
  assign n4399 = ~n4394 & ~n4398 ;
  assign n4400 = n2038 & ~n4399 ;
  assign n4401 = n3203 & n4341 ;
  assign n4402 = n62 & n943 ;
  assign n4403 = n3009 & n4402 ;
  assign n4404 = ~n4401 & ~n4403 ;
  assign n4405 = ~n4400 & n4404 ;
  assign n4406 = n88 & ~n4405 ;
  assign n4407 = ~n1366 & ~n4047 ;
  assign n4408 = ~n364 & ~n2038 ;
  assign n4409 = ~n2181 & n2950 ;
  assign n4410 = ~n4408 & n4409 ;
  assign n4411 = ~n4407 & n4410 ;
  assign n4412 = ~n4406 & ~n4411 ;
  assign n4413 = ~n4397 & n4412 ;
  assign n4414 = ~n4392 & n4413 ;
  assign n4415 = x3 & ~n4414 ;
  assign n4416 = n67 & n3203 ;
  assign n4417 = n4124 & n4416 ;
  assign n4418 = ~x12 & n39 ;
  assign n4419 = ~n603 & ~n3282 ;
  assign n4420 = ~n2587 & n4419 ;
  assign n4421 = ~n3446 & ~n3824 ;
  assign n4422 = ~n4420 & ~n4421 ;
  assign n4423 = ~n817 & ~n2387 ;
  assign n4424 = x11 ^ x9 ;
  assign n4425 = n4424 ^ n4423 ;
  assign n4426 = n3508 ^ x12 ;
  assign n4427 = ~x11 & ~n4426 ;
  assign n4428 = n4427 ^ x12 ;
  assign n4429 = ~n4425 & ~n4428 ;
  assign n4430 = n4429 ^ n4427 ;
  assign n4431 = n4430 ^ x12 ;
  assign n4432 = n4431 ^ x11 ;
  assign n4433 = ~n4423 & n4432 ;
  assign n4434 = n4422 & n4433 ;
  assign n4435 = ~n4418 & n4434 ;
  assign n4436 = ~n4417 & ~n4435 ;
  assign n4437 = ~x8 & n4436 ;
  assign n4438 = ~n4415 & n4437 ;
  assign n4439 = x9 ^ x6 ;
  assign n4440 = n3085 ^ x9 ;
  assign n4441 = n4440 ^ n3085 ;
  assign n4442 = ~x11 & ~n679 ;
  assign n4443 = n4442 ^ n3085 ;
  assign n4444 = n4441 & n4443 ;
  assign n4445 = n4444 ^ n3085 ;
  assign n4446 = n4439 & ~n4445 ;
  assign n4447 = n4446 ^ x6 ;
  assign n4448 = n792 & n4447 ;
  assign n4449 = n252 & n2041 ;
  assign n4450 = n933 & n4449 ;
  assign n4451 = n49 & n3069 ;
  assign n4452 = ~n1728 & ~n4451 ;
  assign n4453 = x12 & n1731 ;
  assign n4454 = n4452 & ~n4453 ;
  assign n4455 = n2661 & ~n4454 ;
  assign n4456 = ~n4450 & ~n4455 ;
  assign n4457 = x9 & ~n4442 ;
  assign n4458 = x6 & n2660 ;
  assign n4459 = n4457 & n4458 ;
  assign n4460 = ~n109 & ~n4383 ;
  assign n4461 = n4460 ^ x9 ;
  assign n4462 = n4461 ^ n4460 ;
  assign n4463 = n4462 ^ n249 ;
  assign n4464 = n819 ^ x11 ;
  assign n4465 = ~n819 & n4464 ;
  assign n4466 = n4465 ^ n4460 ;
  assign n4467 = n4466 ^ n819 ;
  assign n4468 = n4463 & ~n4467 ;
  assign n4469 = n4468 ^ n4465 ;
  assign n4470 = n4469 ^ n819 ;
  assign n4471 = n249 & ~n4470 ;
  assign n4472 = n4471 ^ n249 ;
  assign n4473 = ~n4459 & ~n4472 ;
  assign n4474 = n4456 & n4473 ;
  assign n4475 = ~n4448 & n4474 ;
  assign n4476 = n1786 & ~n4475 ;
  assign n4477 = n38 & n249 ;
  assign n4478 = n34 & n396 ;
  assign n4479 = n4477 & n4478 ;
  assign n4488 = n2548 & n3446 ;
  assign n4489 = ~n99 & n4488 ;
  assign n4490 = n249 ^ x2 ;
  assign n4491 = n4490 ^ n249 ;
  assign n4492 = n2565 & n2647 ;
  assign n4493 = n4492 ^ n249 ;
  assign n4494 = n4491 & n4493 ;
  assign n4495 = n4494 ^ n249 ;
  assign n4496 = x13 & n4495 ;
  assign n4497 = n67 & n4496 ;
  assign n4498 = x1 & n4312 ;
  assign n4499 = x9 & n1438 ;
  assign n4500 = ~x6 & x11 ;
  assign n4501 = n4499 & n4500 ;
  assign n4502 = n2565 & n4341 ;
  assign n4503 = ~n4501 & ~n4502 ;
  assign n4504 = n4498 & ~n4503 ;
  assign n4505 = ~x2 & x12 ;
  assign n4506 = x13 & n4505 ;
  assign n4507 = n4449 & n4506 ;
  assign n4508 = ~n4504 & ~n4507 ;
  assign n4509 = ~n4497 & n4508 ;
  assign n4510 = ~n4489 & n4509 ;
  assign n4480 = ~n3453 & n4449 ;
  assign n4481 = ~n214 & ~n603 ;
  assign n4482 = n571 & ~n4481 ;
  assign n4483 = ~x9 & n3085 ;
  assign n4484 = ~n437 & ~n4483 ;
  assign n4485 = ~n4482 & n4484 ;
  assign n4486 = n249 & ~n4485 ;
  assign n4487 = ~n4480 & ~n4486 ;
  assign n4511 = n4510 ^ n4487 ;
  assign n4512 = n4511 ^ n4510 ;
  assign n4513 = n4510 ^ x2 ;
  assign n4514 = n4513 ^ n4510 ;
  assign n4515 = ~n4512 & n4514 ;
  assign n4516 = n4515 ^ n4510 ;
  assign n4517 = x3 & ~n4516 ;
  assign n4518 = n4517 ^ n4510 ;
  assign n4519 = ~n4479 & n4518 ;
  assign n4520 = x8 & n4519 ;
  assign n4521 = ~n4476 & n4520 ;
  assign n4522 = ~n4438 & ~n4521 ;
  assign n4523 = n775 & n1957 ;
  assign n4524 = x3 & n2079 ;
  assign n4525 = ~x2 & n4524 ;
  assign n4526 = ~n4523 & ~n4525 ;
  assign n4527 = n4477 & ~n4526 ;
  assign n4528 = ~x10 & ~n4527 ;
  assign n4529 = ~n4522 & n4528 ;
  assign n4530 = n2156 & ~n3448 ;
  assign n4531 = ~n2124 & ~n4530 ;
  assign n4532 = ~x3 & ~n4531 ;
  assign n4533 = ~n2505 & ~n4532 ;
  assign n4534 = x11 & n252 ;
  assign n4535 = ~n4533 & n4534 ;
  assign n4536 = ~x9 & n1671 ;
  assign n4537 = n28 & n4536 ;
  assign n4538 = ~n460 & n2223 ;
  assign n4539 = n1599 & ~n3453 ;
  assign n4540 = n4538 & n4539 ;
  assign n4541 = ~n4537 & ~n4540 ;
  assign n4542 = n4541 ^ x4 ;
  assign n4543 = n4542 ^ n4541 ;
  assign n4544 = n4543 ^ n4535 ;
  assign n4545 = ~n34 & ~n604 ;
  assign n4546 = ~n215 & n4545 ;
  assign n4547 = n1671 & ~n4546 ;
  assign n4548 = n1503 & n1728 ;
  assign n4549 = ~n2503 & ~n4548 ;
  assign n4550 = ~n4547 & n4549 ;
  assign n4551 = n4550 ^ x3 ;
  assign n4552 = ~n4550 & ~n4551 ;
  assign n4553 = n4552 ^ n4541 ;
  assign n4554 = n4553 ^ n4550 ;
  assign n4555 = n4544 & n4554 ;
  assign n4556 = n4555 ^ n4552 ;
  assign n4557 = n4556 ^ n4550 ;
  assign n4558 = ~n4535 & ~n4557 ;
  assign n4559 = n4558 ^ n4535 ;
  assign n4560 = n2038 & n4559 ;
  assign n4561 = ~x4 & x9 ;
  assign n4562 = n556 & n4561 ;
  assign n4563 = ~x6 & n88 ;
  assign n4564 = n4562 & n4563 ;
  assign n4565 = n2405 & n4564 ;
  assign n4566 = x10 & ~n4565 ;
  assign n4567 = ~n4560 & n4566 ;
  assign n4568 = ~n3069 & n4341 ;
  assign n4569 = x12 & ~n2565 ;
  assign n4570 = n3422 & ~n4569 ;
  assign n4571 = ~n4568 & ~n4570 ;
  assign n4572 = n2276 & ~n4571 ;
  assign n4573 = x9 & ~x14 ;
  assign n4574 = ~n253 & ~n4573 ;
  assign n4575 = n3162 & ~n4574 ;
  assign n4576 = n4575 ^ n249 ;
  assign n4577 = n3068 ^ n252 ;
  assign n4578 = n4575 ^ n252 ;
  assign n4579 = n4578 ^ n252 ;
  assign n4580 = ~n4577 & ~n4579 ;
  assign n4581 = n4580 ^ n252 ;
  assign n4582 = n4576 & n4581 ;
  assign n4583 = n4582 ^ n249 ;
  assign n4584 = n2277 & n4583 ;
  assign n4585 = ~n4572 & ~n4584 ;
  assign n4586 = n909 & ~n4585 ;
  assign n4587 = x11 & ~n1376 ;
  assign n4588 = n528 & n1298 ;
  assign n4589 = ~x2 & ~n4588 ;
  assign n4590 = n1404 & ~n4589 ;
  assign n4591 = n4587 & n4590 ;
  assign n4592 = ~n49 & ~n62 ;
  assign n4593 = ~x8 & n4592 ;
  assign n4594 = n4134 & n4593 ;
  assign n4595 = n228 & n1669 ;
  assign n4596 = ~n3448 & n4595 ;
  assign n4597 = ~n4594 & ~n4596 ;
  assign n4598 = n2079 & ~n4597 ;
  assign n4599 = ~n4591 & ~n4598 ;
  assign n4600 = x3 & ~n4599 ;
  assign n4601 = n67 & n2601 ;
  assign n4602 = n1404 & n4601 ;
  assign n4603 = ~n4600 & ~n4602 ;
  assign n4604 = ~n4586 & n4603 ;
  assign n4605 = n4604 ^ x1 ;
  assign n4606 = n4605 ^ n4604 ;
  assign n4607 = n4606 ^ n4567 ;
  assign n4608 = ~x3 & x4 ;
  assign n4609 = n528 & n2445 ;
  assign n4610 = n1260 & n4609 ;
  assign n4611 = ~n2503 & ~n4610 ;
  assign n4612 = n4608 & ~n4611 ;
  assign n4613 = ~n153 & ~n2777 ;
  assign n4615 = n4613 ^ x3 ;
  assign n4614 = n4613 ^ n1669 ;
  assign n4616 = n4615 ^ n4614 ;
  assign n4617 = n4616 ^ n4615 ;
  assign n4618 = n4617 ^ n4613 ;
  assign n4619 = x4 & ~n133 ;
  assign n4620 = n4619 ^ n4616 ;
  assign n4621 = ~x9 & n4620 ;
  assign n4622 = n4615 ^ n4613 ;
  assign n4623 = ~n4617 & ~n4622 ;
  assign n4624 = n4623 ^ n4618 ;
  assign n4625 = n4621 & n4624 ;
  assign n4626 = n4625 ^ n4623 ;
  assign n4627 = n4618 & n4626 ;
  assign n4628 = n4627 ^ n4623 ;
  assign n4629 = n4628 ^ x3 ;
  assign n4630 = ~n4612 & n4629 ;
  assign n4631 = x11 & ~n4630 ;
  assign n4632 = n252 & n1404 ;
  assign n4633 = ~x11 & n4632 ;
  assign n4634 = ~n3453 & n4633 ;
  assign n4635 = n4634 ^ x3 ;
  assign n4636 = ~x9 & ~n4588 ;
  assign n4637 = n4587 & ~n4636 ;
  assign n4638 = n1366 & n3824 ;
  assign n4639 = ~n4637 & ~n4638 ;
  assign n4640 = n4639 ^ x8 ;
  assign n4641 = n4640 ^ n4639 ;
  assign n4642 = n890 & n1699 ;
  assign n4643 = n4545 & ~n4642 ;
  assign n4644 = n1376 & ~n4643 ;
  assign n4645 = ~x6 & n570 ;
  assign n4646 = n2877 & n4645 ;
  assign n4647 = n4646 ^ x11 ;
  assign n4648 = n4647 ^ n4646 ;
  assign n4649 = n4648 ^ n4394 ;
  assign n4650 = n2585 ^ n38 ;
  assign n4651 = n2585 & n4650 ;
  assign n4652 = n4651 ^ n4646 ;
  assign n4653 = n4652 ^ n2585 ;
  assign n4654 = n4649 & n4653 ;
  assign n4655 = n4654 ^ n4651 ;
  assign n4656 = n4655 ^ n2585 ;
  assign n4657 = ~n4394 & n4656 ;
  assign n4658 = n4657 ^ n4394 ;
  assign n4659 = ~n4644 & ~n4658 ;
  assign n4660 = n4659 ^ n4639 ;
  assign n4661 = ~n4641 & n4660 ;
  assign n4662 = n4661 ^ n4639 ;
  assign n4663 = n4662 ^ n4634 ;
  assign n4664 = ~n4635 & n4663 ;
  assign n4665 = n4664 ^ n4661 ;
  assign n4666 = n4665 ^ n4639 ;
  assign n4667 = n4666 ^ x3 ;
  assign n4668 = ~n4634 & ~n4667 ;
  assign n4669 = n4668 ^ n4634 ;
  assign n4670 = n4669 ^ n4634 ;
  assign n4671 = ~n4631 & n4670 ;
  assign n4672 = n4671 ^ x2 ;
  assign n4673 = ~n4671 & n4672 ;
  assign n4674 = n4673 ^ n4604 ;
  assign n4675 = n4674 ^ n4671 ;
  assign n4676 = n4607 & n4675 ;
  assign n4677 = n4676 ^ n4673 ;
  assign n4678 = n4677 ^ n4671 ;
  assign n4679 = n4567 & ~n4678 ;
  assign n4680 = n4679 ^ n4567 ;
  assign n4681 = x0 & ~n4680 ;
  assign n4682 = ~n4529 & n4681 ;
  assign n4683 = n1797 & n2447 ;
  assign n4684 = ~n1252 & ~n1367 ;
  assign n4685 = n3021 & ~n4684 ;
  assign n4686 = ~n4683 & ~n4685 ;
  assign n4687 = n308 & ~n4686 ;
  assign n4688 = n1394 & n1797 ;
  assign n4689 = n313 & n4688 ;
  assign n4690 = n425 & n1598 ;
  assign n4691 = x1 & x8 ;
  assign n4692 = n4588 & n4691 ;
  assign n4693 = ~n4690 & ~n4692 ;
  assign n4694 = x3 & n1264 ;
  assign n4695 = ~n4693 & n4694 ;
  assign n4696 = n2640 & n4477 ;
  assign n4697 = x10 & n4696 ;
  assign n4698 = ~n4695 & ~n4697 ;
  assign n4699 = ~n4689 & n4698 ;
  assign n4700 = n1395 & n4113 ;
  assign n4701 = n308 & n1581 ;
  assign n4702 = n679 ^ n49 ;
  assign n4703 = n49 ^ x6 ;
  assign n4704 = n4703 ^ n49 ;
  assign n4705 = n4704 ^ n4701 ;
  assign n4706 = n4702 & n4705 ;
  assign n4707 = n4706 ^ n679 ;
  assign n4708 = n4701 & n4707 ;
  assign n4709 = ~n4700 & ~n4708 ;
  assign n4710 = n4709 ^ x10 ;
  assign n4711 = n4710 ^ n4709 ;
  assign n4712 = n4711 ^ n4699 ;
  assign n4713 = ~x12 & n425 ;
  assign n4714 = ~n1656 & ~n4713 ;
  assign n4715 = x4 & ~n4714 ;
  assign n4716 = n1542 & n3249 ;
  assign n4717 = ~n4715 & ~n4716 ;
  assign n4718 = n2678 & ~n4717 ;
  assign n4719 = n4718 ^ x1 ;
  assign n4720 = x1 & n4719 ;
  assign n4721 = n4720 ^ n4709 ;
  assign n4722 = n4721 ^ x1 ;
  assign n4723 = n4712 & ~n4722 ;
  assign n4724 = n4723 ^ n4720 ;
  assign n4725 = n4724 ^ x1 ;
  assign n4726 = n4699 & n4725 ;
  assign n4727 = n4726 ^ n4699 ;
  assign n4728 = n2079 & ~n4727 ;
  assign n4729 = n308 & n1551 ;
  assign n4730 = n503 & n1790 ;
  assign n4731 = ~n4729 & ~n4730 ;
  assign n4732 = n252 & ~n4731 ;
  assign n4733 = ~n1489 & n2942 ;
  assign n4734 = n550 & n4733 ;
  assign n4735 = ~n4732 & ~n4734 ;
  assign n4736 = n2886 & ~n4735 ;
  assign n4737 = x4 & x9 ;
  assign n4738 = x3 & n1672 ;
  assign n4739 = ~n403 & n2272 ;
  assign n4740 = ~n4738 & ~n4739 ;
  assign n4741 = n3172 & ~n4740 ;
  assign n4742 = n3161 ^ x10 ;
  assign n4743 = n2223 & n4742 ;
  assign n4744 = ~n4741 & ~n4743 ;
  assign n4745 = n4737 & ~n4744 ;
  assign n4746 = ~x1 & x10 ;
  assign n4747 = ~n3172 & ~n4746 ;
  assign n4748 = n1643 & n4747 ;
  assign n4749 = n38 & n4748 ;
  assign n4750 = ~n308 & n4749 ;
  assign n4751 = ~n4745 & ~n4750 ;
  assign n4752 = ~n2656 & ~n4294 ;
  assign n4753 = n153 & n2739 ;
  assign n4754 = x10 & n4753 ;
  assign n4755 = ~n4752 & n4754 ;
  assign n4756 = n1256 & n1619 ;
  assign n4757 = n2424 & n4756 ;
  assign n4758 = ~x10 & n4151 ;
  assign n4759 = ~n4757 & ~n4758 ;
  assign n4760 = ~n4755 & n4759 ;
  assign n4761 = n73 & ~n4760 ;
  assign n4762 = x8 & ~n153 ;
  assign n4763 = n3708 & n4762 ;
  assign n4764 = ~n3659 & ~n4763 ;
  assign n4765 = n3809 & ~n4764 ;
  assign n4766 = ~n550 & ~n4691 ;
  assign n4767 = ~n2410 & n2458 ;
  assign n4768 = ~n1285 & ~n4767 ;
  assign n4769 = ~n4766 & n4768 ;
  assign n4770 = ~n4765 & ~n4769 ;
  assign n4771 = n4561 & ~n4770 ;
  assign n4772 = ~n4761 & ~n4771 ;
  assign n4773 = n4751 & n4772 ;
  assign n4774 = ~x3 & n1256 ;
  assign n4775 = ~x12 & ~n1530 ;
  assign n4776 = n313 & n4775 ;
  assign n4777 = ~n4774 & ~n4776 ;
  assign n4778 = n252 & ~n4777 ;
  assign n4779 = n880 & ~n3708 ;
  assign n4780 = ~n426 & ~n4746 ;
  assign n4781 = ~n926 & n4780 ;
  assign n4782 = n249 & n4781 ;
  assign n4783 = ~n4779 & n4782 ;
  assign n4784 = ~n4778 & ~n4783 ;
  assign n4785 = n1550 & ~n4784 ;
  assign n4786 = ~n556 & n2660 ;
  assign n4787 = n1529 & n2410 ;
  assign n4788 = n4786 & n4787 ;
  assign n4789 = ~n4785 & ~n4788 ;
  assign n4790 = ~x9 & ~n4789 ;
  assign n4791 = n4773 & ~n4790 ;
  assign n4792 = ~n4736 & n4791 ;
  assign n4793 = n4792 ^ x11 ;
  assign n4794 = n4793 ^ n4792 ;
  assign n4795 = n742 & n3926 ;
  assign n4796 = n73 & n3107 ;
  assign n4797 = ~n4752 & n4796 ;
  assign n4798 = ~n4795 & ~n4797 ;
  assign n4799 = n1550 & ~n4798 ;
  assign n4800 = n1559 & n2445 ;
  assign n4801 = x9 & ~x10 ;
  assign n4802 = n4801 ^ n38 ;
  assign n4803 = n4802 ^ n4800 ;
  assign n4804 = n2157 ^ n1546 ;
  assign n4805 = ~n4801 & ~n4804 ;
  assign n4806 = n4805 ^ n1546 ;
  assign n4807 = ~n4803 & ~n4806 ;
  assign n4808 = n4807 ^ n4805 ;
  assign n4809 = n4808 ^ n1546 ;
  assign n4810 = n4809 ^ n4801 ;
  assign n4811 = ~n4800 & n4810 ;
  assign n4812 = n2661 & ~n4811 ;
  assign n4813 = ~n4799 & ~n4812 ;
  assign n4814 = n4477 & n4691 ;
  assign n4815 = n3701 ^ n62 ;
  assign n4816 = n2415 & n4124 ;
  assign n4817 = n4816 ^ n3701 ;
  assign n4818 = n4816 ^ n49 ;
  assign n4819 = ~n4816 & n4818 ;
  assign n4820 = n4819 ^ n4816 ;
  assign n4821 = n4817 & ~n4820 ;
  assign n4822 = n4821 ^ n4819 ;
  assign n4823 = n4822 ^ n4816 ;
  assign n4824 = n4823 ^ n49 ;
  assign n4825 = ~n4815 & n4824 ;
  assign n4826 = n4825 ^ n3701 ;
  assign n4827 = ~n4814 & ~n4826 ;
  assign n4828 = n1758 & ~n4827 ;
  assign n4829 = n4813 & ~n4828 ;
  assign n4830 = n4829 ^ n4792 ;
  assign n4831 = ~n4794 & n4830 ;
  assign n4832 = n4831 ^ n4792 ;
  assign n4833 = ~n4728 & n4832 ;
  assign n4834 = ~n4687 & n4833 ;
  assign n4835 = n1248 & ~n4834 ;
  assign n4836 = ~n4682 & ~n4835 ;
  assign n4837 = ~n4375 & n4836 ;
  assign n4838 = n3724 & n4837 ;
  assign n4839 = n3190 & n4838 ;
  assign n4840 = ~n752 & ~n4839 ;
  assign n4841 = ~n1946 & ~n2877 ;
  assign n4842 = n210 & n1503 ;
  assign n4843 = n1622 & n4842 ;
  assign n4844 = ~n4841 & n4843 ;
  assign n4845 = ~n200 & ~n284 ;
  assign n4846 = ~n1458 & n4845 ;
  assign n4847 = n2556 & n4846 ;
  assign n4848 = ~n4844 & ~n4847 ;
  assign n4849 = n473 & ~n4848 ;
  assign n4850 = n1248 & n1581 ;
  assign n4851 = n2397 ^ n1352 ;
  assign n4852 = n4851 ^ n2351 ;
  assign n4853 = n4852 ^ n2397 ;
  assign n4854 = n4853 ^ n4852 ;
  assign n4855 = n4852 ^ n3868 ;
  assign n4856 = n4855 ^ n4851 ;
  assign n4857 = n4854 & ~n4856 ;
  assign n4858 = n4857 ^ n3868 ;
  assign n4859 = ~n77 & ~n3868 ;
  assign n4860 = n4859 ^ n4851 ;
  assign n4861 = ~n4858 & n4860 ;
  assign n4862 = n4861 ^ n4859 ;
  assign n4863 = n4851 & n4862 ;
  assign n4864 = n4863 ^ n4857 ;
  assign n4865 = n4864 ^ n1352 ;
  assign n4866 = n4865 ^ n3868 ;
  assign n4867 = ~n4850 & ~n4866 ;
  assign n4868 = n2184 & ~n4867 ;
  assign n4869 = ~x0 & n207 ;
  assign n4870 = n3745 & n4869 ;
  assign n4871 = ~n2557 & ~n4870 ;
  assign n4872 = n25 & n88 ;
  assign n4873 = ~n4871 & n4872 ;
  assign n4874 = ~n4868 & ~n4873 ;
  assign n4875 = n207 & n2309 ;
  assign n4876 = n2555 & n4875 ;
  assign n4877 = ~x4 & n3488 ;
  assign n4878 = n207 & n1671 ;
  assign n4879 = ~n4877 & ~n4878 ;
  assign n4880 = n4879 ^ x0 ;
  assign n4881 = n4880 ^ n4879 ;
  assign n4882 = n4881 ^ n4876 ;
  assign n4883 = ~x4 & n2257 ;
  assign n4884 = n4883 ^ x8 ;
  assign n4885 = x8 & n4884 ;
  assign n4886 = n4885 ^ n4879 ;
  assign n4887 = n4886 ^ x8 ;
  assign n4888 = ~n4882 & ~n4887 ;
  assign n4889 = n4888 ^ n4885 ;
  assign n4890 = n4889 ^ x8 ;
  assign n4891 = ~n4876 & n4890 ;
  assign n4892 = n4891 ^ n4876 ;
  assign n4893 = n910 & n4892 ;
  assign n4894 = x5 & n4893 ;
  assign n4895 = n4874 & ~n4894 ;
  assign n4896 = ~n4849 & n4895 ;
  assign n4897 = n905 & ~n4896 ;
  assign n4898 = ~n1293 & n2282 ;
  assign n4899 = n1990 & n2397 ;
  assign n4900 = ~n4898 & ~n4899 ;
  assign n4901 = ~n79 & ~n4900 ;
  assign n4902 = n247 & n2558 ;
  assign n4903 = ~n4875 & ~n4902 ;
  assign n4904 = n25 & ~n4903 ;
  assign n4905 = ~n3462 & n4904 ;
  assign n4906 = ~n4901 & ~n4905 ;
  assign n4907 = n74 & ~n4906 ;
  assign n4908 = n22 & n909 ;
  assign n4909 = ~n2710 & n3317 ;
  assign n4910 = n3283 & n3728 ;
  assign n4911 = n2257 & n2549 ;
  assign n4912 = ~n4910 & ~n4911 ;
  assign n4913 = ~n2197 & ~n4912 ;
  assign n4914 = ~n4909 & ~n4913 ;
  assign n4915 = ~n2755 & n4914 ;
  assign n4916 = n4908 & ~n4915 ;
  assign n4917 = ~n4907 & ~n4916 ;
  assign n4918 = x1 & ~n4917 ;
  assign n4919 = x14 ^ x0 ;
  assign n4920 = n247 & n2386 ;
  assign n4921 = n1470 & n4920 ;
  assign n4922 = n1290 & n2138 ;
  assign n4923 = n74 & n4922 ;
  assign n4924 = n207 & n4923 ;
  assign n4925 = ~n4921 & ~n4924 ;
  assign n4926 = n4925 ^ x14 ;
  assign n4927 = n4926 ^ n4925 ;
  assign n4928 = n74 & n1630 ;
  assign n4929 = n1815 & n4928 ;
  assign n4930 = n1320 & n1611 ;
  assign n4931 = n1834 & n4930 ;
  assign n4932 = n425 & n4931 ;
  assign n4933 = ~n4929 & ~n4932 ;
  assign n4934 = n4933 ^ n4925 ;
  assign n4935 = ~n4927 & n4934 ;
  assign n4936 = n4935 ^ n4925 ;
  assign n4937 = n4919 & ~n4936 ;
  assign n4938 = ~n4918 & ~n4937 ;
  assign n4939 = x15 & ~n4938 ;
  assign n4949 = n292 & n2555 ;
  assign n4950 = n1619 & n4949 ;
  assign n4951 = n247 & n1669 ;
  assign n4952 = n77 & n4951 ;
  assign n4953 = ~n4950 & ~n4952 ;
  assign n4954 = n333 & n909 ;
  assign n4955 = n74 & n2123 ;
  assign n4956 = ~n4954 & ~n4955 ;
  assign n4957 = ~n4953 & ~n4956 ;
  assign n4958 = n2607 ^ x4 ;
  assign n4959 = n4958 ^ n2607 ;
  assign n4960 = n267 & n2397 ;
  assign n4961 = n4960 ^ n2607 ;
  assign n4962 = n4961 ^ n2607 ;
  assign n4963 = n4959 & n4962 ;
  assign n4964 = n4963 ^ n2607 ;
  assign n4965 = ~x0 & n4964 ;
  assign n4966 = n4965 ^ n2607 ;
  assign n4967 = n189 & n4966 ;
  assign n4968 = ~n1253 & n4967 ;
  assign n4969 = ~n4957 & ~n4968 ;
  assign n4940 = ~x1 & n909 ;
  assign n4941 = n266 & n1503 ;
  assign n4942 = ~n78 & ~n3652 ;
  assign n4943 = n4941 & ~n4942 ;
  assign n4944 = ~n269 & ~n1618 ;
  assign n4945 = n278 & n2282 ;
  assign n4946 = ~n4944 & n4945 ;
  assign n4947 = ~n4943 & ~n4946 ;
  assign n4948 = n4940 & ~n4947 ;
  assign n4970 = n4969 ^ n4948 ;
  assign n4971 = n4970 ^ n4969 ;
  assign n4972 = n4969 ^ x7 ;
  assign n4973 = n4972 ^ n4969 ;
  assign n4974 = n4971 & n4973 ;
  assign n4975 = n4974 ^ n4969 ;
  assign n4976 = ~x5 & ~n4975 ;
  assign n4977 = n4976 ^ n4969 ;
  assign n4978 = ~n4939 & n4977 ;
  assign n4979 = ~n4897 & n4978 ;
  assign n4980 = ~n457 & ~n4979 ;
  assign n4981 = n1376 & n2814 ;
  assign n4982 = n189 & n280 ;
  assign n4983 = x8 & n85 ;
  assign n4984 = n4982 & n4983 ;
  assign n4985 = n4981 & n4984 ;
  assign n4995 = n1248 & n4608 ;
  assign n4986 = n31 & n1273 ;
  assign n4987 = n1248 & n2739 ;
  assign n4988 = n4986 & n4987 ;
  assign n4989 = ~n2758 & ~n2867 ;
  assign n4990 = n1787 & ~n4989 ;
  assign n4991 = n1667 & n4990 ;
  assign n4992 = ~n4988 & ~n4991 ;
  assign n4996 = n4995 ^ n4992 ;
  assign n4997 = n4996 ^ n4992 ;
  assign n4993 = n4992 ^ n399 ;
  assign n4994 = n4993 ^ n4992 ;
  assign n4998 = n4997 ^ n4994 ;
  assign n4999 = n4992 ^ n1671 ;
  assign n5000 = n4999 ^ n4992 ;
  assign n5001 = n5000 ^ n4997 ;
  assign n5002 = n4997 & n5001 ;
  assign n5003 = n5002 ^ n4997 ;
  assign n5004 = n4998 & n5003 ;
  assign n5005 = n5004 ^ n5002 ;
  assign n5006 = n5005 ^ n4992 ;
  assign n5007 = n5006 ^ n4997 ;
  assign n5008 = x5 & ~n5007 ;
  assign n5009 = n5008 ^ n4992 ;
  assign n5010 = n4940 & ~n5009 ;
  assign n5011 = ~x2 & n308 ;
  assign n5012 = ~n1293 & n3474 ;
  assign n5013 = n1411 & n3473 ;
  assign n5014 = ~n5012 & ~n5013 ;
  assign n5015 = n5011 & ~n5014 ;
  assign n5016 = n1667 & n5015 ;
  assign n5017 = ~n5010 & ~n5016 ;
  assign n5018 = ~n4985 & n5017 ;
  assign n5019 = ~n2905 & ~n5018 ;
  assign n5020 = n1248 & n2610 ;
  assign n5021 = ~x2 & n3296 ;
  assign n5022 = n3745 & n5021 ;
  assign n5023 = ~n5020 & ~n5022 ;
  assign n5024 = ~n905 & n1085 ;
  assign n5025 = n149 & n892 ;
  assign n5026 = ~n5024 & n5025 ;
  assign n5027 = ~x11 & n475 ;
  assign n5028 = x5 & n5027 ;
  assign n5029 = n2123 & n5028 ;
  assign n5030 = n507 & n5029 ;
  assign n5031 = ~n321 & ~n2233 ;
  assign n5032 = n22 & n5031 ;
  assign n5033 = ~x13 & n918 ;
  assign n5034 = ~n5032 & ~n5033 ;
  assign n5035 = n4524 & ~n5034 ;
  assign n5036 = ~n5030 & ~n5035 ;
  assign n5037 = ~n5026 & n5036 ;
  assign n5038 = ~n5023 & ~n5037 ;
  assign n5039 = ~n2184 & ~n4908 ;
  assign n5040 = ~n4947 & ~n5039 ;
  assign n5041 = ~n4053 & ~n4949 ;
  assign n5042 = ~n2197 & ~n5041 ;
  assign n5043 = n2546 & n2739 ;
  assign n5044 = ~n3251 & ~n5043 ;
  assign n5045 = ~n5042 & n5044 ;
  assign n5046 = n4908 & ~n5045 ;
  assign n5047 = ~n4937 & ~n5046 ;
  assign n5048 = ~n5040 & n5047 ;
  assign n5049 = n2110 & ~n5048 ;
  assign n5050 = ~n5038 & ~n5049 ;
  assign n5051 = ~n5019 & n5050 ;
  assign n5052 = ~n4980 & n5051 ;
  assign n5053 = n1073 & n2218 ;
  assign n5054 = n1583 & n3294 ;
  assign n5055 = n278 & n1254 ;
  assign n5056 = ~n5054 & ~n5055 ;
  assign n5057 = ~n5053 & n5056 ;
  assign n5058 = n42 & ~n5057 ;
  assign n5059 = n291 & n3283 ;
  assign n5060 = x5 & n5059 ;
  assign n5061 = ~n5058 & ~n5060 ;
  assign n5062 = n4954 & ~n5061 ;
  assign n5063 = ~x0 & ~n269 ;
  assign n5064 = n5028 & ~n5063 ;
  assign n5065 = x6 & ~n470 ;
  assign n5066 = n104 & n5065 ;
  assign n5067 = x13 ^ x11 ;
  assign n5068 = n1454 & ~n5067 ;
  assign n5069 = n5068 ^ n5067 ;
  assign n5070 = n5066 & n5069 ;
  assign n5071 = ~n5064 & ~n5070 ;
  assign n5072 = n799 & ~n5071 ;
  assign n5073 = n278 & n1492 ;
  assign n5074 = n2218 ^ n1290 ;
  assign n5075 = ~x0 & ~n5074 ;
  assign n5076 = n5075 ^ n2218 ;
  assign n5077 = ~x4 & ~n5076 ;
  assign n5078 = ~n5073 & ~n5077 ;
  assign n5079 = ~n470 & ~n5078 ;
  assign n5080 = n42 & n5054 ;
  assign n5081 = ~n5079 & ~n5080 ;
  assign n5082 = n5081 ^ n291 ;
  assign n5083 = n5082 ^ n5081 ;
  assign n5084 = n5081 ^ n107 ;
  assign n5085 = n5084 ^ n5081 ;
  assign n5086 = n5083 & n5085 ;
  assign n5087 = n5086 ^ n5081 ;
  assign n5088 = x13 & ~n5087 ;
  assign n5089 = n5088 ^ n5081 ;
  assign n5090 = n571 & ~n5089 ;
  assign n5091 = ~n284 & ~n2233 ;
  assign n5092 = ~n470 & n5091 ;
  assign n5093 = x5 & ~x11 ;
  assign n5094 = n5092 & n5093 ;
  assign n5095 = n3649 & n5094 ;
  assign n5096 = n205 & n5093 ;
  assign n5097 = ~n2234 & n5096 ;
  assign n5098 = n2264 ^ x5 ;
  assign n5099 = n5098 ^ n2264 ;
  assign n5100 = n2264 ^ n320 ;
  assign n5101 = n5100 ^ n2264 ;
  assign n5102 = ~n5099 & ~n5101 ;
  assign n5103 = n5102 ^ n2264 ;
  assign n5104 = x0 & n5103 ;
  assign n5105 = n5104 ^ n2264 ;
  assign n5106 = n4500 & n5105 ;
  assign n5107 = ~n5097 & ~n5106 ;
  assign n5108 = ~n5095 & n5107 ;
  assign n5109 = n1027 & ~n5108 ;
  assign n5110 = ~n5090 & ~n5109 ;
  assign n5111 = ~n5072 & n5110 ;
  assign n5112 = n5111 ^ x7 ;
  assign n5113 = n5112 ^ n5111 ;
  assign n5114 = n5113 ^ n5062 ;
  assign n5115 = n78 & ~n1253 ;
  assign n5116 = ~n1021 & ~n5115 ;
  assign n5117 = n1261 & ~n5116 ;
  assign n5118 = n74 & n1433 ;
  assign n5119 = n104 & n5118 ;
  assign n5120 = ~n5117 & ~n5119 ;
  assign n5121 = n1618 & ~n5120 ;
  assign n5122 = ~x6 & n3296 ;
  assign n5123 = n5093 & n5122 ;
  assign n5124 = ~x5 & ~n1352 ;
  assign n5125 = ~n470 & n1021 ;
  assign n5126 = n5124 & n5125 ;
  assign n5127 = ~n5123 & ~n5126 ;
  assign n5128 = ~n2234 & ~n5127 ;
  assign n5129 = ~n5121 & ~n5128 ;
  assign n5130 = n5129 ^ x1 ;
  assign n5131 = x1 & ~n5130 ;
  assign n5132 = n5131 ^ n5111 ;
  assign n5133 = n5132 ^ x1 ;
  assign n5134 = n5114 & ~n5133 ;
  assign n5135 = n5134 ^ n5131 ;
  assign n5136 = n5135 ^ x1 ;
  assign n5137 = ~n5062 & n5136 ;
  assign n5138 = n5137 ^ n5062 ;
  assign n5139 = n2682 & n5138 ;
  assign n5140 = n222 & n3421 ;
  assign n5141 = n1994 & n5027 ;
  assign n5142 = n5140 & n5141 ;
  assign n5143 = n258 & n2756 ;
  assign n5144 = ~n1352 & n5143 ;
  assign n5145 = n74 & n2106 ;
  assign n5146 = n1261 & n5145 ;
  assign n5147 = ~n5144 & ~n5146 ;
  assign n5148 = ~n470 & ~n5147 ;
  assign n5149 = x15 & n281 ;
  assign n5150 = ~x4 & n1583 ;
  assign n5151 = n354 & n1728 ;
  assign n5152 = n5150 & n5151 ;
  assign n5153 = n5149 & n5152 ;
  assign n5154 = ~x2 & ~n5153 ;
  assign n5155 = ~n5148 & n5154 ;
  assign n5156 = ~x6 & n1456 ;
  assign n5157 = n310 & n5151 ;
  assign n5158 = n5156 & n5157 ;
  assign n5159 = n66 & n74 ;
  assign n5160 = n263 & n5159 ;
  assign n5161 = n394 & n5160 ;
  assign n5162 = ~n5144 & ~n5161 ;
  assign n5163 = ~n43 & ~n5162 ;
  assign n5164 = x2 & ~n5163 ;
  assign n5165 = ~n5158 & n5164 ;
  assign n5166 = ~n5155 & ~n5165 ;
  assign n5167 = ~n5142 & ~n5166 ;
  assign n5168 = x7 & ~n5167 ;
  assign n5169 = n140 & n5151 ;
  assign n5170 = n308 & n2809 ;
  assign n5171 = ~n5169 & ~n5170 ;
  assign n5172 = n256 & ~n5171 ;
  assign n5173 = n247 & n267 ;
  assign n5174 = n207 & n269 ;
  assign n5175 = ~n5173 & ~n5174 ;
  assign n5176 = x15 & n5170 ;
  assign n5177 = ~n5175 & n5176 ;
  assign n5178 = ~n5172 & ~n5177 ;
  assign n5179 = n640 & ~n5178 ;
  assign n5180 = n1253 ^ n909 ;
  assign n5181 = x1 & ~n5180 ;
  assign n5182 = n5181 ^ n909 ;
  assign n5183 = n3317 & n5182 ;
  assign n5184 = ~n20 & ~n394 ;
  assign n5185 = ~n221 & ~n792 ;
  assign n5186 = n5184 & ~n5185 ;
  assign n5187 = n74 & n5186 ;
  assign n5188 = ~n4247 & n5187 ;
  assign n5189 = ~n5183 & ~n5188 ;
  assign n5190 = n66 & n592 ;
  assign n5191 = ~n5189 & n5190 ;
  assign n5192 = ~n5179 & ~n5191 ;
  assign n5193 = ~n5168 & n5192 ;
  assign n5194 = ~n2710 & ~n5193 ;
  assign n5195 = ~n5139 & ~n5194 ;
  assign n5196 = n5052 & n5195 ;
  assign n5197 = n2876 & n4940 ;
  assign n5198 = n3009 & n5197 ;
  assign n5199 = n1599 & n2168 ;
  assign n5200 = n1823 & n5199 ;
  assign n5201 = n3809 & n5200 ;
  assign n5202 = n5201 ^ x4 ;
  assign n5203 = n5202 ^ n5201 ;
  assign n5204 = n5203 ^ n5198 ;
  assign n5205 = n507 & n5182 ;
  assign n5206 = n372 & n2079 ;
  assign n5207 = ~n5205 & ~n5206 ;
  assign n5208 = n1642 & ~n5207 ;
  assign n5209 = n2501 & n5199 ;
  assign n5210 = ~n5208 & ~n5209 ;
  assign n5211 = n5210 ^ x2 ;
  assign n5212 = x2 & ~n5211 ;
  assign n5213 = n5212 ^ n5201 ;
  assign n5214 = n5213 ^ x2 ;
  assign n5215 = n5204 & n5214 ;
  assign n5216 = n5215 ^ n5212 ;
  assign n5217 = n5216 ^ x2 ;
  assign n5218 = ~n5198 & n5217 ;
  assign n5219 = n5218 ^ n5198 ;
  assign n5220 = n165 & n5219 ;
  assign n5221 = n107 & n394 ;
  assign n5222 = x1 & ~n2278 ;
  assign n5223 = n2756 & n5222 ;
  assign n5224 = n2253 & n5199 ;
  assign n5225 = ~n5223 & ~n5224 ;
  assign n5226 = n5221 & ~n5225 ;
  assign n5227 = ~x9 & n1630 ;
  assign n5228 = ~n1253 & n5227 ;
  assign n5229 = n1376 & n1942 ;
  assign n5230 = n5228 & n5229 ;
  assign n5231 = ~n5226 & ~n5230 ;
  assign n5232 = n260 & n2867 ;
  assign n5233 = x5 & ~n4989 ;
  assign n5234 = ~n5055 & ~n5233 ;
  assign n5235 = n1084 & ~n5234 ;
  assign n5236 = x5 & n2868 ;
  assign n5237 = n249 & n318 ;
  assign n5238 = n165 & n5237 ;
  assign n5239 = ~n5236 & ~n5238 ;
  assign n5240 = ~n5235 & n5239 ;
  assign n5241 = ~x11 & ~n5240 ;
  assign n5242 = ~n5232 & ~n5241 ;
  assign n5243 = ~n2865 & ~n5242 ;
  assign n5244 = n5231 & ~n5243 ;
  assign n5245 = ~n5220 & n5244 ;
  assign n5246 = ~n43 & ~n5245 ;
  assign n5247 = n2615 & n2833 ;
  assign n5248 = n2832 ^ n2809 ;
  assign n5249 = n5248 ^ n2832 ;
  assign n5250 = n3264 ^ n2832 ;
  assign n5251 = n5250 ^ n2832 ;
  assign n5252 = n5249 & ~n5251 ;
  assign n5253 = n5252 ^ n2832 ;
  assign n5254 = ~n2282 & n5253 ;
  assign n5255 = n5254 ^ n2832 ;
  assign n5256 = ~x3 & n5255 ;
  assign n5257 = ~n5247 & ~n5256 ;
  assign n5258 = n5122 & ~n5257 ;
  assign n5259 = n425 & n2950 ;
  assign n5260 = n4348 & n5259 ;
  assign n5261 = n2445 & n5260 ;
  assign n5262 = ~n5258 & ~n5261 ;
  assign n5263 = ~n745 & ~n5262 ;
  assign n5264 = ~x9 & n263 ;
  assign n5265 = n1150 & n2041 ;
  assign n5266 = x6 & n5265 ;
  assign n5267 = ~n5264 & ~n5266 ;
  assign n5268 = ~n2197 & ~n5267 ;
  assign n5269 = n1715 & n5268 ;
  assign n5270 = ~x2 & n816 ;
  assign n5271 = n291 & ~n2743 ;
  assign n5272 = ~n1506 & ~n5271 ;
  assign n5273 = n642 & ~n5272 ;
  assign n5274 = x6 & n5227 ;
  assign n5275 = ~n5273 & ~n5274 ;
  assign n5276 = n5270 & ~n5275 ;
  assign n5277 = n228 & n1671 ;
  assign n5278 = ~n1670 & ~n5277 ;
  assign n5279 = x0 & ~n5277 ;
  assign n5280 = ~n5278 & ~n5279 ;
  assign n5281 = n5264 & n5280 ;
  assign n5282 = n3809 & n4573 ;
  assign n5283 = n1123 & n3060 ;
  assign n5284 = n5282 & n5283 ;
  assign n5285 = ~n5281 & ~n5284 ;
  assign n5286 = ~n5276 & n5285 ;
  assign n5287 = n206 & n2739 ;
  assign n5288 = n394 & ~n2743 ;
  assign n5289 = ~n2687 & ~n5288 ;
  assign n5290 = ~n5287 & n5289 ;
  assign n5291 = x2 & ~n5290 ;
  assign n5292 = ~x4 & n4214 ;
  assign n5293 = ~n5291 & ~n5292 ;
  assign n5294 = n875 & ~n5293 ;
  assign n5295 = n1715 & n3161 ;
  assign n5296 = ~x4 & n642 ;
  assign n5297 = ~n1433 & ~n4737 ;
  assign n5298 = ~x14 & n1254 ;
  assign n5299 = ~x9 & n1290 ;
  assign n5300 = ~n5298 & ~n5299 ;
  assign n5301 = ~n5297 & ~n5300 ;
  assign n5302 = ~n5296 & ~n5301 ;
  assign n5303 = n5295 & ~n5302 ;
  assign n5304 = ~n5294 & ~n5303 ;
  assign n5305 = n5286 & n5304 ;
  assign n5306 = ~n5269 & n5305 ;
  assign n5307 = n2786 & ~n5306 ;
  assign n5308 = ~n5263 & ~n5307 ;
  assign n5309 = x15 & ~n5308 ;
  assign n5310 = ~n79 & n3009 ;
  assign n5311 = ~n3295 & ~n3595 ;
  assign n5312 = n5311 ^ n77 ;
  assign n5313 = n5312 ^ n5311 ;
  assign n5314 = ~n1826 & ~n2758 ;
  assign n5315 = n5314 ^ n5311 ;
  assign n5316 = n5315 ^ n5311 ;
  assign n5317 = ~n5313 & ~n5316 ;
  assign n5318 = n5317 ^ n5311 ;
  assign n5319 = ~x2 & n5318 ;
  assign n5320 = n5319 ^ n5311 ;
  assign n5321 = ~n5310 & ~n5320 ;
  assign n5322 = n551 & ~n5321 ;
  assign n5323 = n2257 & n5296 ;
  assign n5324 = ~n5322 & ~n5323 ;
  assign n5325 = n2857 & ~n5324 ;
  assign n5326 = n254 & n1702 ;
  assign n5327 = ~x4 & ~n3982 ;
  assign n5328 = n5326 & ~n5327 ;
  assign n5329 = n1248 & ~n3983 ;
  assign n5330 = n251 & n5329 ;
  assign n5331 = ~n208 & ~n2929 ;
  assign n5332 = ~n5330 & n5331 ;
  assign n5333 = ~n5328 & n5332 ;
  assign n5334 = n551 & ~n5333 ;
  assign n5335 = n287 & n3294 ;
  assign n5336 = ~n431 & n1456 ;
  assign n5337 = ~n5299 & ~n5336 ;
  assign n5338 = n210 & ~n5337 ;
  assign n5339 = ~n5335 & ~n5338 ;
  assign n5340 = ~n5334 & n5339 ;
  assign n5341 = n1608 & ~n5340 ;
  assign n5342 = ~n5325 & ~n5341 ;
  assign n5343 = n571 & ~n5342 ;
  assign n5344 = x5 & ~x8 ;
  assign n5345 = n210 & n394 ;
  assign n5346 = n5344 & n5345 ;
  assign n5347 = n1634 & n3452 ;
  assign n5348 = n1518 & n5174 ;
  assign n5349 = x0 & n5348 ;
  assign n5350 = ~n5347 & ~n5349 ;
  assign n5351 = ~n5346 & n5350 ;
  assign n5352 = n1366 & ~n5351 ;
  assign n5353 = ~x13 & n551 ;
  assign n5354 = n4966 & n5353 ;
  assign n5355 = n1261 & n4573 ;
  assign n5356 = n425 & n4064 ;
  assign n5357 = n5355 & n5356 ;
  assign n5358 = ~n5354 & ~n5357 ;
  assign n5359 = ~n5352 & n5358 ;
  assign n5360 = n5359 ^ x11 ;
  assign n5361 = n5360 ^ n5359 ;
  assign n5362 = n5361 ^ x1 ;
  assign n5363 = n210 & n2776 ;
  assign n5364 = n281 & n5363 ;
  assign n5365 = n1366 & n1667 ;
  assign n5366 = n3220 & n5365 ;
  assign n5367 = n1503 ^ x0 ;
  assign n5368 = n5367 ^ n2168 ;
  assign n5369 = ~n1078 & ~n1433 ;
  assign n5370 = n5369 ^ n394 ;
  assign n5371 = n1503 & n5370 ;
  assign n5372 = n5371 ^ n394 ;
  assign n5373 = ~n5368 & n5372 ;
  assign n5374 = n5373 ^ n5371 ;
  assign n5375 = n5374 ^ n394 ;
  assign n5376 = n5375 ^ n1503 ;
  assign n5377 = n2168 & n5376 ;
  assign n5378 = ~n5366 & ~n5377 ;
  assign n5379 = x2 & ~n5378 ;
  assign n5380 = ~n5364 & ~n5379 ;
  assign n5381 = n5380 ^ x5 ;
  assign n5382 = x5 & ~n5381 ;
  assign n5383 = n5382 ^ n5359 ;
  assign n5384 = n5383 ^ x5 ;
  assign n5385 = n5362 & ~n5384 ;
  assign n5386 = n5385 ^ n5382 ;
  assign n5387 = n5386 ^ x5 ;
  assign n5388 = ~x1 & n5387 ;
  assign n5389 = ~n5343 & ~n5388 ;
  assign n5390 = n63 & ~n5389 ;
  assign n5391 = ~n5309 & ~n5390 ;
  assign n5392 = n1775 & n2639 ;
  assign n5393 = n24 & ~n2865 ;
  assign n5394 = ~n3763 & ~n5393 ;
  assign n5395 = ~n5392 & n5394 ;
  assign n5396 = n1582 & ~n5395 ;
  assign n5397 = n214 & n1669 ;
  assign n5398 = n2253 & n5397 ;
  assign n5399 = n1942 & n3761 ;
  assign n5400 = ~n5398 & ~n5399 ;
  assign n5401 = ~n5396 & n5400 ;
  assign n5402 = n1123 & ~n5401 ;
  assign n5403 = ~x6 & n792 ;
  assign n5404 = ~n2865 & n5403 ;
  assign n5405 = n291 & n3763 ;
  assign n5406 = ~n5404 & ~n5405 ;
  assign n5407 = ~x0 & ~n5406 ;
  assign n5408 = x9 & n394 ;
  assign n5409 = ~x8 & n1941 ;
  assign n5410 = n5408 & n5409 ;
  assign n5411 = ~n5407 & ~n5410 ;
  assign n5412 = n1138 & ~n5411 ;
  assign n5413 = ~x2 & n222 ;
  assign n5414 = ~n284 & n4214 ;
  assign n5415 = n2695 & n5414 ;
  assign n5416 = n214 & n313 ;
  assign n5417 = n1672 & n5416 ;
  assign n5418 = ~n5415 & ~n5417 ;
  assign n5419 = n5413 & ~n5418 ;
  assign n5420 = ~n5412 & ~n5419 ;
  assign n5421 = ~n5402 & n5420 ;
  assign n5422 = ~x11 & ~n5421 ;
  assign n5423 = n909 & n2005 ;
  assign n5424 = n74 & n286 ;
  assign n5425 = ~n5423 & ~n5424 ;
  assign n5426 = n3161 & ~n5425 ;
  assign n5427 = n2038 & n5199 ;
  assign n5428 = ~n5426 & ~n5427 ;
  assign n5429 = x3 & ~n5428 ;
  assign n5430 = ~n5223 & ~n5429 ;
  assign n5431 = n5054 & ~n5430 ;
  assign n5432 = x5 & ~n1352 ;
  assign n5433 = n1857 ^ n507 ;
  assign n5434 = n5433 ^ n5159 ;
  assign n5435 = n5434 ^ n1857 ;
  assign n5436 = n5435 ^ n5434 ;
  assign n5437 = ~n1253 & n2632 ;
  assign n5438 = n5437 ^ n5434 ;
  assign n5439 = n5438 ^ n5433 ;
  assign n5440 = n5436 & ~n5439 ;
  assign n5441 = n5440 ^ n5437 ;
  assign n5442 = ~n909 & ~n5437 ;
  assign n5443 = n5442 ^ n5433 ;
  assign n5444 = ~n5441 & ~n5443 ;
  assign n5445 = n5444 ^ n5442 ;
  assign n5446 = ~n5433 & n5445 ;
  assign n5447 = n5446 ^ n5440 ;
  assign n5448 = n5447 ^ n507 ;
  assign n5449 = n5448 ^ n5437 ;
  assign n5450 = ~x8 & ~n5449 ;
  assign n5451 = n50 & n2782 ;
  assign n5452 = n2075 & n5451 ;
  assign n5453 = ~n5450 & ~n5452 ;
  assign n5454 = n5432 & ~n5453 ;
  assign n5455 = n104 & ~n5207 ;
  assign n5456 = n2724 & n5455 ;
  assign n5457 = ~n5454 & ~n5456 ;
  assign n5458 = ~n5431 & n5457 ;
  assign n5459 = ~n470 & ~n5458 ;
  assign n5460 = ~n5422 & ~n5459 ;
  assign n5461 = n5391 & n5460 ;
  assign n5462 = ~n5246 & n5461 ;
  assign n5463 = n5462 ^ x7 ;
  assign n5464 = n5463 ^ n5462 ;
  assign n5465 = ~n431 & ~n2342 ;
  assign n5466 = n5259 & n5465 ;
  assign n5467 = n4500 & n4737 ;
  assign n5468 = n1138 & n5467 ;
  assign n5469 = ~n5466 & ~n5468 ;
  assign n5470 = n3283 & ~n5469 ;
  assign n5471 = ~x0 & n1123 ;
  assign n5472 = ~n528 & n2105 ;
  assign n5473 = n5471 & n5472 ;
  assign n5474 = ~x11 & n5473 ;
  assign n5475 = ~n5470 & ~n5474 ;
  assign n5476 = n2277 & ~n5475 ;
  assign n5477 = x11 & n294 ;
  assign n5478 = n2256 & n5477 ;
  assign n5479 = n1634 & n5478 ;
  assign n5480 = n2005 & n5479 ;
  assign n5481 = ~n5476 & ~n5480 ;
  assign n5482 = n550 & ~n5481 ;
  assign n5483 = ~n2756 & ~n5159 ;
  assign n5484 = n1073 & n3981 ;
  assign n5485 = ~n3250 & ~n5484 ;
  assign n5486 = n263 & n2405 ;
  assign n5487 = ~n5485 & n5486 ;
  assign n5488 = n1290 & n2558 ;
  assign n5489 = n221 & n1073 ;
  assign n5490 = n5488 & n5489 ;
  assign n5491 = n1630 & n2075 ;
  assign n5492 = n5059 & n5491 ;
  assign n5493 = ~n5490 & ~n5492 ;
  assign n5494 = ~n5487 & n5493 ;
  assign n5495 = ~n5483 & ~n5494 ;
  assign n5496 = n41 & n3649 ;
  assign n5497 = n1609 & n5496 ;
  assign n5505 = ~x3 & n394 ;
  assign n5506 = x11 & n1550 ;
  assign n5507 = n5505 & n5506 ;
  assign n5498 = n2775 & ~n3725 ;
  assign n5499 = ~n1669 & n2786 ;
  assign n5500 = ~n5498 & ~n5499 ;
  assign n5501 = ~x6 & ~n2276 ;
  assign n5502 = ~n228 & ~n5501 ;
  assign n5503 = ~n5500 & n5502 ;
  assign n5504 = ~n117 & n5503 ;
  assign n5508 = n5507 ^ n5504 ;
  assign n5509 = n5508 ^ n5504 ;
  assign n5510 = ~x4 & n2223 ;
  assign n5511 = n74 & n2558 ;
  assign n5512 = n5510 & n5511 ;
  assign n5513 = n5512 ^ n5504 ;
  assign n5514 = n5513 ^ n5504 ;
  assign n5515 = ~n5509 & ~n5514 ;
  assign n5516 = n5515 ^ n5504 ;
  assign n5517 = n210 & ~n5516 ;
  assign n5518 = n5517 ^ n5504 ;
  assign n5519 = ~n5497 & ~n5518 ;
  assign n5520 = n943 & ~n5519 ;
  assign n5521 = ~x8 & n2302 ;
  assign n5522 = n228 & n5477 ;
  assign n5523 = n5521 & n5522 ;
  assign n5524 = n5523 ^ n2786 ;
  assign n5525 = n5524 ^ x0 ;
  assign n5540 = n5525 ^ n5524 ;
  assign n5526 = x2 & n291 ;
  assign n5527 = ~x6 & n2739 ;
  assign n5528 = n228 & n5527 ;
  assign n5529 = ~n5526 & ~n5528 ;
  assign n5530 = ~x0 & ~n5529 ;
  assign n5531 = ~n1669 & ~n5288 ;
  assign n5532 = n210 & ~n5531 ;
  assign n5533 = ~n5530 & ~n5532 ;
  assign n5534 = n5533 ^ n5525 ;
  assign n5535 = n5534 ^ n5524 ;
  assign n5536 = n5525 ^ n5523 ;
  assign n5537 = n5536 ^ n5533 ;
  assign n5538 = n5537 ^ n5535 ;
  assign n5539 = ~n5535 & ~n5538 ;
  assign n5541 = n5540 ^ n5539 ;
  assign n5542 = n5541 ^ n5535 ;
  assign n5543 = ~x6 & ~n2282 ;
  assign n5544 = ~n4052 & n5543 ;
  assign n5545 = ~x4 & n20 ;
  assign n5546 = ~n5271 & ~n5545 ;
  assign n5547 = ~x2 & ~n2739 ;
  assign n5548 = ~n5546 & ~n5547 ;
  assign n5549 = ~n5544 & ~n5548 ;
  assign n5550 = n5549 ^ n5524 ;
  assign n5551 = n5539 ^ n5535 ;
  assign n5552 = n5550 & ~n5551 ;
  assign n5553 = n5552 ^ n5524 ;
  assign n5554 = n5542 & n5553 ;
  assign n5555 = n5554 ^ n5524 ;
  assign n5556 = n5555 ^ n2786 ;
  assign n5557 = n5556 ^ n5524 ;
  assign n5558 = n2041 & n5557 ;
  assign n5559 = x0 & n3725 ;
  assign n5560 = ~n4987 & ~n5559 ;
  assign n5561 = n291 & ~n5560 ;
  assign n5562 = ~n2256 & n2598 ;
  assign n5563 = ~n4052 & n5562 ;
  assign n5564 = ~x0 & n2276 ;
  assign n5565 = x6 & n5564 ;
  assign n5566 = ~n5563 & ~n5565 ;
  assign n5567 = ~n5561 & n5566 ;
  assign n5568 = n74 & n365 ;
  assign n5569 = ~n5567 & n5568 ;
  assign n5570 = ~n5558 & ~n5569 ;
  assign n5571 = ~n5520 & n5570 ;
  assign n5572 = n5571 ^ x5 ;
  assign n5573 = n5572 ^ n5571 ;
  assign n5574 = n450 & n909 ;
  assign n5575 = n77 & n5182 ;
  assign n5576 = ~n5574 & ~n5575 ;
  assign n5577 = n228 & n2272 ;
  assign n5578 = n2105 & n5577 ;
  assign n5579 = ~n5576 & n5578 ;
  assign n5580 = ~n2278 & ~n5311 ;
  assign n5581 = ~n3319 & ~n5580 ;
  assign n5582 = n817 & ~n5581 ;
  assign n5583 = n21 & n3245 ;
  assign n5584 = n528 & n5583 ;
  assign n5585 = ~n5582 & ~n5584 ;
  assign n5586 = n29 & ~n5585 ;
  assign n5587 = n308 & n2079 ;
  assign n5588 = ~n3557 & ~n3789 ;
  assign n5589 = n5588 ^ n252 ;
  assign n5590 = n5589 ^ n5588 ;
  assign n5591 = n5588 ^ n528 ;
  assign n5592 = n5591 ^ n5588 ;
  assign n5593 = n5590 & n5592 ;
  assign n5594 = n5593 ^ n5588 ;
  assign n5595 = ~x2 & ~n5594 ;
  assign n5596 = n5595 ^ n5588 ;
  assign n5597 = n3643 & ~n5596 ;
  assign n5598 = n528 & n1669 ;
  assign n5599 = n5021 & n5598 ;
  assign n5600 = ~n5597 & ~n5599 ;
  assign n5601 = n5587 & ~n5600 ;
  assign n5602 = ~n5586 & ~n5601 ;
  assign n5603 = n2005 & n5574 ;
  assign n5604 = n3701 & n5603 ;
  assign n5605 = n790 & ~n1352 ;
  assign n5606 = n2590 & n5605 ;
  assign n5607 = n24 & n5606 ;
  assign n5608 = ~n5604 & ~n5607 ;
  assign n5609 = n1957 & n5477 ;
  assign n5610 = ~n5159 & ~n5609 ;
  assign n5611 = n2704 & ~n5610 ;
  assign n5612 = x0 & n1786 ;
  assign n5613 = n2809 & n5612 ;
  assign n5614 = n909 & n2119 ;
  assign n5615 = n1715 & n3069 ;
  assign n5616 = n5614 & n5615 ;
  assign n5617 = ~n5613 & ~n5616 ;
  assign n5618 = ~n5200 & n5617 ;
  assign n5619 = n469 & n1611 ;
  assign n5620 = n78 & n5619 ;
  assign n5621 = ~n2006 & n5620 ;
  assign n5622 = n5618 & ~n5621 ;
  assign n5623 = ~n5611 & n5622 ;
  assign n5624 = n2656 & ~n5623 ;
  assign n5625 = n5608 & ~n5624 ;
  assign n5626 = n5602 & n5625 ;
  assign n5627 = ~n5579 & n5626 ;
  assign n5628 = n5627 ^ n5571 ;
  assign n5629 = ~n5573 & n5628 ;
  assign n5630 = n5629 ^ n5571 ;
  assign n5631 = ~n5495 & n5630 ;
  assign n5632 = x15 & ~n5631 ;
  assign n5633 = ~x0 & n1027 ;
  assign n5634 = ~x11 & n1630 ;
  assign n5635 = n5633 & n5634 ;
  assign n5636 = ~x14 & n1027 ;
  assign n5637 = n107 & n1611 ;
  assign n5638 = n5636 & n5637 ;
  assign n5639 = ~n2739 & ~n4691 ;
  assign n5640 = ~x5 & n1073 ;
  assign n5641 = ~n538 & ~n571 ;
  assign n5642 = n5640 & ~n5641 ;
  assign n5643 = ~n5639 & n5642 ;
  assign n5644 = ~n5638 & ~n5643 ;
  assign n5645 = ~n5635 & n5644 ;
  assign n5646 = n1582 & ~n5645 ;
  assign n5647 = ~x5 & ~x8 ;
  assign n5648 = x1 & n259 ;
  assign n5649 = ~n5485 & n5648 ;
  assign n5650 = ~n278 & ~n1073 ;
  assign n5651 = ~n450 & ~n5650 ;
  assign n5652 = x13 & n3249 ;
  assign n5653 = ~n5641 & n5652 ;
  assign n5654 = n5651 & n5653 ;
  assign n5655 = ~n5649 & ~n5654 ;
  assign n5656 = n5647 & ~n5655 ;
  assign n5657 = ~n5646 & ~n5656 ;
  assign n5658 = n286 & ~n5657 ;
  assign n5659 = n2877 & n5096 ;
  assign n5660 = n74 & n3249 ;
  assign n5661 = n5471 & n5660 ;
  assign n5662 = n701 & n909 ;
  assign n5663 = n2867 & n5662 ;
  assign n5664 = ~n5661 & ~n5663 ;
  assign n5665 = ~n5659 & n5664 ;
  assign n5666 = n3417 & ~n5665 ;
  assign n5667 = ~n214 & ~n4573 ;
  assign n5668 = n20 & n1599 ;
  assign n5669 = n258 & n1073 ;
  assign n5670 = n21 & n1456 ;
  assign n5671 = ~n5669 & ~n5670 ;
  assign n5672 = n5668 & ~n5671 ;
  assign n5673 = ~n5667 & n5672 ;
  assign n5674 = ~n5666 & ~n5673 ;
  assign n5675 = ~n5658 & n5674 ;
  assign n5676 = x3 & ~n5675 ;
  assign n5677 = ~x2 & n5182 ;
  assign n5678 = x2 & ~x13 ;
  assign n5679 = n571 & n5678 ;
  assign n5680 = ~n5677 & ~n5679 ;
  assign n5681 = ~x5 & n1642 ;
  assign n5682 = n235 & n5681 ;
  assign n5683 = ~n5680 & n5682 ;
  assign n5684 = n357 & n5683 ;
  assign n5685 = n2075 & n2156 ;
  assign n5686 = n5140 & n5685 ;
  assign n5687 = n2109 & n5124 ;
  assign n5688 = n1397 & n2695 ;
  assign n5689 = ~n5687 & ~n5688 ;
  assign n5690 = ~n2278 & ~n5689 ;
  assign n5691 = ~n5686 & ~n5690 ;
  assign n5692 = n1021 & ~n5691 ;
  assign n5693 = ~n2415 & ~n3161 ;
  assign n5694 = n295 & n5496 ;
  assign n5695 = n2809 & n5694 ;
  assign n5696 = ~n5693 & n5695 ;
  assign n5697 = ~n5692 & ~n5696 ;
  assign n5698 = ~n5684 & n5697 ;
  assign n5699 = ~n470 & ~n5698 ;
  assign n5700 = ~n5676 & ~n5699 ;
  assign n5701 = ~n5632 & n5700 ;
  assign n5702 = ~n5482 & n5701 ;
  assign n5703 = n5702 ^ n5462 ;
  assign n5704 = ~n5464 & n5703 ;
  assign n5705 = n5704 ^ n5462 ;
  assign n5706 = n5196 & n5705 ;
  assign n5707 = n2677 & ~n5706 ;
  assign n5708 = ~n4840 & ~n5707 ;
  assign n5709 = n2534 & n5708 ;
  assign n5793 = n1255 & ~n1702 ;
  assign n5794 = ~n85 & ~n2119 ;
  assign n5795 = n5793 & ~n5794 ;
  assign n5796 = n5150 ^ n3462 ;
  assign n5797 = n5796 ^ n5150 ;
  assign n5798 = n5150 ^ n222 ;
  assign n5799 = n5798 ^ n5150 ;
  assign n5800 = ~n5797 & n5799 ;
  assign n5801 = n5800 ^ n5150 ;
  assign n5802 = x2 & n5801 ;
  assign n5803 = n5802 ^ n5150 ;
  assign n5804 = n2272 & n5803 ;
  assign n5805 = n5804 ^ x7 ;
  assign n5806 = n5805 ^ n5804 ;
  assign n5807 = n5806 ^ n5795 ;
  assign n5808 = n2302 & n5413 ;
  assign n5809 = n2218 & n2582 ;
  assign n5810 = ~n104 & n5809 ;
  assign n5811 = n1261 ^ x6 ;
  assign n5812 = n5811 ^ n1261 ;
  assign n5813 = n1985 & ~n5812 ;
  assign n5814 = n5813 ^ n1261 ;
  assign n5815 = ~n2127 & n5814 ;
  assign n5816 = n1702 & n5815 ;
  assign n5714 = n31 & n1290 ;
  assign n5817 = ~x6 & n41 ;
  assign n5818 = ~x5 & n5817 ;
  assign n5819 = ~n5714 & ~n5818 ;
  assign n5820 = n210 & ~n5819 ;
  assign n5821 = ~n5816 & ~n5820 ;
  assign n5822 = x14 & ~n5821 ;
  assign n5823 = ~n5810 & ~n5822 ;
  assign n5824 = ~n5808 & n5823 ;
  assign n5825 = n5824 ^ x8 ;
  assign n5826 = ~n5824 & n5825 ;
  assign n5827 = n5826 ^ n5804 ;
  assign n5828 = n5827 ^ n5824 ;
  assign n5829 = n5807 & ~n5828 ;
  assign n5830 = n5829 ^ n5826 ;
  assign n5831 = n5830 ^ n5824 ;
  assign n5832 = ~n5795 & ~n5831 ;
  assign n5833 = n5832 ^ n5795 ;
  assign n5710 = n3991 & n4251 ;
  assign n5711 = n2587 & ~n2602 ;
  assign n5712 = ~n5710 & ~n5711 ;
  assign n5713 = n1518 & ~n5712 ;
  assign n5715 = ~n2586 & n2704 ;
  assign n5716 = n5714 & n5715 ;
  assign n5717 = ~n3297 & ~n4124 ;
  assign n5718 = x2 & n5647 ;
  assign n5719 = ~n5717 & n5718 ;
  assign n5720 = ~n861 & n5719 ;
  assign n5721 = ~n5716 & ~n5720 ;
  assign n5722 = ~n5713 & n5721 ;
  assign n5723 = n257 & ~n5722 ;
  assign n5724 = n2503 & n4995 ;
  assign n5725 = n217 & n5724 ;
  assign n5726 = n210 & n235 ;
  assign n5727 = n22 & n2442 ;
  assign n5728 = n5726 & n5727 ;
  assign n5729 = ~n5725 & ~n5728 ;
  assign n5730 = ~n5723 & n5729 ;
  assign n5834 = n5833 ^ n5730 ;
  assign n5731 = n107 & n2599 ;
  assign n5732 = n466 & n5731 ;
  assign n5741 = ~n3803 & n5640 ;
  assign n5742 = n3294 & n5488 ;
  assign n5743 = ~n1630 & ~n5527 ;
  assign n5744 = n278 & ~n5743 ;
  assign n5745 = ~n1492 & n5744 ;
  assign n5746 = ~n5742 & ~n5745 ;
  assign n5747 = ~n5741 & n5746 ;
  assign n5748 = n1786 & ~n5747 ;
  assign n5749 = n1926 & n2289 ;
  assign n5750 = ~n3249 & n5749 ;
  assign n5751 = n2223 & n4052 ;
  assign n5752 = n132 & n5751 ;
  assign n5753 = ~n5750 & ~n5752 ;
  assign n5754 = n165 & ~n2309 ;
  assign n5755 = n249 & n5754 ;
  assign n5756 = ~n104 & n267 ;
  assign n5757 = n1581 & n5756 ;
  assign n5758 = n5647 ^ n1630 ;
  assign n5759 = n5758 ^ n394 ;
  assign n5760 = n1630 ^ x14 ;
  assign n5761 = n1630 ^ x0 ;
  assign n5762 = n5761 ^ n5760 ;
  assign n5763 = ~n5760 & n5762 ;
  assign n5764 = n5763 ^ n1630 ;
  assign n5765 = n5764 ^ n5760 ;
  assign n5766 = n5759 & ~n5765 ;
  assign n5767 = n5766 ^ n5763 ;
  assign n5768 = n5767 ^ n5760 ;
  assign n5769 = n394 & ~n5768 ;
  assign n5770 = ~n5757 & ~n5769 ;
  assign n5771 = ~n5755 & n5770 ;
  assign n5772 = n1823 & ~n5771 ;
  assign n5773 = n100 & n2277 ;
  assign n5774 = n3649 ^ n1433 ;
  assign n5775 = n5774 ^ n1433 ;
  assign n5776 = n5369 ^ n1433 ;
  assign n5777 = n5775 & n5776 ;
  assign n5778 = n5777 ^ n1433 ;
  assign n5779 = n5773 & n5778 ;
  assign n5780 = ~n5772 & ~n5779 ;
  assign n5781 = n5753 & n5780 ;
  assign n5782 = ~n5748 & n5781 ;
  assign n5733 = ~n210 & n394 ;
  assign n5734 = n2558 & n5733 ;
  assign n5735 = ~n3728 & ~n5173 ;
  assign n5736 = n2709 & ~n5735 ;
  assign n5737 = ~n268 & ~n394 ;
  assign n5738 = n3643 & ~n5737 ;
  assign n5739 = ~n5736 & ~n5738 ;
  assign n5740 = ~n5734 & n5739 ;
  assign n5783 = n5782 ^ n5740 ;
  assign n5784 = n5783 ^ n5782 ;
  assign n5785 = n5782 ^ n129 ;
  assign n5786 = n5785 ^ n5782 ;
  assign n5787 = ~n5784 & n5786 ;
  assign n5788 = n5787 ^ n5782 ;
  assign n5789 = ~x7 & ~n5788 ;
  assign n5790 = n5789 ^ n5782 ;
  assign n5791 = ~n5732 & n5790 ;
  assign n5792 = n5791 ^ n5730 ;
  assign n5835 = n5834 ^ n5792 ;
  assign n5836 = n5792 ^ x9 ;
  assign n5837 = n5836 ^ n5792 ;
  assign n5838 = ~n5835 & n5837 ;
  assign n5839 = n5838 ^ n5792 ;
  assign n5840 = ~x13 & n5839 ;
  assign n5841 = n5840 ^ n5730 ;
  assign n5842 = x1 & ~n5841 ;
  assign n5843 = n25 & n1902 ;
  assign n5844 = ~x14 & n5843 ;
  assign n5845 = n4218 & n5844 ;
  assign n5846 = n294 & n5471 ;
  assign n5847 = n1101 & n5846 ;
  assign n5848 = ~n5845 & ~n5847 ;
  assign n5849 = ~x2 & ~n5848 ;
  assign n5850 = n22 & n214 ;
  assign n5851 = ~n5843 & ~n5850 ;
  assign n5852 = n41 & n210 ;
  assign n5853 = n927 & n5852 ;
  assign n5854 = ~n5851 & n5853 ;
  assign n5855 = n3759 & n5844 ;
  assign n5856 = ~n5854 & ~n5855 ;
  assign n5857 = ~n5849 & n5856 ;
  assign n5858 = ~n2289 & ~n5857 ;
  assign n5859 = ~n5842 & ~n5858 ;
  assign n5860 = n1256 & ~n5859 ;
  assign n5861 = n1395 & n3728 ;
  assign n5862 = ~n292 & ~n3314 ;
  assign n5863 = n277 & n5862 ;
  assign n5864 = n2857 & n5863 ;
  assign n5865 = ~n5861 & ~n5864 ;
  assign n5866 = n41 & n101 ;
  assign n5867 = ~n5865 & n5866 ;
  assign n5868 = n1246 & ~n1546 ;
  assign n5869 = n206 & n5868 ;
  assign n5870 = n1602 & n3421 ;
  assign n5871 = n3821 & n5870 ;
  assign n5872 = ~n5869 & ~n5871 ;
  assign n5873 = n1366 & ~n5872 ;
  assign n5874 = ~n2387 & ~n3314 ;
  assign n5875 = n5122 & n5874 ;
  assign n5876 = ~n830 & n5875 ;
  assign n5877 = n1457 & n4348 ;
  assign n5878 = ~n5876 & ~n5877 ;
  assign n5879 = n5878 ^ x8 ;
  assign n5880 = n5879 ^ n5878 ;
  assign n5881 = n5880 ^ n603 ;
  assign n5882 = n85 & n394 ;
  assign n5883 = n5678 ^ n603 ;
  assign n5884 = n5882 & ~n5883 ;
  assign n5885 = n5884 ^ n5878 ;
  assign n5886 = ~n5881 & ~n5885 ;
  assign n5887 = n5886 ^ n5884 ;
  assign n5888 = ~n603 & n5887 ;
  assign n5889 = n5888 ^ n5884 ;
  assign n5890 = n5889 ^ n5886 ;
  assign n5891 = ~n5873 & ~n5890 ;
  assign n5892 = ~n5867 & n5891 ;
  assign n5893 = n1779 & ~n5892 ;
  assign n5894 = x10 ^ x7 ;
  assign n5895 = n49 & n2445 ;
  assign n5896 = n1608 & n3068 ;
  assign n5897 = ~n5895 & ~n5896 ;
  assign n5898 = n206 & n1829 ;
  assign n5899 = n1340 & n4251 ;
  assign n5902 = n5899 ^ n5862 ;
  assign n5903 = n5902 ^ n5899 ;
  assign n5900 = n5899 ^ n466 ;
  assign n5901 = n5900 ^ n5899 ;
  assign n5904 = n5903 ^ n5901 ;
  assign n5905 = n5899 ^ n3296 ;
  assign n5906 = n5905 ^ n5899 ;
  assign n5907 = n5906 ^ n5903 ;
  assign n5908 = ~n5903 & ~n5907 ;
  assign n5909 = n5908 ^ n5903 ;
  assign n5910 = ~n5904 & ~n5909 ;
  assign n5911 = n5910 ^ n5908 ;
  assign n5912 = n5911 ^ n5899 ;
  assign n5913 = n5912 ^ n5903 ;
  assign n5914 = ~x6 & ~n5913 ;
  assign n5915 = n5914 ^ n5899 ;
  assign n5916 = ~n5898 & ~n5915 ;
  assign n5917 = ~n5897 & ~n5916 ;
  assign n5918 = n206 & n284 ;
  assign n5919 = ~n1252 & ~n2156 ;
  assign n5920 = n1786 & ~n5919 ;
  assign n5921 = ~n2863 & ~n5920 ;
  assign n5922 = n5918 & ~n5921 ;
  assign n5923 = n2006 & ~n3728 ;
  assign n5924 = n117 & n294 ;
  assign n5925 = n4052 & n5924 ;
  assign n5926 = n5923 & n5925 ;
  assign n5927 = n2586 & n2679 ;
  assign n5928 = ~x3 & n286 ;
  assign n5929 = ~n5927 & ~n5928 ;
  assign n5930 = ~x13 & n5122 ;
  assign n5931 = ~n5929 & n5930 ;
  assign n5932 = ~n5926 & ~n5931 ;
  assign n5933 = ~n5922 & n5932 ;
  assign n5934 = n587 & ~n5933 ;
  assign n5935 = ~x8 & n1702 ;
  assign n5936 = n1276 & n4608 ;
  assign n5937 = n5935 & n5936 ;
  assign n5938 = n1366 & n5937 ;
  assign n5939 = ~n5934 & ~n5938 ;
  assign n5940 = n210 & n291 ;
  assign n5941 = ~n2458 & ~n2678 ;
  assign n5942 = n3808 & ~n5941 ;
  assign n5943 = n5940 & n5942 ;
  assign n5944 = n5939 & ~n5943 ;
  assign n5945 = ~n5917 & n5944 ;
  assign n5946 = n5945 ^ n5894 ;
  assign n5947 = n5946 ^ x10 ;
  assign n5948 = n5947 ^ n5946 ;
  assign n5949 = ~x8 & n3967 ;
  assign n5950 = n86 & n117 ;
  assign n5951 = n1484 & n5950 ;
  assign n5952 = n1433 & n2555 ;
  assign n5953 = ~n830 & n5952 ;
  assign n5954 = x12 & n5953 ;
  assign n5955 = ~n5951 & ~n5954 ;
  assign n5956 = n5949 & ~n5955 ;
  assign n5957 = n639 & n5545 ;
  assign n5958 = n1365 & n5957 ;
  assign n5959 = n210 & n1581 ;
  assign n5960 = n425 & n5959 ;
  assign n5961 = n394 & n1702 ;
  assign n5962 = ~n1550 & n5961 ;
  assign n5963 = ~n5960 & ~n5962 ;
  assign n5964 = n890 & ~n5963 ;
  assign n5965 = n294 & n1394 ;
  assign n5966 = n5940 & n5965 ;
  assign n5967 = ~n5964 & ~n5966 ;
  assign n5968 = ~n5958 & n5967 ;
  assign n5969 = x3 & ~n5968 ;
  assign n5970 = ~x2 & n5951 ;
  assign n5971 = ~n5969 & ~n5970 ;
  assign n5972 = n1991 & ~n5971 ;
  assign n5973 = ~x13 & n1433 ;
  assign n5974 = n2277 & n5973 ;
  assign n5975 = n2555 & n5974 ;
  assign n5976 = n5940 ^ n2309 ;
  assign n5977 = x13 ^ x8 ;
  assign n5978 = n5977 ^ x13 ;
  assign n5979 = n609 ^ x13 ;
  assign n5980 = n5978 & n5979 ;
  assign n5981 = n5980 ^ x13 ;
  assign n5982 = n5981 ^ n5940 ;
  assign n5983 = ~n5976 & ~n5982 ;
  assign n5984 = n5983 ^ n5980 ;
  assign n5985 = n5984 ^ x13 ;
  assign n5986 = n5985 ^ n2309 ;
  assign n5987 = n5940 & n5986 ;
  assign n5988 = n5987 ^ n5940 ;
  assign n5989 = ~n5975 & ~n5988 ;
  assign n5990 = n1256 & ~n5989 ;
  assign n5991 = n66 & n5990 ;
  assign n5992 = ~x12 & n2277 ;
  assign n5993 = n5918 & n5992 ;
  assign n5994 = ~x8 & n38 ;
  assign n5995 = n206 & n5994 ;
  assign n5996 = ~n2857 & n5122 ;
  assign n5997 = n1529 & n5996 ;
  assign n5998 = ~n5995 & ~n5997 ;
  assign n5999 = n3264 & ~n5998 ;
  assign n6000 = ~x8 & ~n529 ;
  assign n6001 = ~n1608 & n5940 ;
  assign n6002 = ~n6000 & n6001 ;
  assign n6003 = ~n5999 & ~n6002 ;
  assign n6004 = ~n5993 & n6003 ;
  assign n6005 = n1859 & ~n6004 ;
  assign n6006 = ~n5991 & ~n6005 ;
  assign n6007 = ~n5972 & n6006 ;
  assign n6008 = ~n5956 & n6007 ;
  assign n6009 = n6008 ^ n5946 ;
  assign n6010 = n6009 ^ n5894 ;
  assign n6011 = ~n5948 & ~n6010 ;
  assign n6012 = n6011 ^ n6008 ;
  assign n6013 = ~n3069 & ~n4573 ;
  assign n6014 = n1528 & ~n6013 ;
  assign n6015 = n6014 ^ x9 ;
  assign n6016 = n6015 ^ n6014 ;
  assign n6017 = n6014 ^ n1394 ;
  assign n6018 = n6017 ^ n6014 ;
  assign n6019 = n6016 & ~n6018 ;
  assign n6020 = n6019 ^ n6014 ;
  assign n6021 = ~x3 & n6020 ;
  assign n6022 = n6021 ^ n6014 ;
  assign n6023 = n5122 & n6022 ;
  assign n6024 = ~x4 & ~n3069 ;
  assign n6025 = n117 & ~n570 ;
  assign n6026 = ~n2126 & n6025 ;
  assign n6027 = n6024 & n6026 ;
  assign n6028 = ~n1528 & n6027 ;
  assign n6029 = ~n6023 & ~n6028 ;
  assign n6030 = n4312 & ~n6029 ;
  assign n6031 = n2857 & n5882 ;
  assign n6032 = ~n1642 & n3294 ;
  assign n6033 = ~n1582 & n6032 ;
  assign n6034 = ~n830 & n6033 ;
  assign n6035 = ~n6031 & ~n6034 ;
  assign n6036 = n86 & n2548 ;
  assign n6037 = ~n6035 & n6036 ;
  assign n6038 = ~x0 & n3249 ;
  assign n6039 = n395 & n3277 ;
  assign n6040 = ~n6038 & ~n6039 ;
  assign n6041 = ~x14 & ~n31 ;
  assign n6042 = n286 & n2857 ;
  assign n6043 = ~n6041 & n6042 ;
  assign n6044 = ~n6040 & n6043 ;
  assign n6045 = n2556 & n5973 ;
  assign n6046 = n1059 & n4941 ;
  assign n6047 = ~n6045 & ~n6046 ;
  assign n6048 = ~n457 & ~n6047 ;
  assign n6049 = ~n6044 & ~n6048 ;
  assign n6050 = ~n6037 & n6049 ;
  assign n6051 = ~n6030 & n6050 ;
  assign n6052 = n6008 & n6051 ;
  assign n6053 = n6052 ^ n5894 ;
  assign n6054 = n6012 & ~n6053 ;
  assign n6055 = n6054 ^ n6052 ;
  assign n6056 = ~n5894 & n6055 ;
  assign n6057 = n6056 ^ n6011 ;
  assign n6058 = n6057 ^ x7 ;
  assign n6059 = n6058 ^ n6008 ;
  assign n6060 = ~n5893 & n6059 ;
  assign n6061 = ~n745 & ~n6060 ;
  assign n6062 = ~x4 & n2351 ;
  assign n6063 = n86 & n6062 ;
  assign n6064 = n2253 & n6063 ;
  assign n6065 = n394 & n550 ;
  assign n6066 = n3260 & n6065 ;
  assign n6067 = ~x1 & n3296 ;
  assign n6068 = ~n3049 & ~n3509 ;
  assign n6069 = n6067 & ~n6068 ;
  assign n6070 = n221 & n4132 ;
  assign n6071 = ~n6069 & ~n6070 ;
  assign n6072 = n3421 & ~n6071 ;
  assign n6073 = ~n6066 & ~n6072 ;
  assign n6074 = ~n6064 & n6073 ;
  assign n6075 = n22 & ~n6074 ;
  assign n6076 = ~n1276 & ~n2351 ;
  assign n6077 = ~n148 & ~n6076 ;
  assign n6078 = ~x14 & n731 ;
  assign n6079 = n3017 & n6078 ;
  assign n6080 = n6077 & n6079 ;
  assign n6081 = n1340 & n1917 ;
  assign n6082 = n403 & n1266 ;
  assign n6083 = n6081 & n6082 ;
  assign n6084 = ~n6080 & ~n6083 ;
  assign n6085 = ~n6075 & n6084 ;
  assign n6086 = n1366 & ~n6085 ;
  assign n6087 = x0 & n185 ;
  assign n6088 = n1902 & n6087 ;
  assign n6089 = n5815 & n6088 ;
  assign n6090 = n3049 & n6089 ;
  assign n6091 = n861 & n1267 ;
  assign n6092 = ~x5 & n294 ;
  assign n6093 = n1438 & n6092 ;
  assign n6094 = n3203 & n6093 ;
  assign n6095 = n6091 & n6094 ;
  assign n6096 = ~n6090 & ~n6095 ;
  assign n6097 = ~n6086 & n6096 ;
  assign n6098 = ~x8 & ~n6097 ;
  assign n6099 = ~x3 & n24 ;
  assign n6100 = ~n248 & n6099 ;
  assign n6101 = n49 & n674 ;
  assign n6102 = n1267 & n1518 ;
  assign n6103 = n6101 & n6102 ;
  assign n6104 = n6100 & n6103 ;
  assign n6105 = ~n691 & n3217 ;
  assign n6106 = n3044 & n6105 ;
  assign n6107 = ~n6104 & ~n6106 ;
  assign n6108 = ~n6098 & n6107 ;
  assign n6109 = ~n6061 & n6108 ;
  assign n6110 = ~n1493 & ~n2857 ;
  assign n6111 = n2075 ^ n1267 ;
  assign n6112 = n21 & n31 ;
  assign n6113 = x2 & n6112 ;
  assign n6114 = n6113 ^ n6111 ;
  assign n6115 = n6114 ^ n1267 ;
  assign n6116 = n6115 ^ n6114 ;
  assign n6117 = n235 & n1312 ;
  assign n6118 = ~n5936 & ~n6117 ;
  assign n6119 = ~x0 & ~n6118 ;
  assign n6120 = n6119 ^ n6114 ;
  assign n6121 = n6120 ^ n6111 ;
  assign n6122 = n6116 & ~n6121 ;
  assign n6123 = n6122 ^ n6119 ;
  assign n6124 = ~x4 & n85 ;
  assign n6125 = ~n6119 & ~n6124 ;
  assign n6126 = n6125 ^ n6111 ;
  assign n6127 = ~n6123 & ~n6126 ;
  assign n6128 = n6127 ^ n6125 ;
  assign n6129 = ~n6111 & n6128 ;
  assign n6130 = n6129 ^ n6122 ;
  assign n6131 = n6130 ^ n2075 ;
  assign n6132 = n6131 ^ n6119 ;
  assign n6133 = ~n6110 & ~n6132 ;
  assign n6134 = ~n5667 & n6133 ;
  assign n6135 = n189 & n425 ;
  assign n6136 = ~x7 & n2906 ;
  assign n6137 = n284 & n6136 ;
  assign n6138 = ~n6135 & ~n6137 ;
  assign n6139 = ~x4 & n2156 ;
  assign n6140 = n4251 & n6139 ;
  assign n6141 = ~n6138 & n6140 ;
  assign n6142 = ~n6134 & ~n6141 ;
  assign n6143 = ~x5 & ~n6142 ;
  assign n6144 = n280 & n1276 ;
  assign n6145 = n2659 & n6144 ;
  assign n6146 = n354 & ~n528 ;
  assign n6147 = n6145 & n6146 ;
  assign n6148 = ~n1538 & n6147 ;
  assign n6149 = ~n6143 & ~n6148 ;
  assign n6223 = n1273 & n1715 ;
  assign n6224 = n2886 & n6223 ;
  assign n6225 = n258 & n6224 ;
  assign n6152 = ~n1667 & ~n2857 ;
  assign n6153 = n2105 & n6152 ;
  assign n6226 = n684 & n6153 ;
  assign n6227 = n2038 & n6226 ;
  assign n6228 = n674 & ~n1084 ;
  assign n6229 = n1702 & n6228 ;
  assign n6230 = ~n5693 & n6229 ;
  assign n6231 = ~x2 & ~n609 ;
  assign n6232 = ~n2642 & n6231 ;
  assign n6233 = ~n6230 & ~n6232 ;
  assign n6234 = n2308 & ~n6233 ;
  assign n6235 = ~n6227 & ~n6234 ;
  assign n6236 = ~n6225 & n6235 ;
  assign n6189 = n2386 & n2871 ;
  assign n6190 = n129 & n6189 ;
  assign n6191 = n354 & n2500 ;
  assign n6192 = n199 & ~n5919 ;
  assign n6193 = ~n6191 & ~n6192 ;
  assign n6194 = n1266 & ~n2857 ;
  assign n6195 = ~n6193 & n6194 ;
  assign n6196 = ~n6190 & ~n6195 ;
  assign n6197 = n2352 & ~n6196 ;
  assign n6168 = n294 & n2075 ;
  assign n6198 = x8 & n2038 ;
  assign n6199 = ~n284 & n6198 ;
  assign n6200 = ~n6168 & ~n6199 ;
  assign n6201 = n85 & ~n6200 ;
  assign n6202 = n2038 & n5924 ;
  assign n6203 = ~n6201 & ~n6202 ;
  assign n6204 = n1254 & n1482 ;
  assign n6205 = ~n6203 & n6204 ;
  assign n6206 = ~n6197 & ~n6205 ;
  assign n6207 = n2698 & n5227 ;
  assign n6208 = n231 & n2641 ;
  assign n6209 = ~n6207 & ~n6208 ;
  assign n6210 = ~n609 & ~n6209 ;
  assign n6211 = n77 & n934 ;
  assign n6212 = n1138 & n6211 ;
  assign n6213 = ~n6210 & ~n6212 ;
  assign n6214 = ~x7 & ~n6213 ;
  assign n6215 = n768 & n2640 ;
  assign n6216 = ~x5 & n397 ;
  assign n6217 = n6215 & n6216 ;
  assign n6218 = ~n457 & n6217 ;
  assign n6219 = ~n6214 & ~n6218 ;
  assign n6220 = n20 & ~n6219 ;
  assign n6221 = n6206 & ~n6220 ;
  assign n6237 = n6236 ^ n6221 ;
  assign n6164 = ~x6 & ~n609 ;
  assign n6165 = n22 & n1252 ;
  assign n6166 = n2038 & n6165 ;
  assign n6167 = n6164 & n6166 ;
  assign n6169 = ~n1020 & ~n1482 ;
  assign n6170 = n2328 & n6169 ;
  assign n6171 = ~n642 & n6170 ;
  assign n6172 = ~n6165 & ~n6171 ;
  assign n6173 = n6168 & ~n6172 ;
  assign n6174 = n1945 & n2886 ;
  assign n6175 = ~n4376 & n6174 ;
  assign n6176 = n2181 & n4114 ;
  assign n6177 = n4982 & n6176 ;
  assign n6178 = ~n6175 & ~n6177 ;
  assign n6179 = ~n6173 & n6178 ;
  assign n6180 = ~n6167 & n6179 ;
  assign n6150 = n1273 & n2075 ;
  assign n6151 = n4609 & n6150 ;
  assign n6154 = n189 & n6153 ;
  assign n6155 = ~x6 & n927 ;
  assign n6156 = n1482 & ~n1550 ;
  assign n6157 = n6155 & n6156 ;
  assign n6158 = n1493 & n2906 ;
  assign n6159 = n264 & n6158 ;
  assign n6160 = ~n6157 & ~n6159 ;
  assign n6161 = ~n6154 & n6160 ;
  assign n6162 = x2 & ~n6161 ;
  assign n6163 = ~n6151 & ~n6162 ;
  assign n6181 = n6180 ^ n6163 ;
  assign n6182 = n6181 ^ n6180 ;
  assign n6183 = n6180 ^ x5 ;
  assign n6184 = n6183 ^ n6180 ;
  assign n6185 = ~n6182 & n6184 ;
  assign n6186 = n6185 ^ n6180 ;
  assign n6187 = x0 & ~n6186 ;
  assign n6188 = n6187 ^ n6180 ;
  assign n6222 = n6221 ^ n6188 ;
  assign n6238 = n6237 ^ n6222 ;
  assign n6239 = n6222 ^ x3 ;
  assign n6240 = n6239 ^ n6222 ;
  assign n6241 = n6238 & n6240 ;
  assign n6242 = n6241 ^ n6222 ;
  assign n6243 = x4 & n6242 ;
  assign n6244 = n6243 ^ n6221 ;
  assign n6245 = n6244 ^ x12 ;
  assign n6246 = n6245 ^ n6244 ;
  assign n6247 = n6246 ^ n6149 ;
  assign n6248 = ~x8 & n1267 ;
  assign n6249 = n222 & n6248 ;
  assign n6250 = n50 & n6249 ;
  assign n6251 = n222 & n6223 ;
  assign n6252 = n2678 & n6251 ;
  assign n6253 = n280 & n338 ;
  assign n6254 = ~n249 & ~n1669 ;
  assign n6255 = n6253 & n6254 ;
  assign n6256 = ~n1503 & ~n2276 ;
  assign n6257 = n522 & n1261 ;
  assign n6258 = ~n6256 & n6257 ;
  assign n6259 = ~n6255 & ~n6258 ;
  assign n6260 = ~x0 & ~n6259 ;
  assign n6261 = ~n6252 & ~n6260 ;
  assign n6262 = ~n6250 & n6261 ;
  assign n6263 = n2168 & ~n6262 ;
  assign n6264 = n2397 & n2687 ;
  assign n6265 = n1073 & n3264 ;
  assign n6266 = ~n1671 & n6265 ;
  assign n6267 = n3249 & n5959 ;
  assign n6268 = ~n6266 & ~n6267 ;
  assign n6269 = ~n6264 & n6268 ;
  assign n6272 = n6269 ^ n5184 ;
  assign n6273 = n6272 ^ n6269 ;
  assign n6270 = n6269 ^ n2558 ;
  assign n6271 = n6270 ^ n6269 ;
  assign n6274 = n6273 ^ n6271 ;
  assign n6275 = n6269 ^ x0 ;
  assign n6276 = n6275 ^ n6269 ;
  assign n6277 = n6276 ^ n6273 ;
  assign n6278 = ~n6273 & n6277 ;
  assign n6279 = n6278 ^ n6273 ;
  assign n6280 = ~n6274 & ~n6279 ;
  assign n6281 = n6280 ^ n6278 ;
  assign n6282 = n6281 ^ n6269 ;
  assign n6283 = n6282 ^ n6273 ;
  assign n6284 = ~x7 & n6283 ;
  assign n6285 = n6284 ^ n6269 ;
  assign n6286 = n230 & ~n6285 ;
  assign n6287 = ~n1507 & ~n2752 ;
  assign n6288 = ~n3462 & ~n6287 ;
  assign n6289 = n78 & ~n5278 ;
  assign n6290 = ~n6288 & ~n6289 ;
  assign n6291 = n1111 & ~n6290 ;
  assign n6292 = n640 & n1715 ;
  assign n6293 = n1670 & n6292 ;
  assign n6294 = n2304 & ~n3314 ;
  assign n6295 = n5221 & n6294 ;
  assign n6296 = ~n6293 & ~n6295 ;
  assign n6297 = n6296 ^ x3 ;
  assign n6298 = n6297 ^ n6296 ;
  assign n6299 = n6298 ^ n6291 ;
  assign n6300 = n408 & ~n2197 ;
  assign n6301 = n2352 & n6300 ;
  assign n6302 = ~n2138 & ~n2386 ;
  assign n6303 = n1877 & ~n6302 ;
  assign n6304 = ~x7 & n2558 ;
  assign n6305 = ~n1340 & ~n6304 ;
  assign n6306 = n1702 & ~n2309 ;
  assign n6307 = ~n6305 & n6306 ;
  assign n6308 = ~n6303 & ~n6307 ;
  assign n6309 = ~x6 & ~n6308 ;
  assign n6310 = ~n6301 & ~n6309 ;
  assign n6311 = n6310 ^ x5 ;
  assign n6312 = x5 & ~n6311 ;
  assign n6313 = n6312 ^ n6296 ;
  assign n6314 = n6313 ^ x5 ;
  assign n6315 = n6299 & ~n6314 ;
  assign n6316 = n6315 ^ n6312 ;
  assign n6317 = n6316 ^ x5 ;
  assign n6318 = ~n6291 & n6317 ;
  assign n6319 = n6318 ^ n6291 ;
  assign n6320 = ~n6286 & ~n6319 ;
  assign n6321 = n214 & ~n6320 ;
  assign n6322 = n210 & n4272 ;
  assign n6323 = n2549 & n3701 ;
  assign n6324 = ~n247 & n3328 ;
  assign n6325 = ~n2687 & ~n6324 ;
  assign n6326 = n2678 & ~n6325 ;
  assign n6327 = ~n6323 & ~n6326 ;
  assign n6328 = ~n6322 & n6327 ;
  assign n6331 = n6328 ^ n2368 ;
  assign n6332 = n6331 ^ n6328 ;
  assign n6329 = n6328 ^ x3 ;
  assign n6330 = n6329 ^ n6328 ;
  assign n6333 = n6332 ^ n6330 ;
  assign n6334 = n6328 ^ x4 ;
  assign n6335 = n6334 ^ n6328 ;
  assign n6336 = n6335 ^ n6332 ;
  assign n6337 = n6332 & ~n6336 ;
  assign n6338 = n6337 ^ n6332 ;
  assign n6339 = ~n6333 & n6338 ;
  assign n6340 = n6339 ^ n6337 ;
  assign n6341 = n6340 ^ n6328 ;
  assign n6342 = n6341 ^ n6332 ;
  assign n6343 = x13 & ~n6342 ;
  assign n6344 = n6343 ^ n6328 ;
  assign n6345 = n52 & ~n6344 ;
  assign n6346 = ~n6321 & ~n6345 ;
  assign n6347 = ~n6263 & n6346 ;
  assign n6348 = n6347 ^ x1 ;
  assign n6349 = ~n6347 & n6348 ;
  assign n6350 = n6349 ^ n6244 ;
  assign n6351 = n6350 ^ n6347 ;
  assign n6352 = n6247 & n6351 ;
  assign n6353 = n6352 ^ n6349 ;
  assign n6354 = n6353 ^ n6347 ;
  assign n6355 = n6149 & ~n6354 ;
  assign n6356 = n6355 ^ n6149 ;
  assign n6357 = x10 & ~n6356 ;
  assign n6358 = ~x5 & n214 ;
  assign n6359 = ~n5353 & ~n6358 ;
  assign n6360 = ~x14 & n4052 ;
  assign n6361 = n2218 & n6360 ;
  assign n6362 = ~x5 & n267 ;
  assign n6363 = n214 & n1506 ;
  assign n6364 = n6362 & n6363 ;
  assign n6365 = ~n6361 & ~n6364 ;
  assign n6366 = ~n2677 & ~n6365 ;
  assign n6367 = ~n6359 & n6366 ;
  assign n6368 = ~x10 & n281 ;
  assign n6369 = ~n4325 & ~n6368 ;
  assign n6370 = n1598 & ~n4801 ;
  assign n6371 = ~n6369 & n6370 ;
  assign n6372 = ~n1366 & ~n1706 ;
  assign n6373 = n1365 & ~n1760 ;
  assign n6374 = ~n281 & n6373 ;
  assign n6375 = ~n6372 & n6374 ;
  assign n6376 = ~n6371 & ~n6375 ;
  assign n6377 = n6376 ^ n1303 ;
  assign n6378 = n6377 ^ n6376 ;
  assign n6379 = n6376 ^ n2156 ;
  assign n6380 = n6379 ^ n6376 ;
  assign n6381 = n6378 & n6380 ;
  assign n6382 = n6381 ^ n6376 ;
  assign n6383 = ~x6 & ~n6382 ;
  assign n6384 = n6383 ^ n6376 ;
  assign n6385 = n1261 & ~n6384 ;
  assign n6386 = n2699 ^ x10 ;
  assign n6387 = n6386 ^ n2699 ;
  assign n6388 = n269 & ~n1370 ;
  assign n6389 = n6388 ^ n2699 ;
  assign n6390 = n6387 & n6389 ;
  assign n6391 = n6390 ^ n2699 ;
  assign n6392 = n1456 & n6391 ;
  assign n6393 = ~n6385 & ~n6392 ;
  assign n6394 = ~n6367 & n6393 ;
  assign n6395 = n199 & ~n6394 ;
  assign n6396 = ~n1706 & ~n1708 ;
  assign n6397 = n1420 & n1642 ;
  assign n6398 = ~n3954 & ~n6397 ;
  assign n6399 = n6396 & ~n6398 ;
  assign n6400 = n25 & n6399 ;
  assign n6401 = n18 & n86 ;
  assign n6402 = n6401 ^ n640 ;
  assign n6403 = n6402 ^ n5150 ;
  assign n6404 = n6403 ^ n6401 ;
  assign n6405 = n6404 ^ n6403 ;
  assign n6406 = n1257 & n1669 ;
  assign n6407 = n6406 ^ n6403 ;
  assign n6408 = n6407 ^ n6402 ;
  assign n6409 = n6405 & ~n6408 ;
  assign n6410 = n6409 ^ n6406 ;
  assign n6411 = ~n394 & ~n6406 ;
  assign n6412 = n6411 ^ n6402 ;
  assign n6413 = ~n6410 & ~n6412 ;
  assign n6414 = n6413 ^ n6411 ;
  assign n6415 = ~n6402 & n6414 ;
  assign n6416 = n6415 ^ n6409 ;
  assign n6417 = n6416 ^ n640 ;
  assign n6418 = n6417 ^ n6406 ;
  assign n6419 = ~n86 & n1671 ;
  assign n6420 = n2677 & n6419 ;
  assign n6421 = ~x10 & n1642 ;
  assign n6422 = ~n3267 & ~n6421 ;
  assign n6423 = ~n6420 & n6422 ;
  assign n6424 = n1456 & ~n6423 ;
  assign n6425 = n6424 ^ x5 ;
  assign n6426 = n6425 ^ n6424 ;
  assign n6427 = n1257 & n1581 ;
  assign n6428 = ~x14 & n1528 ;
  assign n6429 = ~n1772 & ~n2977 ;
  assign n6430 = ~n394 & ~n6429 ;
  assign n6431 = n6428 & ~n6430 ;
  assign n6432 = ~n6427 & ~n6431 ;
  assign n6433 = n6432 ^ n6424 ;
  assign n6434 = n6433 ^ n6424 ;
  assign n6435 = ~n6426 & ~n6434 ;
  assign n6436 = n6435 ^ n6424 ;
  assign n6437 = ~x7 & n6436 ;
  assign n6438 = n6437 ^ n6424 ;
  assign n6439 = n6418 & ~n6438 ;
  assign n6440 = ~n6400 & n6439 ;
  assign n6441 = n1714 & ~n6440 ;
  assign n6442 = x10 & ~n1394 ;
  assign n6443 = ~n3851 & ~n6442 ;
  assign n6444 = n1714 & ~n6443 ;
  assign n6445 = n1902 & n3174 ;
  assign n6446 = x14 & n6445 ;
  assign n6447 = x14 & n354 ;
  assign n6448 = n1256 & n1366 ;
  assign n6449 = ~x13 & n1404 ;
  assign n6450 = ~n1551 & n6449 ;
  assign n6451 = ~n6448 & ~n6450 ;
  assign n6452 = n6447 & ~n6451 ;
  assign n6453 = ~n6446 & ~n6452 ;
  assign n6454 = ~n6444 & n6453 ;
  assign n6455 = n1990 & ~n6454 ;
  assign n6456 = ~n1257 & ~n3217 ;
  assign n6457 = ~n2289 & n6429 ;
  assign n6458 = ~n6456 & n6457 ;
  assign n6459 = ~n1672 & ~n6429 ;
  assign n6460 = n1438 ^ n1234 ;
  assign n6461 = ~x14 & n6460 ;
  assign n6462 = n6461 ^ n1234 ;
  assign n6463 = n6459 & n6462 ;
  assign n6464 = ~n1352 & ~n1624 ;
  assign n6465 = ~n6463 & ~n6464 ;
  assign n6466 = ~n6458 & n6465 ;
  assign n6467 = n308 & ~n6466 ;
  assign n6468 = n5843 & n6467 ;
  assign n6469 = ~n6455 & ~n6468 ;
  assign n6470 = ~n6441 & n6469 ;
  assign n6471 = ~n1619 & ~n2225 ;
  assign n6472 = ~n222 & n6471 ;
  assign n6473 = n294 & ~n5344 ;
  assign n6474 = ~n6472 & n6473 ;
  assign n6475 = ~n1502 & n6474 ;
  assign n6476 = ~x4 & n1597 ;
  assign n6477 = n1608 & n6476 ;
  assign n6478 = n6477 ^ x14 ;
  assign n6479 = n6478 ^ n6477 ;
  assign n6480 = n6479 ^ n6475 ;
  assign n6481 = n1597 & n2877 ;
  assign n6482 = n6481 ^ x8 ;
  assign n6483 = n6481 & n6482 ;
  assign n6484 = n6483 ^ n6477 ;
  assign n6485 = n6484 ^ n6481 ;
  assign n6486 = ~n6480 & n6485 ;
  assign n6487 = n6486 ^ n6483 ;
  assign n6488 = n6487 ^ n6481 ;
  assign n6489 = ~n6475 & n6488 ;
  assign n6490 = n6489 ^ n6475 ;
  assign n6491 = n1298 & n6490 ;
  assign n6492 = ~n62 & ~n2331 ;
  assign n6493 = n1619 & ~n6492 ;
  assign n6494 = n609 & n6493 ;
  assign n6495 = n17 & ~n5369 ;
  assign n6496 = ~n891 & n6495 ;
  assign n6497 = ~n6494 & ~n6496 ;
  assign n6498 = n1290 & ~n6497 ;
  assign n6499 = n1671 & n2331 ;
  assign n6500 = ~n528 & n6499 ;
  assign n6501 = x5 & n6500 ;
  assign n6502 = ~n5369 & n6501 ;
  assign n6503 = ~n6498 & ~n6502 ;
  assign n6504 = ~n6491 & n6503 ;
  assign n6505 = n264 & ~n6504 ;
  assign n6506 = n1256 & n4052 ;
  assign n6507 = ~n3982 & ~n6506 ;
  assign n6508 = ~n2183 & n6507 ;
  assign n6509 = ~n4247 & ~n4756 ;
  assign n6510 = x5 & ~n6509 ;
  assign n6511 = ~n6508 & n6510 ;
  assign n6512 = ~n1256 & n3234 ;
  assign n6513 = n1456 & n6512 ;
  assign n6514 = ~n6511 & ~n6513 ;
  assign n6515 = n2168 & ~n6514 ;
  assign n6516 = x7 & n6515 ;
  assign n6517 = ~n6505 & ~n6516 ;
  assign n6518 = n354 & ~n6517 ;
  assign n6519 = n6470 & ~n6518 ;
  assign n6520 = ~n6395 & n6519 ;
  assign n6521 = ~n1716 & ~n6520 ;
  assign n6526 = ~n609 & n6165 ;
  assign n6522 = n253 & n1231 ;
  assign n6523 = n1482 & n6522 ;
  assign n6527 = n6526 ^ n6523 ;
  assign n6528 = n6527 ^ n6523 ;
  assign n6524 = n6523 ^ x4 ;
  assign n6525 = n6524 ^ n6523 ;
  assign n6529 = n6528 ^ n6525 ;
  assign n6530 = n6523 ^ n403 ;
  assign n6531 = n6530 ^ n6523 ;
  assign n6532 = n6531 ^ n6528 ;
  assign n6533 = n6528 & ~n6532 ;
  assign n6534 = n6533 ^ n6528 ;
  assign n6535 = n6529 & n6534 ;
  assign n6536 = n6535 ^ n6533 ;
  assign n6537 = n6536 ^ n6523 ;
  assign n6538 = n6537 ^ n6528 ;
  assign n6539 = ~n1582 & n6538 ;
  assign n6540 = n6539 ^ n6523 ;
  assign n6541 = n119 & n5465 ;
  assign n6542 = n1310 & n5296 ;
  assign n6543 = x9 & n1521 ;
  assign n6544 = ~n6542 & ~n6543 ;
  assign n6545 = ~n6541 & n6544 ;
  assign n6546 = n1267 & ~n6545 ;
  assign n6547 = x13 & n3497 ;
  assign n6548 = ~n1656 & ~n6547 ;
  assign n6549 = n222 & ~n6548 ;
  assign n6550 = n133 & n1123 ;
  assign n6551 = n4247 & n6550 ;
  assign n6552 = ~n6549 & ~n6551 ;
  assign n6553 = n264 & ~n6552 ;
  assign n6554 = ~x12 & n264 ;
  assign n6555 = ~n609 & n6554 ;
  assign n6556 = n121 & n674 ;
  assign n6557 = ~n6555 & ~n6556 ;
  assign n6558 = n5156 & ~n6557 ;
  assign n6559 = ~n6553 & ~n6558 ;
  assign n6560 = ~n6546 & n6559 ;
  assign n6561 = n6560 ^ x8 ;
  assign n6562 = n6561 ^ n6560 ;
  assign n6563 = n6562 ^ n6540 ;
  assign n6564 = x7 & ~x13 ;
  assign n6565 = n1433 & n2219 ;
  assign n6566 = ~n5299 & ~n6565 ;
  assign n6567 = n6564 & ~n6566 ;
  assign n6568 = ~n119 & ~n1078 ;
  assign n6569 = n257 & n1254 ;
  assign n6570 = ~n6568 & n6569 ;
  assign n6571 = ~n6567 & ~n6570 ;
  assign n6572 = n6571 ^ x12 ;
  assign n6573 = ~n6571 & ~n6572 ;
  assign n6574 = n6573 ^ n6560 ;
  assign n6575 = n6574 ^ n6571 ;
  assign n6576 = n6563 & n6575 ;
  assign n6577 = n6576 ^ n6573 ;
  assign n6578 = n6577 ^ n6571 ;
  assign n6579 = ~n6540 & ~n6578 ;
  assign n6580 = n6579 ^ n6540 ;
  assign n6581 = n2271 & n6580 ;
  assign n6582 = n1298 & n2309 ;
  assign n6583 = n62 & n1669 ;
  assign n6584 = ~n6582 & ~n6583 ;
  assign n6585 = n1886 & ~n6584 ;
  assign n6586 = n3453 & n4922 ;
  assign n6587 = ~n6585 & ~n6586 ;
  assign n6588 = x9 & ~n6587 ;
  assign n6589 = n264 & n5488 ;
  assign n6590 = ~n49 & n6589 ;
  assign n6591 = ~n6588 & ~n6590 ;
  assign n6592 = n228 & ~n6591 ;
  assign n6593 = n4569 ^ n890 ;
  assign n6594 = n6593 ^ x9 ;
  assign n6595 = n6594 ^ n6593 ;
  assign n6596 = n6595 ^ x5 ;
  assign n6597 = n4569 ^ x14 ;
  assign n6598 = ~x14 & ~n6597 ;
  assign n6599 = n6598 ^ n6593 ;
  assign n6600 = n6599 ^ x14 ;
  assign n6601 = ~n6596 & ~n6600 ;
  assign n6602 = n6601 ^ n6598 ;
  assign n6603 = n6602 ^ x14 ;
  assign n6604 = ~x5 & ~n6603 ;
  assign n6605 = n6604 ^ n4569 ;
  assign n6606 = n6564 & n6605 ;
  assign n6607 = n1310 & n2174 ;
  assign n6608 = ~n6606 & ~n6607 ;
  assign n6609 = n1503 & ~n6608 ;
  assign n6610 = n2308 & n4451 ;
  assign n6611 = x5 & n425 ;
  assign n6612 = n399 & n603 ;
  assign n6613 = ~n6554 & ~n6612 ;
  assign n6614 = n6611 & ~n6613 ;
  assign n6615 = ~n891 & n6569 ;
  assign n6616 = ~n257 & ~n264 ;
  assign n6617 = n267 & n1231 ;
  assign n6618 = ~n6616 & n6617 ;
  assign n6619 = ~n6615 & ~n6618 ;
  assign n6620 = ~n6614 & n6619 ;
  assign n6621 = n6620 ^ x8 ;
  assign n6622 = n6621 ^ n6620 ;
  assign n6623 = n6622 ^ n6610 ;
  assign n6624 = n52 & n1177 ;
  assign n6625 = ~n5850 & ~n6624 ;
  assign n6626 = n6625 ^ x6 ;
  assign n6627 = ~n6625 & n6626 ;
  assign n6628 = n6627 ^ n6620 ;
  assign n6629 = n6628 ^ n6625 ;
  assign n6630 = n6623 & n6629 ;
  assign n6631 = n6630 ^ n6627 ;
  assign n6632 = n6631 ^ n6625 ;
  assign n6633 = ~n6610 & ~n6632 ;
  assign n6634 = n6633 ^ n6610 ;
  assign n6635 = ~n6609 & ~n6634 ;
  assign n6636 = n247 & ~n6635 ;
  assign n6637 = ~n6592 & ~n6636 ;
  assign n6638 = n1732 & ~n6637 ;
  assign n6639 = ~n2699 & ~n2729 ;
  assign n6640 = n4022 & ~n6639 ;
  assign n6641 = n2387 & n3553 ;
  assign n6642 = n2126 & n6641 ;
  assign n6643 = ~n6640 & ~n6642 ;
  assign n6644 = n1230 & ~n6643 ;
  assign n6645 = n780 & n5363 ;
  assign n6646 = n1273 & n2445 ;
  assign n6647 = ~x4 & n1702 ;
  assign n6648 = n3453 & n6647 ;
  assign n6649 = n6646 & n6648 ;
  assign n6650 = ~n6645 & ~n6649 ;
  assign n6651 = ~n6644 & n6650 ;
  assign n6652 = ~x5 & ~n6651 ;
  assign n6653 = ~n6638 & ~n6652 ;
  assign n6654 = ~n6581 & n6653 ;
  assign n6655 = n355 & ~n6654 ;
  assign n6656 = n1623 ^ n1257 ;
  assign n6657 = n6656 ^ n1623 ;
  assign n6658 = n1623 ^ x8 ;
  assign n6659 = n6658 ^ n1623 ;
  assign n6660 = n6657 & n6659 ;
  assign n6661 = n6660 ^ n1623 ;
  assign n6662 = ~x5 & n6661 ;
  assign n6663 = n6662 ^ n1623 ;
  assign n6664 = n3728 & n6663 ;
  assign n6665 = n17 & n3048 ;
  assign n6666 = n6362 & n6665 ;
  assign n6667 = ~n6664 & ~n6666 ;
  assign n6668 = n450 & ~n6667 ;
  assign n6669 = ~x6 & n1801 ;
  assign n6670 = x1 & x10 ;
  assign n6671 = n4117 & n6670 ;
  assign n6672 = n6669 & n6671 ;
  assign n6673 = n1492 & n3267 ;
  assign n6674 = ~x2 & n1583 ;
  assign n6675 = n6401 & n6674 ;
  assign n6676 = ~n6673 & ~n6675 ;
  assign n6677 = n24 & ~n6676 ;
  assign n6678 = n2276 & n3196 ;
  assign n6679 = n1254 & n6678 ;
  assign n6680 = n503 & n1562 ;
  assign n6681 = n6674 & n6680 ;
  assign n6682 = n18 & n3282 ;
  assign n6683 = ~n1266 & n6682 ;
  assign n6684 = ~x6 & n6683 ;
  assign n6685 = ~n6681 & ~n6684 ;
  assign n6686 = ~n6679 & n6685 ;
  assign n6687 = n21 & ~n6686 ;
  assign n6688 = ~n6677 & ~n6687 ;
  assign n6689 = ~n6672 & n6688 ;
  assign n6690 = ~n6668 & n6689 ;
  assign n6691 = n41 & ~n6690 ;
  assign n6692 = n1917 & n6401 ;
  assign n6693 = n1256 & n4691 ;
  assign n6694 = ~x0 & n2592 ;
  assign n6695 = ~n3277 & ~n6694 ;
  assign n6696 = ~n1757 & n6695 ;
  assign n6697 = n6693 & ~n6696 ;
  assign n6698 = ~n6692 & ~n6697 ;
  assign n6699 = n1634 & ~n6698 ;
  assign n6700 = n1625 & n1715 ;
  assign n6701 = n78 & n6682 ;
  assign n6702 = n17 & n3049 ;
  assign n6703 = ~n3261 & ~n6702 ;
  assign n6704 = ~n6701 & n6703 ;
  assign n6705 = ~n6700 & n6704 ;
  assign n6706 = n2280 & ~n6705 ;
  assign n6707 = n1261 & n6706 ;
  assign n6708 = ~x1 & n280 ;
  assign n6709 = n3267 & n6708 ;
  assign n6710 = n1583 & n2038 ;
  assign n6711 = n6401 & n6710 ;
  assign n6712 = ~n6709 & ~n6711 ;
  assign n6713 = ~x0 & ~n6712 ;
  assign n6714 = x1 & n3981 ;
  assign n6715 = n295 & ~n3643 ;
  assign n6716 = ~n1624 & n6715 ;
  assign n6717 = n6714 & n6716 ;
  assign n6718 = ~n6713 & ~n6717 ;
  assign n6719 = n4608 & ~n6718 ;
  assign n6720 = ~x7 & ~n6719 ;
  assign n6721 = ~x6 & n2282 ;
  assign n6722 = n3154 & n6721 ;
  assign n6723 = n2319 & n6722 ;
  assign n6724 = ~x4 & n6723 ;
  assign n6725 = n6720 & ~n6724 ;
  assign n6726 = ~n6707 & n6725 ;
  assign n6727 = ~n6699 & n6726 ;
  assign n6728 = ~n6691 & n6727 ;
  assign n6729 = n24 & n2309 ;
  assign n6730 = ~n984 & n2704 ;
  assign n6731 = ~n6729 & ~n6730 ;
  assign n6732 = n4774 & ~n6731 ;
  assign n6733 = n1123 & n6732 ;
  assign n6734 = n1256 & n1518 ;
  assign n6735 = n50 & n792 ;
  assign n6736 = n6734 & n6735 ;
  assign n6737 = x12 & ~n2309 ;
  assign n6738 = x10 & n6737 ;
  assign n6739 = ~n926 & ~n2640 ;
  assign n6740 = n6738 & n6739 ;
  assign n6741 = n223 & n6740 ;
  assign n6742 = ~n6736 & ~n6741 ;
  assign n6745 = n6671 ^ n132 ;
  assign n6746 = n6745 ^ n6671 ;
  assign n6743 = n6671 ^ n18 ;
  assign n6744 = n6743 ^ n6671 ;
  assign n6747 = n6746 ^ n6744 ;
  assign n6748 = n6671 ^ n533 ;
  assign n6749 = n6748 ^ n6671 ;
  assign n6750 = n6749 ^ n6746 ;
  assign n6751 = ~n6746 & ~n6750 ;
  assign n6752 = n6751 ^ n6746 ;
  assign n6753 = ~n6747 & ~n6752 ;
  assign n6754 = n6753 ^ n6751 ;
  assign n6755 = n6754 ^ n6671 ;
  assign n6756 = n6755 ^ n6746 ;
  assign n6757 = ~n165 & ~n6756 ;
  assign n6758 = n6757 ^ n6671 ;
  assign n6759 = n4608 & n6758 ;
  assign n6760 = n6742 & ~n6759 ;
  assign n6761 = ~n6733 & n6760 ;
  assign n6762 = n2598 & ~n6761 ;
  assign n6763 = n1625 ^ x4 ;
  assign n6764 = n6763 ^ n1625 ;
  assign n6765 = n6738 ^ n1625 ;
  assign n6766 = ~n6764 & n6765 ;
  assign n6767 = n6766 ^ n1625 ;
  assign n6768 = ~n1943 & n6767 ;
  assign n6769 = ~n1483 & ~n1620 ;
  assign n6770 = n6769 ^ n1716 ;
  assign n6771 = n6770 ^ n6769 ;
  assign n6772 = ~x12 & ~n1733 ;
  assign n6773 = ~n3569 & ~n6772 ;
  assign n6774 = n1506 & n6773 ;
  assign n6775 = n6774 ^ n6769 ;
  assign n6776 = n6771 & ~n6775 ;
  assign n6777 = n6776 ^ n6769 ;
  assign n6778 = n6447 & ~n6777 ;
  assign n6779 = ~n6768 & ~n6778 ;
  assign n6780 = n1290 & ~n6779 ;
  assign n6781 = x1 & n1623 ;
  assign n6782 = n1757 & n6781 ;
  assign n6783 = n3708 & n4117 ;
  assign n6784 = n24 & n6783 ;
  assign n6785 = ~n6782 & ~n6784 ;
  assign n6786 = n5150 & ~n6785 ;
  assign n6787 = ~x4 & n2038 ;
  assign n6788 = ~x3 & n6787 ;
  assign n6789 = ~n2974 & ~n6788 ;
  assign n6790 = n1583 & ~n6789 ;
  assign n6791 = n3267 & n6790 ;
  assign n6792 = x7 & ~n6791 ;
  assign n6793 = ~n6786 & n6792 ;
  assign n6794 = n6708 ^ n2555 ;
  assign n6795 = x4 & n3217 ;
  assign n6796 = n6795 ^ n2272 ;
  assign n6797 = n6796 ^ n6795 ;
  assign n6798 = ~n224 & n2558 ;
  assign n6799 = n1256 & ~n4052 ;
  assign n6800 = ~n6041 & n6799 ;
  assign n6801 = ~n6798 & n6800 ;
  assign n6802 = n6801 ^ n6795 ;
  assign n6803 = ~n6797 & n6802 ;
  assign n6804 = n6803 ^ n6795 ;
  assign n6805 = n6804 ^ n6708 ;
  assign n6806 = n6794 & n6805 ;
  assign n6807 = n6806 ^ n6803 ;
  assign n6808 = n6807 ^ n6795 ;
  assign n6809 = n6808 ^ n2555 ;
  assign n6810 = n6708 & n6809 ;
  assign n6811 = n6810 ^ n6708 ;
  assign n6812 = n6793 & ~n6811 ;
  assign n6813 = ~x8 & n890 ;
  assign n6814 = n1073 & n2257 ;
  assign n6815 = n6813 & n6814 ;
  assign n6816 = n1332 & n6815 ;
  assign n6817 = x12 ^ x10 ;
  assign n6818 = n3364 ^ x12 ;
  assign n6819 = n6818 ^ n3364 ;
  assign n6820 = n3365 & n6819 ;
  assign n6821 = n6820 ^ n3364 ;
  assign n6822 = ~n6817 & n6821 ;
  assign n6823 = n1376 & n6822 ;
  assign n6824 = n1503 & n1551 ;
  assign n6825 = n4869 & n6824 ;
  assign n6826 = n1483 & n2546 ;
  assign n6827 = ~n6825 & ~n6826 ;
  assign n6828 = ~n6823 & n6827 ;
  assign n6829 = n3864 ^ n1702 ;
  assign n6830 = n6829 ^ n3864 ;
  assign n6831 = n3864 ^ n1257 ;
  assign n6832 = n6831 ^ n3864 ;
  assign n6833 = n6830 & n6832 ;
  assign n6834 = n6833 ^ n3864 ;
  assign n6835 = ~x4 & n6834 ;
  assign n6836 = n6835 ^ n3864 ;
  assign n6837 = n2289 & n6836 ;
  assign n6838 = n6828 & ~n6837 ;
  assign n6839 = n6838 ^ x5 ;
  assign n6840 = n6839 ^ n6838 ;
  assign n6841 = n3439 & n5345 ;
  assign n6842 = n6841 ^ n6838 ;
  assign n6843 = ~n6840 & ~n6842 ;
  assign n6844 = n6843 ^ n6838 ;
  assign n6845 = ~n6816 & n6844 ;
  assign n6846 = ~n558 & ~n6845 ;
  assign n6847 = n6812 & ~n6846 ;
  assign n6848 = ~n6780 & n6847 ;
  assign n6849 = ~n6762 & n6848 ;
  assign n6850 = ~n6728 & ~n6849 ;
  assign n6851 = ~n2169 & n6850 ;
  assign n6852 = ~n6655 & ~n6851 ;
  assign n6853 = ~n6521 & n6852 ;
  assign n6854 = ~n6357 & n6853 ;
  assign n6855 = n6109 & n6854 ;
  assign n6856 = ~n5860 & n6855 ;
  assign n6857 = n6856 ^ x10 ;
  assign n6858 = n5598 & n6647 ;
  assign n6859 = ~n4505 & ~n5678 ;
  assign n6860 = n278 & n3234 ;
  assign n6861 = ~n6859 & n6860 ;
  assign n6862 = ~n6858 & ~n6861 ;
  assign n6863 = n2123 & ~n6862 ;
  assign n6864 = n799 & n1814 ;
  assign n6865 = n1669 & n6864 ;
  assign n6866 = ~x8 & n1312 ;
  assign n6867 = x4 & n450 ;
  assign n6868 = n6866 & n6867 ;
  assign n6869 = n185 & ~n252 ;
  assign n6870 = ~n266 & n6869 ;
  assign n6871 = ~n6150 & ~n6870 ;
  assign n6872 = n2256 & ~n6871 ;
  assign n6873 = ~n6868 & ~n6872 ;
  assign n6874 = ~n6865 & n6873 ;
  assign n6875 = n62 & ~n6874 ;
  assign n6876 = n72 & ~n6302 ;
  assign n6877 = ~n1814 & ~n2257 ;
  assign n6878 = n792 & n6877 ;
  assign n6879 = n6876 & n6878 ;
  assign n6880 = ~n2687 & ~n5059 ;
  assign n6881 = n591 & n3740 ;
  assign n6882 = ~n6880 & n6881 ;
  assign n6883 = ~n6879 & ~n6882 ;
  assign n6884 = ~n6875 & n6883 ;
  assign n6885 = x13 & ~n6884 ;
  assign n6886 = ~n6863 & ~n6885 ;
  assign n6887 = n230 & ~n6886 ;
  assign n6888 = n550 & n6045 ;
  assign n6889 = x3 & n1702 ;
  assign n6890 = n1484 & n2640 ;
  assign n6891 = n284 & n1365 ;
  assign n6892 = n5403 & n6891 ;
  assign n6893 = ~n6890 & ~n6892 ;
  assign n6894 = n6889 & ~n6893 ;
  assign n6895 = n2038 & n5510 ;
  assign n6896 = ~x0 & ~n253 ;
  assign n6897 = n5011 & ~n6896 ;
  assign n6898 = n3462 & n6897 ;
  assign n6899 = ~n6895 & ~n6898 ;
  assign n6900 = n1498 & ~n6899 ;
  assign n6901 = ~n6894 & ~n6900 ;
  assign n6902 = ~n6888 & n6901 ;
  assign n6903 = ~x0 & n404 ;
  assign n6904 = ~n87 & ~n250 ;
  assign n6905 = n3649 & n6904 ;
  assign n6906 = ~n6903 & ~n6905 ;
  assign n6907 = ~n6062 & n6906 ;
  assign n6908 = n4312 & ~n6907 ;
  assign n6912 = ~n120 & ~n1420 ;
  assign n6909 = n61 & n394 ;
  assign n6910 = n503 & n6909 ;
  assign n6911 = ~n5918 & ~n6910 ;
  assign n6913 = n6912 ^ n6911 ;
  assign n6914 = n6913 ^ n6911 ;
  assign n6915 = n6911 ^ n6038 ;
  assign n6916 = n6915 ^ n6911 ;
  assign n6917 = ~n6914 & n6916 ;
  assign n6918 = n6917 ^ n6911 ;
  assign n6919 = ~x2 & ~n6918 ;
  assign n6920 = n6919 ^ n6911 ;
  assign n6921 = ~n6908 & n6920 ;
  assign n6922 = n550 & ~n6921 ;
  assign n6923 = ~x6 & n49 ;
  assign n6924 = ~x14 & n4185 ;
  assign n6925 = ~n6923 & ~n6924 ;
  assign n6926 = x1 & ~n6925 ;
  assign n6927 = n717 & n2424 ;
  assign n6928 = ~n6926 & ~n6927 ;
  assign n6929 = n278 & ~n6928 ;
  assign n6930 = x6 & n529 ;
  assign n6931 = ~x4 & n6930 ;
  assign n6932 = ~n1299 & ~n6931 ;
  assign n6933 = n24 & ~n6932 ;
  assign n6934 = ~n6929 & ~n6933 ;
  assign n6935 = n1786 & ~n6934 ;
  assign n6936 = ~n6922 & ~n6935 ;
  assign n6937 = n6936 ^ x8 ;
  assign n6938 = n6937 ^ n6936 ;
  assign n6939 = n1715 & n6462 ;
  assign n6940 = n394 & n3049 ;
  assign n6941 = ~n6939 & ~n6940 ;
  assign n6942 = n3797 & ~n6941 ;
  assign n6943 = n6942 ^ n6936 ;
  assign n6944 = n6938 & ~n6943 ;
  assign n6945 = n6944 ^ n6936 ;
  assign n6946 = n6902 & n6945 ;
  assign n6947 = n640 & ~n6946 ;
  assign n6948 = ~n6887 & ~n6947 ;
  assign n6949 = n354 & n2304 ;
  assign n6950 = n308 & n2186 ;
  assign n6951 = ~n6949 & ~n6950 ;
  assign n6952 = n4869 & ~n6951 ;
  assign n6953 = n1299 & n6952 ;
  assign n6954 = n1669 & n4348 ;
  assign n6955 = ~n2289 & n6889 ;
  assign n6956 = ~n6954 & ~n6955 ;
  assign n6957 = ~x14 & ~n6956 ;
  assign n6958 = ~x6 & n1702 ;
  assign n6959 = n2678 & n6958 ;
  assign n6960 = ~n6957 & ~n6959 ;
  assign n6961 = n2660 & ~n6960 ;
  assign n6962 = ~n1669 & ~n6360 ;
  assign n6963 = ~n1943 & ~n6962 ;
  assign n6964 = ~n6961 & ~n6963 ;
  assign n6965 = n153 & ~n6964 ;
  assign n6966 = ~x14 & n1438 ;
  assign n6967 = n6966 ^ x6 ;
  assign n6968 = n6967 ^ n6966 ;
  assign n6969 = n6966 ^ n1234 ;
  assign n6970 = n6969 ^ n6966 ;
  assign n6971 = n6968 & ~n6970 ;
  assign n6972 = n6971 ^ n6966 ;
  assign n6973 = x2 & n6972 ;
  assign n6974 = n6973 ^ n6966 ;
  assign n6975 = n6099 & n6974 ;
  assign n6976 = n503 & n2914 ;
  assign n6977 = ~n6975 & ~n6976 ;
  assign n6978 = n1550 & ~n6977 ;
  assign n6979 = ~n251 & n6099 ;
  assign n6980 = ~x2 & n6112 ;
  assign n6981 = ~n6979 & ~n6980 ;
  assign n6982 = n2124 & ~n6981 ;
  assign n6983 = ~n4047 & n6982 ;
  assign n6984 = ~n6978 & ~n6983 ;
  assign n6985 = ~n2368 & ~n3043 ;
  assign n6986 = n753 & ~n6985 ;
  assign n6987 = n244 & n5678 ;
  assign n6988 = ~n5369 & n6987 ;
  assign n6989 = n247 & n3283 ;
  assign n6990 = n49 & n6989 ;
  assign n6991 = ~x0 & n4505 ;
  assign n6992 = ~n6568 & n6991 ;
  assign n6993 = ~n6990 & ~n6992 ;
  assign n6994 = ~n6988 & n6993 ;
  assign n6995 = n1671 & ~n6994 ;
  assign n6996 = ~n6986 & ~n6995 ;
  assign n6997 = n5369 & n5935 ;
  assign n6998 = n2558 & n4869 ;
  assign n6999 = ~n6997 & ~n6998 ;
  assign n7000 = n4185 & ~n6999 ;
  assign n7001 = ~x13 & n1438 ;
  assign n7002 = n3452 & n7001 ;
  assign n7003 = ~n7000 & ~n7002 ;
  assign n7004 = n6996 & n7003 ;
  assign n7005 = n355 & ~n7004 ;
  assign n7006 = n6984 & ~n7005 ;
  assign n7007 = n396 & n4311 ;
  assign n7008 = ~n3059 & ~n4003 ;
  assign n7009 = n252 & n6447 ;
  assign n7010 = ~n7008 & n7009 ;
  assign n7011 = ~n7007 & ~n7010 ;
  assign n7012 = n3740 & n4254 ;
  assign n7013 = n3643 & ~n4247 ;
  assign n7014 = ~n1642 & ~n7013 ;
  assign n7015 = n2039 & ~n7014 ;
  assign n7016 = ~n1642 & ~n4960 ;
  assign n7017 = n2037 & ~n7016 ;
  assign n7018 = ~n1503 & ~n3249 ;
  assign n7019 = ~n2309 & n7018 ;
  assign n7020 = n1919 & ~n7019 ;
  assign n7021 = ~n7017 & ~n7020 ;
  assign n7022 = ~n7015 & n7021 ;
  assign n7023 = ~n7012 & n7022 ;
  assign n7024 = n1330 & ~n7023 ;
  assign n7025 = n7011 & ~n7024 ;
  assign n7026 = ~x13 & ~n7025 ;
  assign n7027 = n7006 & ~n7026 ;
  assign n7028 = ~n6965 & n7027 ;
  assign n7029 = x7 & ~n7028 ;
  assign n7030 = n210 & n2660 ;
  assign n7031 = n86 & n1503 ;
  assign n7032 = ~n830 & n7031 ;
  assign n7033 = n7030 & n7032 ;
  assign n7034 = ~n7029 & ~n7033 ;
  assign n7035 = n7034 ^ x5 ;
  assign n7036 = n7035 ^ n7034 ;
  assign n7037 = n7036 ^ n6953 ;
  assign n7038 = ~n529 & n2257 ;
  assign n7039 = n717 & n3728 ;
  assign n7040 = ~n7038 & ~n7039 ;
  assign n7041 = n6087 & ~n7040 ;
  assign n7042 = ~x6 & n586 ;
  assign n7043 = n2586 & n7042 ;
  assign n7044 = n49 & n399 ;
  assign n7045 = n284 & n587 ;
  assign n7046 = ~n7044 & ~n7045 ;
  assign n7047 = n2598 & ~n7046 ;
  assign n7048 = ~n7043 & ~n7047 ;
  assign n7049 = n21 & ~n7048 ;
  assign n7050 = n529 & n1312 ;
  assign n7051 = ~n7045 & ~n7050 ;
  assign n7052 = n2001 & ~n7051 ;
  assign n7053 = ~n7049 & ~n7052 ;
  assign n7054 = n1582 & n1702 ;
  assign n7055 = n210 & n717 ;
  assign n7056 = n3728 & n4123 ;
  assign n7057 = ~n7055 & ~n7056 ;
  assign n7058 = ~n7054 & n7057 ;
  assign n7059 = n189 & ~n7058 ;
  assign n7060 = n333 & n2469 ;
  assign n7061 = n3264 & n7060 ;
  assign n7062 = ~n7059 & ~n7061 ;
  assign n7063 = n7053 & n7062 ;
  assign n7064 = ~n7041 & n7063 ;
  assign n7065 = n1619 & ~n7064 ;
  assign n7066 = n153 & n2304 ;
  assign n7067 = ~n2187 & ~n7066 ;
  assign n7068 = n7067 ^ n2124 ;
  assign n7069 = n7068 ^ n7067 ;
  assign n7070 = n7067 ^ x7 ;
  assign n7071 = n7070 ^ n7067 ;
  assign n7072 = n7069 & n7071 ;
  assign n7073 = n7072 ^ n7067 ;
  assign n7074 = ~x1 & ~n7073 ;
  assign n7075 = n7074 ^ n7067 ;
  assign n7076 = n3249 & ~n7075 ;
  assign n7077 = n189 & n5598 ;
  assign n7078 = n399 & n1394 ;
  assign n7079 = ~n1085 & n7078 ;
  assign n7080 = ~n7077 & ~n7079 ;
  assign n7081 = ~n7076 & n7080 ;
  assign n7082 = n6647 & ~n7081 ;
  assign n7083 = n291 & n816 ;
  assign n7084 = n1493 & n7083 ;
  assign n7085 = n3509 & n7084 ;
  assign n7086 = ~n7082 & ~n7085 ;
  assign n7087 = ~x1 & n2598 ;
  assign n7088 = n7044 & n7087 ;
  assign n7089 = n333 & n2586 ;
  assign n7090 = n768 & n7089 ;
  assign n7091 = n1084 & ~n2257 ;
  assign n7092 = x7 & ~n210 ;
  assign n7093 = n7091 & n7092 ;
  assign n7094 = n721 & n1715 ;
  assign n7095 = n3756 & n7094 ;
  assign n7096 = ~n7093 & ~n7095 ;
  assign n7097 = ~n7090 & n7096 ;
  assign n7098 = ~x12 & ~n7097 ;
  assign n7099 = ~n7088 & ~n7098 ;
  assign n7100 = n1506 & ~n7099 ;
  assign n7101 = n62 & n1503 ;
  assign n7102 = ~n86 & ~n7101 ;
  assign n7103 = ~x1 & n2387 ;
  assign n7104 = n1073 & n7103 ;
  assign n7105 = ~n7102 & n7104 ;
  assign n7106 = ~n6302 & n7105 ;
  assign n7107 = ~n7100 & ~n7106 ;
  assign n7108 = n7086 & n7107 ;
  assign n7109 = ~n7065 & n7108 ;
  assign n7110 = n7109 ^ x3 ;
  assign n7111 = x3 & ~n7110 ;
  assign n7112 = n7111 ^ n7034 ;
  assign n7113 = n7112 ^ x3 ;
  assign n7114 = n7037 & ~n7113 ;
  assign n7115 = n7114 ^ n7111 ;
  assign n7116 = n7115 ^ x3 ;
  assign n7117 = ~n6953 & n7116 ;
  assign n7118 = n7117 ^ n6953 ;
  assign n7119 = n6948 & ~n7118 ;
  assign n7120 = n7119 ^ x9 ;
  assign n7121 = n7120 ^ n7119 ;
  assign n7122 = n318 & n1528 ;
  assign n7123 = n117 & n7122 ;
  assign n7124 = n1414 & n7123 ;
  assign n7125 = n586 & n6112 ;
  assign n7126 = n6669 & n7125 ;
  assign n7127 = ~x8 & n7126 ;
  assign n7128 = ~n7124 & ~n7127 ;
  assign n7129 = n1598 & n3649 ;
  assign n7130 = ~n1669 & n1932 ;
  assign n7131 = n1438 & n7130 ;
  assign n7132 = ~n7129 & ~n7131 ;
  assign n7133 = x7 & ~n1622 ;
  assign n7134 = ~n7132 & n7133 ;
  assign n7135 = n1291 & n1932 ;
  assign n7136 = ~x8 & n7135 ;
  assign n7137 = ~n7134 & ~n7136 ;
  assign n7138 = n354 & ~n7137 ;
  assign n7139 = n153 & n453 ;
  assign n7140 = ~n1581 & n7139 ;
  assign n7141 = n316 & n1498 ;
  assign n7142 = n763 & n2186 ;
  assign n7143 = ~n7141 & ~n7142 ;
  assign n7144 = n7143 ^ x7 ;
  assign n7145 = n7144 ^ n7143 ;
  assign n7146 = n230 & n1598 ;
  assign n7147 = n829 & ~n1630 ;
  assign n7148 = ~x12 & n7147 ;
  assign n7149 = ~n7146 & ~n7148 ;
  assign n7150 = n7149 ^ n7143 ;
  assign n7151 = n7150 ^ n7143 ;
  assign n7152 = ~n7145 & ~n7151 ;
  assign n7153 = n7152 ^ n7143 ;
  assign n7154 = x4 & ~n7153 ;
  assign n7155 = n7154 ^ n7143 ;
  assign n7156 = ~n7140 & n7155 ;
  assign n7157 = ~x6 & ~n7156 ;
  assign n7158 = ~x4 & n731 ;
  assign n7159 = ~x5 & n252 ;
  assign n7160 = n2186 & n7159 ;
  assign n7161 = ~n7158 & ~n7160 ;
  assign n7162 = n1125 & ~n7161 ;
  assign n7163 = ~x7 & n2289 ;
  assign n7164 = n7163 ^ n1503 ;
  assign n7165 = n7162 & n7164 ;
  assign n7166 = ~n7157 & ~n7165 ;
  assign n7167 = n21 & ~n7166 ;
  assign n7168 = ~n2194 & ~n7042 ;
  assign n7169 = n1073 & ~n7168 ;
  assign n7170 = ~n252 & ~n587 ;
  assign n7171 = n638 & ~n1273 ;
  assign n7172 = ~n7170 & n7171 ;
  assign n7173 = ~n7169 & ~n7172 ;
  assign n7174 = n5647 & ~n7173 ;
  assign n7175 = n3649 & n7066 ;
  assign n7176 = ~n1622 & n7175 ;
  assign n7177 = ~x7 & n132 ;
  assign n7178 = n1598 & n7177 ;
  assign n7179 = ~n867 & ~n5647 ;
  assign n7180 = n1932 & ~n2138 ;
  assign n7181 = ~n7179 & n7180 ;
  assign n7182 = ~n7178 & ~n7181 ;
  assign n7183 = ~n1352 & ~n7182 ;
  assign n7184 = ~n7176 & ~n7183 ;
  assign n7185 = ~n7174 & n7184 ;
  assign n7186 = n313 & ~n7185 ;
  assign n7187 = ~n7167 & ~n7186 ;
  assign n7188 = ~n7138 & n7187 ;
  assign n7189 = n7188 ^ x2 ;
  assign n7190 = n7189 ^ n7188 ;
  assign n7191 = n7190 ^ n7128 ;
  assign n7192 = n2186 & n2687 ;
  assign n7193 = ~x12 & n2304 ;
  assign n7194 = n6062 & n7193 ;
  assign n7195 = ~n7192 & ~n7194 ;
  assign n7196 = n230 & ~n7195 ;
  assign n7197 = n85 & n1312 ;
  assign n7198 = n1261 & n7197 ;
  assign n7199 = n1365 & n7198 ;
  assign n7200 = ~n7196 & ~n7199 ;
  assign n7201 = x1 & ~n7200 ;
  assign n7202 = n85 & ~n2218 ;
  assign n7203 = ~n2314 & ~n7202 ;
  assign n7204 = n799 & n7193 ;
  assign n7205 = ~n7203 & n7204 ;
  assign n7206 = n100 & n337 ;
  assign n7212 = x6 ^ x4 ;
  assign n7213 = n7212 ^ x0 ;
  assign n7207 = x6 ^ x0 ;
  assign n7208 = n7207 ^ x6 ;
  assign n7219 = n7208 ^ n2304 ;
  assign n7220 = n7219 ^ x6 ;
  assign n7209 = ~n1073 & n2710 ;
  assign n7210 = ~x7 & n7209 ;
  assign n7211 = n7210 ^ n7208 ;
  assign n7214 = n7213 ^ n7211 ;
  assign n7221 = n7220 ^ n7214 ;
  assign n7222 = n7221 ^ n7213 ;
  assign n7223 = n7213 & n7222 ;
  assign n7224 = n7223 ^ n7208 ;
  assign n7225 = n7224 ^ n7214 ;
  assign n7226 = n7225 ^ n7213 ;
  assign n7227 = n7226 ^ x6 ;
  assign n7228 = n7214 ^ n7213 ;
  assign n7229 = n7228 ^ x6 ;
  assign n7230 = n7225 & n7229 ;
  assign n7231 = n7230 ^ n7208 ;
  assign n7232 = n7231 ^ n7214 ;
  assign n7233 = n7232 ^ n7213 ;
  assign n7234 = n7233 ^ x6 ;
  assign n7235 = n7227 & n7234 ;
  assign n7215 = n7214 ^ n7208 ;
  assign n7216 = n7215 ^ n7213 ;
  assign n7217 = n7216 ^ x6 ;
  assign n7218 = n7216 & n7217 ;
  assign n7236 = n7235 ^ n7218 ;
  assign n7237 = n7236 ^ n7223 ;
  assign n7238 = n7237 ^ n7208 ;
  assign n7239 = n7238 ^ n7214 ;
  assign n7240 = n7239 ^ n7213 ;
  assign n7241 = n7240 ^ x6 ;
  assign n7242 = n7206 & n7241 ;
  assign n7243 = ~n7205 & ~n7242 ;
  assign n7244 = ~n7201 & n7243 ;
  assign n7245 = n7244 ^ x13 ;
  assign n7246 = ~x13 & n7245 ;
  assign n7247 = n7246 ^ n7188 ;
  assign n7248 = n7247 ^ x13 ;
  assign n7249 = n7191 & n7248 ;
  assign n7250 = n7249 ^ n7246 ;
  assign n7251 = n7250 ^ x13 ;
  assign n7252 = n7128 & ~n7251 ;
  assign n7253 = n7252 ^ n7128 ;
  assign n7254 = ~x14 & ~n7253 ;
  assign n7255 = n466 & n5669 ;
  assign n7256 = x0 & n2138 ;
  assign n7257 = ~n798 & ~n7256 ;
  assign n7258 = n7257 ^ x7 ;
  assign n7259 = n7257 ^ x1 ;
  assign n7260 = n7259 ^ x1 ;
  assign n7261 = x8 & n21 ;
  assign n7262 = n7261 ^ x1 ;
  assign n7263 = n7260 & n7262 ;
  assign n7264 = n7263 ^ x1 ;
  assign n7265 = n7258 & ~n7264 ;
  assign n7266 = n7265 ^ x7 ;
  assign n7267 = n100 & ~n7266 ;
  assign n7268 = n309 & n1619 ;
  assign n7269 = ~n7267 & ~n7268 ;
  assign n7270 = ~n7255 & n7269 ;
  assign n7271 = n2257 & ~n7270 ;
  assign n7272 = n1630 & n6081 ;
  assign n7273 = n1492 & n5564 ;
  assign n7274 = n107 & ~n2397 ;
  assign n7275 = ~n2257 & n7274 ;
  assign n7276 = ~n7273 & ~n7275 ;
  assign n7277 = n189 & ~n7276 ;
  assign n7278 = x14 & n1801 ;
  assign n7279 = ~n280 & ~n7278 ;
  assign n7280 = ~x6 & n4691 ;
  assign n7281 = n429 & n7280 ;
  assign n7282 = ~n7279 & n7281 ;
  assign n7283 = ~n7277 & ~n7282 ;
  assign n7284 = n41 & ~n7283 ;
  assign n7285 = n640 & n3981 ;
  assign n7286 = ~n217 & ~n7285 ;
  assign n7287 = x2 & ~n7286 ;
  assign n7288 = ~n6144 & ~n7287 ;
  assign n7289 = n1506 & n2698 ;
  assign n7290 = ~n7288 & n7289 ;
  assign n7291 = ~n7284 & ~n7290 ;
  assign n7292 = ~n7272 & n7291 ;
  assign n7293 = x14 & n1340 ;
  assign n7294 = ~n565 & n7293 ;
  assign n7295 = ~n130 & ~n7294 ;
  assign n7296 = n5295 & ~n7295 ;
  assign n7297 = n22 & n41 ;
  assign n7298 = n7297 ^ n7261 ;
  assign n7299 = n7298 ^ n7296 ;
  assign n7300 = ~x4 & n6253 ;
  assign n7301 = n7300 ^ n2632 ;
  assign n7302 = ~n7297 & ~n7301 ;
  assign n7303 = n7302 ^ n2632 ;
  assign n7304 = ~n7299 & ~n7303 ;
  assign n7305 = n7304 ^ n7302 ;
  assign n7306 = n7305 ^ n2632 ;
  assign n7307 = n7306 ^ n7297 ;
  assign n7308 = ~n7296 & n7307 ;
  assign n7309 = x6 & ~n7308 ;
  assign n7310 = n7292 & ~n7309 ;
  assign n7311 = ~n7271 & n7310 ;
  assign n7312 = n153 & ~n7311 ;
  assign n7313 = ~n7254 & ~n7312 ;
  assign n7314 = n2975 & n6428 ;
  assign n7315 = ~x5 & n7314 ;
  assign n7316 = ~x6 & ~n86 ;
  assign n7317 = n5640 & ~n7316 ;
  assign n7318 = ~n3508 & n7317 ;
  assign n7319 = ~x5 & n1702 ;
  assign n7320 = x6 & n87 ;
  assign n7321 = n7319 & ~n7320 ;
  assign n7322 = x4 & n7321 ;
  assign n7323 = ~n7318 & ~n7322 ;
  assign n7324 = n7322 ^ n207 ;
  assign n7325 = n3649 & n6078 ;
  assign n7326 = n244 & n6362 ;
  assign n7327 = ~n7325 & ~n7326 ;
  assign n7328 = n1214 & ~n3462 ;
  assign n7329 = n7327 & ~n7328 ;
  assign n7330 = n7329 ^ n7323 ;
  assign n7331 = ~n7324 & n7330 ;
  assign n7332 = n7331 ^ n7329 ;
  assign n7333 = n7323 & n7332 ;
  assign n7334 = n2678 & ~n7333 ;
  assign n7335 = ~n3220 & ~n3240 ;
  assign n7336 = n149 & n3509 ;
  assign n7337 = ~n7335 & n7336 ;
  assign n7338 = ~n7334 & ~n7337 ;
  assign n7339 = n1376 & ~n3048 ;
  assign n7340 = n249 & ~n5862 ;
  assign n7341 = ~n2570 & ~n7340 ;
  assign n7342 = n7341 ^ x12 ;
  assign n7343 = n7342 ^ n7341 ;
  assign n7344 = n7343 ^ n7339 ;
  assign n7345 = n2601 ^ x14 ;
  assign n7346 = ~x14 & ~n7345 ;
  assign n7347 = n7346 ^ n7341 ;
  assign n7348 = n7347 ^ x14 ;
  assign n7349 = n7344 & n7348 ;
  assign n7350 = n7349 ^ n7346 ;
  assign n7351 = n7350 ^ x14 ;
  assign n7352 = ~n7339 & ~n7351 ;
  assign n7353 = n7352 ^ n7339 ;
  assign n7354 = x0 & n7353 ;
  assign n7355 = n62 & ~n249 ;
  assign n7356 = n210 & n7355 ;
  assign n7357 = ~n2915 & ~n7356 ;
  assign n7358 = ~n7354 & n7357 ;
  assign n7359 = n149 & ~n7358 ;
  assign n7360 = x5 & n2351 ;
  assign n7361 = ~n266 & ~n1775 ;
  assign n7362 = n7360 & ~n7361 ;
  assign n7363 = n7362 ^ n62 ;
  assign n7364 = n7362 ^ n1246 ;
  assign n7365 = n7364 ^ n1246 ;
  assign n7366 = n7365 ^ n7363 ;
  assign n7367 = x6 & ~n3294 ;
  assign n7368 = ~n1702 & n7367 ;
  assign n7369 = ~n2600 & ~n7368 ;
  assign n7370 = n7369 ^ n230 ;
  assign n7371 = n230 & ~n7370 ;
  assign n7372 = n7371 ^ n1246 ;
  assign n7373 = n7372 ^ n230 ;
  assign n7374 = ~n7366 & ~n7373 ;
  assign n7375 = n7374 ^ n7371 ;
  assign n7376 = n7375 ^ n230 ;
  assign n7377 = n7363 & n7376 ;
  assign n7378 = n7377 ^ n7362 ;
  assign n7379 = ~n7359 & ~n7378 ;
  assign n7380 = n7379 ^ x8 ;
  assign n7381 = n7380 ^ n7379 ;
  assign n7382 = n7381 ^ n7338 ;
  assign n7383 = n731 & n3249 ;
  assign n7384 = n4869 & n7383 ;
  assign n7385 = n6522 & n6958 ;
  assign n7386 = ~x2 & n434 ;
  assign n7387 = ~n649 & ~n1266 ;
  assign n7388 = n3282 & n7387 ;
  assign n7389 = ~n7386 & ~n7388 ;
  assign n7390 = n6062 & ~n7389 ;
  assign n7391 = ~n7385 & ~n7390 ;
  assign n7392 = ~n7384 & n7391 ;
  assign n7393 = n7392 ^ x3 ;
  assign n7394 = ~n7392 & n7393 ;
  assign n7395 = n7394 ^ n7379 ;
  assign n7396 = n7395 ^ n7392 ;
  assign n7397 = ~n7382 & n7396 ;
  assign n7398 = n7397 ^ n7394 ;
  assign n7399 = n7398 ^ n7392 ;
  assign n7400 = n7338 & ~n7399 ;
  assign n7401 = n7400 ^ n7338 ;
  assign n7402 = ~x1 & ~n7401 ;
  assign n7403 = n2352 & n6813 ;
  assign n7404 = n3254 & n6991 ;
  assign n7405 = ~n7403 & ~n7404 ;
  assign n7406 = n1456 & ~n7405 ;
  assign n7407 = ~x14 & n1365 ;
  assign n7408 = n6958 & n7407 ;
  assign n7409 = n210 & n1394 ;
  assign n7410 = n1528 & n1702 ;
  assign n7411 = ~n7409 & ~n7410 ;
  assign n7412 = ~n267 & ~n7411 ;
  assign n7413 = ~n7408 & ~n7412 ;
  assign n7414 = n1261 & ~n7413 ;
  assign n7415 = ~n7406 & ~n7414 ;
  assign n7416 = n308 & ~n7415 ;
  assign n7417 = n2743 & n3282 ;
  assign n7418 = ~x2 & ~n1528 ;
  assign n7419 = ~n7417 & ~n7418 ;
  assign n7420 = n7419 ^ n1394 ;
  assign n7421 = n7420 ^ n7419 ;
  assign n7422 = n7419 ^ n292 ;
  assign n7423 = n7422 ^ n7419 ;
  assign n7424 = n7421 & n7423 ;
  assign n7425 = n7424 ^ n7419 ;
  assign n7426 = ~x4 & ~n7425 ;
  assign n7427 = n7426 ^ n7419 ;
  assign n7428 = n1583 & ~n7427 ;
  assign n7429 = n228 & ~n1528 ;
  assign n7430 = ~n86 & ~n4117 ;
  assign n7431 = ~n248 & ~n7430 ;
  assign n7432 = ~n7429 & ~n7431 ;
  assign n7433 = n1254 & ~n7432 ;
  assign n7434 = n5413 & n6582 ;
  assign n7435 = n434 & n4877 ;
  assign n7436 = ~n7434 & ~n7435 ;
  assign n7437 = ~n7433 & n7436 ;
  assign n7438 = ~n7428 & n7437 ;
  assign n7439 = n2698 & ~n7438 ;
  assign n7440 = n291 & ~n1394 ;
  assign n7441 = n1698 & n1826 ;
  assign n7442 = ~n7440 & ~n7441 ;
  assign n7443 = n107 & ~n7442 ;
  assign n7444 = n4117 & n7159 ;
  assign n7445 = ~n87 & n4214 ;
  assign n7446 = n7445 ^ x5 ;
  assign n7447 = n7446 ^ n7445 ;
  assign n7448 = n7447 ^ n7444 ;
  assign n7449 = n6582 ^ n3296 ;
  assign n7450 = n3296 & n7449 ;
  assign n7451 = n7450 ^ n7445 ;
  assign n7452 = n7451 ^ n3296 ;
  assign n7453 = ~n7448 & n7452 ;
  assign n7454 = n7453 ^ n7450 ;
  assign n7455 = n7454 ^ n3296 ;
  assign n7456 = ~n7444 & n7455 ;
  assign n7457 = n7456 ^ n7444 ;
  assign n7458 = ~n7443 & ~n7457 ;
  assign n7459 = n2039 & ~n7458 ;
  assign n7460 = ~n7439 & ~n7459 ;
  assign n7461 = ~n7416 & n7460 ;
  assign n7462 = ~n7402 & n7461 ;
  assign n7463 = n7462 ^ x7 ;
  assign n7464 = n7463 ^ n7462 ;
  assign n7465 = x5 & ~n7019 ;
  assign n7466 = ~n5298 & ~n7465 ;
  assign n7467 = n1330 & ~n7466 ;
  assign n7468 = n1630 & n2942 ;
  assign n7469 = ~n7467 & ~n7468 ;
  assign n7470 = n2974 & ~n7469 ;
  assign n7471 = n1433 & ~n1503 ;
  assign n7472 = n1698 & n7471 ;
  assign n7473 = ~n7440 & ~n7472 ;
  assign n7474 = ~x5 & n24 ;
  assign n7475 = ~n7473 & n7474 ;
  assign n7476 = n279 & n2558 ;
  assign n7477 = n6062 & n6428 ;
  assign n7478 = ~n7476 & ~n7477 ;
  assign n7479 = n7478 ^ x5 ;
  assign n7480 = n7479 ^ n7478 ;
  assign n7481 = n7480 ^ n982 ;
  assign n7482 = n1675 ^ n244 ;
  assign n7483 = n244 & n7482 ;
  assign n7484 = n7483 ^ n7478 ;
  assign n7485 = n7484 ^ n244 ;
  assign n7486 = n7481 & ~n7485 ;
  assign n7487 = n7486 ^ n7483 ;
  assign n7488 = n7487 ^ n244 ;
  assign n7489 = n982 & n7488 ;
  assign n7490 = ~n7475 & ~n7489 ;
  assign n7491 = n1775 & ~n7490 ;
  assign n7492 = ~x6 & n1394 ;
  assign n7493 = n3228 & n7492 ;
  assign n7494 = n4883 & n6428 ;
  assign n7495 = ~n7493 & ~n7494 ;
  assign n7496 = x0 & ~n7495 ;
  assign n7497 = n3896 & n7031 ;
  assign n7498 = ~n7496 & ~n7497 ;
  assign n7499 = n974 & ~n7498 ;
  assign n7500 = ~n7491 & ~n7499 ;
  assign n7501 = ~n7470 & n7500 ;
  assign n7502 = n7501 ^ n7462 ;
  assign n7503 = n7464 & n7502 ;
  assign n7504 = n7503 ^ n7462 ;
  assign n7505 = ~n7315 & n7504 ;
  assign n7506 = x13 & ~n7505 ;
  assign n7507 = ~x12 & n2558 ;
  assign n7508 = n355 & n7507 ;
  assign n7509 = n1411 & n1702 ;
  assign n7510 = n7508 & n7509 ;
  assign n7511 = n466 & ~n1352 ;
  assign n7512 = ~n4986 & ~n7511 ;
  assign n7513 = n7512 ^ n451 ;
  assign n7514 = n7513 ^ n7512 ;
  assign n7515 = n7512 ^ n291 ;
  assign n7516 = n7515 ^ n7512 ;
  assign n7517 = n7514 & n7516 ;
  assign n7518 = n7517 ^ n7512 ;
  assign n7519 = x1 & ~n7518 ;
  assign n7520 = n7519 ^ n7512 ;
  assign n7521 = n200 & ~n7520 ;
  assign n7522 = n3868 & n7521 ;
  assign n7523 = ~n7510 & ~n7522 ;
  assign n7524 = ~n7506 & n7523 ;
  assign n7525 = n7313 & n7524 ;
  assign n7526 = n7525 ^ n7119 ;
  assign n7527 = n7121 & n7526 ;
  assign n7528 = n7527 ^ n7119 ;
  assign n7529 = n7528 ^ n6856 ;
  assign n7530 = ~n6857 & ~n7529 ;
  assign n7531 = n7530 ^ n7527 ;
  assign n7532 = n7531 ^ n7119 ;
  assign n7533 = n7532 ^ x10 ;
  assign n7534 = n6856 & n7533 ;
  assign n7535 = n7534 ^ n6856 ;
  assign n7536 = n7535 ^ n6856 ;
  assign n7537 = x15 & ~n7536 ;
  assign n7538 = n1264 & n7492 ;
  assign n7539 = n1715 & n7538 ;
  assign n7540 = n1260 & n1562 ;
  assign n7541 = ~x4 & n7540 ;
  assign n7542 = n1248 & n7541 ;
  assign n7543 = ~n7539 & ~n7542 ;
  assign n7544 = n2472 & ~n7543 ;
  assign n7545 = x7 & ~n558 ;
  assign n7546 = ~n199 & ~n7545 ;
  assign n7549 = ~n167 & ~n603 ;
  assign n7547 = ~x8 & n1706 ;
  assign n7548 = n6814 & n7547 ;
  assign n7550 = n7549 ^ n7548 ;
  assign n7551 = n7550 ^ n7548 ;
  assign n7552 = n1877 & n3018 ;
  assign n7553 = n7552 ^ n7548 ;
  assign n7554 = ~n7551 & n7553 ;
  assign n7555 = n7554 ^ n7548 ;
  assign n7556 = ~n7546 & n7555 ;
  assign n7557 = ~n7544 & ~n7556 ;
  assign n7558 = ~x8 & n1790 ;
  assign n7559 = ~n2157 & ~n7558 ;
  assign n7560 = x12 & n2351 ;
  assign n7561 = ~n7559 & n7560 ;
  assign n7562 = n1733 & n2302 ;
  assign n7563 = n1365 & n7562 ;
  assign n7564 = ~n7561 & ~n7563 ;
  assign n7565 = n207 & n2123 ;
  assign n7566 = ~n7564 & n7565 ;
  assign n7567 = n7557 & ~n7566 ;
  assign n7568 = n1670 & n3107 ;
  assign n7569 = n394 & n1528 ;
  assign n7570 = n1708 & n7569 ;
  assign n7571 = ~n7568 & ~n7570 ;
  assign n7572 = ~n1716 & ~n7571 ;
  assign n7573 = n3267 & n5940 ;
  assign n7574 = n5961 & n6401 ;
  assign n7575 = ~n7573 & ~n7574 ;
  assign n7576 = ~n7572 & n7575 ;
  assign n7577 = n189 & ~n7576 ;
  assign n7578 = n1312 & n3314 ;
  assign n7579 = n291 ^ x2 ;
  assign n7580 = n7579 ^ n291 ;
  assign n7581 = ~n1276 & n2535 ;
  assign n7582 = n7581 ^ n291 ;
  assign n7583 = ~n7580 & ~n7582 ;
  assign n7584 = n7583 ^ n291 ;
  assign n7585 = ~n7578 & ~n7584 ;
  assign n7586 = n3969 & ~n7585 ;
  assign n7587 = ~x7 & ~n250 ;
  assign n7588 = ~n6896 & n7492 ;
  assign n7589 = x2 & n7588 ;
  assign n7590 = ~n7587 & n7589 ;
  assign n7591 = ~n7586 & ~n7590 ;
  assign n7592 = n3172 & ~n7591 ;
  assign n7593 = n1267 & n3282 ;
  assign n7594 = n4048 & n7593 ;
  assign n7595 = n1230 & n1503 ;
  assign n7596 = n72 & n7595 ;
  assign n7597 = n655 & ~n1433 ;
  assign n7598 = n1642 & n7597 ;
  assign n7599 = ~n7596 & ~n7598 ;
  assign n7602 = n7599 ^ x0 ;
  assign n7603 = n7602 ^ n7599 ;
  assign n7600 = n7599 ^ x12 ;
  assign n7601 = n7600 ^ n7599 ;
  assign n7604 = n7603 ^ n7601 ;
  assign n7605 = ~n2138 & ~n2309 ;
  assign n7606 = n7605 ^ n2304 ;
  assign n7607 = n7606 ^ n2304 ;
  assign n7608 = n2304 ^ n1230 ;
  assign n7609 = n7608 ^ n2304 ;
  assign n7610 = ~n7607 & ~n7609 ;
  assign n7611 = n7610 ^ n2304 ;
  assign n7612 = x6 & n7611 ;
  assign n7613 = n7612 ^ n2304 ;
  assign n7614 = n7613 ^ n7599 ;
  assign n7615 = n7614 ^ n7599 ;
  assign n7616 = n7615 ^ n7603 ;
  assign n7617 = ~n7603 & ~n7616 ;
  assign n7618 = n7617 ^ n7603 ;
  assign n7619 = n7604 & ~n7618 ;
  assign n7620 = n7619 ^ n7617 ;
  assign n7621 = n7620 ^ n7599 ;
  assign n7622 = n7621 ^ n7603 ;
  assign n7623 = ~x2 & n7622 ;
  assign n7624 = n7623 ^ n7599 ;
  assign n7625 = ~n7594 & n7624 ;
  assign n7626 = n6670 & ~n7625 ;
  assign n7627 = ~n7592 & ~n7626 ;
  assign n7628 = ~n7577 & n7627 ;
  assign n7629 = n384 & ~n7628 ;
  assign n7630 = n17 & n277 ;
  assign n7631 = n5021 & n7630 ;
  assign n7632 = n1671 & n4775 ;
  assign n7633 = ~x0 & n247 ;
  assign n7634 = n7632 & n7633 ;
  assign n7635 = n207 & ~n1489 ;
  assign n7636 = n2360 & n7635 ;
  assign n7637 = ~n7634 & ~n7636 ;
  assign n7638 = ~x7 & ~n7637 ;
  assign n7639 = ~n7631 & ~n7638 ;
  assign n7640 = n364 & ~n7639 ;
  assign n7641 = ~n7629 & ~n7640 ;
  assign n7642 = n7567 & n7641 ;
  assign n7643 = ~x5 & ~n7642 ;
  assign n7644 = n247 & n1256 ;
  assign n7645 = n1058 & n7644 ;
  assign n7646 = n1482 & n1551 ;
  assign n7647 = n5852 & n7646 ;
  assign n7648 = ~n7645 & ~n7647 ;
  assign n7649 = n1503 & ~n7648 ;
  assign n7650 = n1256 & n2304 ;
  assign n7651 = n2181 & n2929 ;
  assign n7652 = n7650 & n7651 ;
  assign n7653 = n556 & n1264 ;
  assign n7654 = n264 & n2362 ;
  assign n7655 = n7653 & n7654 ;
  assign n7656 = ~n7652 & ~n7655 ;
  assign n7657 = ~n7649 & n7656 ;
  assign n7658 = x1 & ~n7657 ;
  assign n7659 = ~x7 & n3508 ;
  assign n7660 = n5496 & n7659 ;
  assign n7661 = ~n338 & ~n1137 ;
  assign n7662 = n404 & n1716 ;
  assign n7663 = ~n7661 & n7662 ;
  assign n7664 = ~n7660 & ~n7663 ;
  assign n7665 = n17 & ~n7664 ;
  assign n7666 = n1248 & n1551 ;
  assign n7667 = n5936 & n7666 ;
  assign n7668 = n7667 ^ x8 ;
  assign n7669 = n7668 ^ n7667 ;
  assign n7670 = n7669 ^ n7665 ;
  assign n7671 = n395 ^ x0 ;
  assign n7672 = n7671 ^ n395 ;
  assign n7676 = n3056 ^ n404 ;
  assign n7673 = n7672 ^ n395 ;
  assign n7674 = n7672 ^ n404 ;
  assign n7675 = ~n7673 & n7674 ;
  assign n7677 = n7676 ^ n7675 ;
  assign n7678 = n7672 & n7677 ;
  assign n7679 = n7678 ^ n3056 ;
  assign n7680 = n7679 ^ n7672 ;
  assign n7681 = n7680 ^ x0 ;
  assign n7682 = n338 & n7681 ;
  assign n7683 = n1420 & n7197 ;
  assign n7684 = ~n7682 & ~n7683 ;
  assign n7685 = n7684 ^ n1952 ;
  assign n7686 = ~n7684 & ~n7685 ;
  assign n7687 = n7686 ^ n7667 ;
  assign n7688 = n7687 ^ n7684 ;
  assign n7689 = n7670 & ~n7688 ;
  assign n7690 = n7689 ^ n7686 ;
  assign n7691 = n7690 ^ n7684 ;
  assign n7692 = ~n7665 & ~n7691 ;
  assign n7693 = n7692 ^ n7665 ;
  assign n7694 = n364 & n7693 ;
  assign n7695 = ~n7658 & ~n7694 ;
  assign n7696 = n31 & n1483 ;
  assign n7697 = x6 & n7696 ;
  assign n7698 = n1020 & n1248 ;
  assign n7699 = n7697 & n7698 ;
  assign n7700 = ~x2 & n357 ;
  assign n7701 = ~n4738 & ~n5521 ;
  assign n7702 = n1265 & ~n7701 ;
  assign n7703 = ~n7697 & ~n7702 ;
  assign n7704 = n7700 & ~n7703 ;
  assign n7705 = n18 & n3068 ;
  assign n7706 = n5505 & n7705 ;
  assign n7707 = n73 & n1652 ;
  assign n7708 = n1285 & n7707 ;
  assign n7709 = ~n7706 & ~n7708 ;
  assign n7710 = n1248 & ~n7709 ;
  assign n7711 = x9 & ~n2225 ;
  assign n7712 = ~n1562 & ~n7711 ;
  assign n7713 = n2582 & n7560 ;
  assign n7714 = ~n7712 & n7713 ;
  assign n7715 = ~n7710 & ~n7714 ;
  assign n7716 = ~n7704 & n7715 ;
  assign n7717 = n189 & ~n7716 ;
  assign n7718 = n4869 & n7632 ;
  assign n7719 = n3439 & n6814 ;
  assign n7720 = ~n7718 & ~n7719 ;
  assign n7721 = ~n558 & ~n7720 ;
  assign n7722 = n1623 & ~n1943 ;
  assign n7723 = n394 & n7722 ;
  assign n7724 = ~n7721 & ~n7723 ;
  assign n7725 = n6169 & ~n7724 ;
  assign n7726 = n3437 & n5345 ;
  assign n7727 = ~n7719 & ~n7726 ;
  assign n7728 = n308 & n1482 ;
  assign n7729 = ~n1101 & ~n7728 ;
  assign n7730 = ~n7727 & ~n7729 ;
  assign n7731 = ~n7725 & ~n7730 ;
  assign n7732 = ~n7717 & n7731 ;
  assign n7733 = ~n7699 & n7732 ;
  assign n7734 = n7695 & n7733 ;
  assign n7735 = ~n1489 & ~n2452 ;
  assign n7736 = ~n1283 & ~n7735 ;
  assign n7737 = n3532 & ~n7736 ;
  assign n7738 = x12 & ~n6396 ;
  assign n7739 = n1669 & n7738 ;
  assign n7740 = ~n3095 & ~n7739 ;
  assign n7741 = ~x4 & ~n7740 ;
  assign n7742 = n18 & n1438 ;
  assign n7743 = n1264 & n2558 ;
  assign n7744 = ~n1265 & ~n6427 ;
  assign n7745 = ~n7743 & n7744 ;
  assign n7746 = n7745 ^ x6 ;
  assign n7747 = n7746 ^ n7745 ;
  assign n7748 = n7747 ^ n7742 ;
  assign n7749 = ~x8 & n1256 ;
  assign n7750 = n7749 ^ n253 ;
  assign n7751 = n253 & n7750 ;
  assign n7752 = n7751 ^ n7745 ;
  assign n7753 = n7752 ^ n253 ;
  assign n7754 = ~n7748 & ~n7753 ;
  assign n7755 = n7754 ^ n7751 ;
  assign n7756 = n7755 ^ n253 ;
  assign n7757 = ~n7742 & n7756 ;
  assign n7758 = n7757 ^ n7742 ;
  assign n7759 = ~n7741 & ~n7758 ;
  assign n7760 = n7759 ^ x8 ;
  assign n7761 = n7760 ^ x7 ;
  assign n7762 = n7761 ^ n7759 ;
  assign n7763 = n7762 ^ n7761 ;
  assign n7764 = n7763 ^ n7760 ;
  assign n7765 = n7764 ^ n7761 ;
  assign n7766 = n7765 ^ n7760 ;
  assign n7767 = n7766 ^ n7764 ;
  assign n7768 = n2977 ^ x6 ;
  assign n7769 = n2977 ^ x12 ;
  assign n7770 = n7769 ^ x12 ;
  assign n7771 = n1435 ^ x12 ;
  assign n7772 = ~n7770 & n7771 ;
  assign n7773 = n7772 ^ x12 ;
  assign n7774 = n7768 & ~n7773 ;
  assign n7775 = n7774 ^ x6 ;
  assign n7776 = n7775 ^ n7760 ;
  assign n7777 = n7776 ^ n7766 ;
  assign n7778 = n7767 & ~n7777 ;
  assign n7779 = n7778 ^ n7760 ;
  assign n7780 = n7779 ^ n7766 ;
  assign n7781 = n7780 ^ n7764 ;
  assign n7782 = n1234 & n1779 ;
  assign n7783 = ~n2909 & ~n7782 ;
  assign n7784 = n7783 ^ n7778 ;
  assign n7785 = n7784 ^ n7760 ;
  assign n7786 = n7764 & ~n7785 ;
  assign n7787 = n7786 ^ n7766 ;
  assign n7788 = n7787 ^ n7764 ;
  assign n7789 = ~n7781 & n7788 ;
  assign n7790 = n7789 ^ n7778 ;
  assign n7791 = n7790 ^ n7760 ;
  assign n7792 = n7791 ^ n7766 ;
  assign n7793 = n7792 ^ n7764 ;
  assign n7794 = n7793 ^ x8 ;
  assign n7795 = n221 & ~n7794 ;
  assign n7796 = ~n7737 & ~n7795 ;
  assign n7797 = n692 & ~n7796 ;
  assign n7798 = ~n1503 & ~n6304 ;
  assign n7799 = n3643 ^ n1747 ;
  assign n7800 = n1312 & n7799 ;
  assign n7801 = n7800 ^ n1747 ;
  assign n7802 = ~n7798 & n7801 ;
  assign n7803 = n4499 & n7802 ;
  assign n7804 = n1758 ^ x0 ;
  assign n7805 = n7804 ^ x7 ;
  assign n7812 = n7805 ^ n7804 ;
  assign n7806 = n7805 ^ n4801 ;
  assign n7807 = n7806 ^ n7804 ;
  assign n7808 = n7805 ^ n1758 ;
  assign n7809 = n7808 ^ n4801 ;
  assign n7810 = n7809 ^ n7807 ;
  assign n7811 = ~n7807 & ~n7810 ;
  assign n7813 = n7812 ^ n7811 ;
  assign n7814 = n7813 ^ n7807 ;
  assign n7815 = n7804 ^ n1530 ;
  assign n7816 = n7811 ^ n7807 ;
  assign n7817 = n7815 & ~n7816 ;
  assign n7818 = n7817 ^ n7804 ;
  assign n7819 = ~n7814 & n7818 ;
  assign n7820 = n7819 ^ n7804 ;
  assign n7821 = n7820 ^ x0 ;
  assign n7822 = n7821 ^ n7804 ;
  assign n7823 = n1598 & n7822 ;
  assign n7824 = ~x0 & n2225 ;
  assign n7825 = n587 & n7824 ;
  assign n7826 = x9 & n587 ;
  assign n7827 = x0 & ~n3069 ;
  assign n7828 = ~n7826 & ~n7827 ;
  assign n7829 = n17 & ~n7828 ;
  assign n7830 = ~n244 & n7829 ;
  assign n7831 = ~n7825 & ~n7830 ;
  assign n7834 = n6616 ^ x9 ;
  assign n7835 = n7834 ^ n6616 ;
  assign n7832 = n6616 ^ n1259 ;
  assign n7833 = n7832 ^ n6616 ;
  assign n7836 = n7835 ^ n7833 ;
  assign n7837 = ~x7 & n1489 ;
  assign n7838 = n7837 ^ n6616 ;
  assign n7839 = n7838 ^ n6616 ;
  assign n7840 = n7839 ^ n7835 ;
  assign n7841 = n7835 & ~n7840 ;
  assign n7842 = n7841 ^ n7835 ;
  assign n7843 = ~n7836 & n7842 ;
  assign n7844 = n7843 ^ n7841 ;
  assign n7845 = n7844 ^ n6616 ;
  assign n7846 = n7845 ^ n7835 ;
  assign n7847 = x0 & ~n7846 ;
  assign n7848 = n7847 ^ n6616 ;
  assign n7849 = n1528 & ~n7848 ;
  assign n7850 = n7831 & ~n7849 ;
  assign n7851 = ~n7823 & n7850 ;
  assign n7852 = n394 & ~n7851 ;
  assign n7853 = ~x4 & x10 ;
  assign n7854 = n403 & ~n2709 ;
  assign n7855 = x7 & n7854 ;
  assign n7856 = ~n1404 & n7855 ;
  assign n7857 = n86 & n1252 ;
  assign n7858 = n1312 & n7857 ;
  assign n7859 = n277 & ~n5919 ;
  assign n7860 = ~n7858 & ~n7859 ;
  assign n7863 = n7860 ^ n7605 ;
  assign n7864 = n7863 ^ n7860 ;
  assign n7861 = n7860 ^ n277 ;
  assign n7862 = n7861 ^ n7860 ;
  assign n7865 = n7864 ^ n7862 ;
  assign n7866 = n7860 ^ x9 ;
  assign n7867 = n7866 ^ n7860 ;
  assign n7868 = n7867 ^ n7864 ;
  assign n7869 = n7864 & n7868 ;
  assign n7870 = n7869 ^ n7864 ;
  assign n7871 = n7865 & n7870 ;
  assign n7872 = n7871 ^ n7869 ;
  assign n7873 = n7872 ^ n7860 ;
  assign n7874 = n7873 ^ n7864 ;
  assign n7875 = ~x0 & ~n7874 ;
  assign n7876 = n7875 ^ n7860 ;
  assign n7877 = ~n7856 & n7876 ;
  assign n7878 = n7853 & ~n7877 ;
  assign n7879 = n403 & n2386 ;
  assign n7880 = n692 & n7879 ;
  assign n7881 = n7880 ^ x4 ;
  assign n7882 = n7881 ^ n7880 ;
  assign n7883 = n7882 ^ n7878 ;
  assign n7884 = ~x12 & n4801 ;
  assign n7885 = n3643 & n7884 ;
  assign n7886 = ~n17 & ~n6428 ;
  assign n7887 = n257 & ~n1435 ;
  assign n7888 = ~n7886 & n7887 ;
  assign n7889 = n2186 & n3196 ;
  assign n7890 = ~n7888 & ~n7889 ;
  assign n7891 = n7890 ^ x0 ;
  assign n7892 = n7891 ^ n7890 ;
  assign n7893 = n7892 ^ n7885 ;
  assign n7894 = n86 & n257 ;
  assign n7895 = n7894 ^ n2225 ;
  assign n7896 = n2225 & n7895 ;
  assign n7897 = n7896 ^ n7890 ;
  assign n7898 = n7897 ^ n2225 ;
  assign n7899 = n7893 & ~n7898 ;
  assign n7900 = n7899 ^ n7896 ;
  assign n7901 = n7900 ^ n2225 ;
  assign n7902 = ~n7885 & n7901 ;
  assign n7903 = n7902 ^ n7885 ;
  assign n7904 = n7903 ^ x6 ;
  assign n7905 = n7903 & n7904 ;
  assign n7906 = n7905 ^ n7880 ;
  assign n7907 = n7906 ^ n7903 ;
  assign n7908 = ~n7883 & n7907 ;
  assign n7909 = n7908 ^ n7905 ;
  assign n7910 = n7909 ^ n7903 ;
  assign n7911 = ~n7878 & n7910 ;
  assign n7912 = n7911 ^ n7878 ;
  assign n7913 = ~n7852 & ~n7912 ;
  assign n7914 = ~n7803 & n7913 ;
  assign n7915 = n2038 & ~n7914 ;
  assign n7916 = n18 & n1320 ;
  assign n7917 = n533 & n7916 ;
  assign n7918 = n532 & n4052 ;
  assign n7919 = ~n1489 & ~n1779 ;
  assign n7920 = n7918 & n7919 ;
  assign n7921 = ~n7917 & ~n7920 ;
  assign n7922 = n20 & ~n7921 ;
  assign n7923 = ~n926 & n1772 ;
  assign n7924 = ~x6 & ~n7923 ;
  assign n7925 = ~x7 & n1530 ;
  assign n7926 = ~n3228 & ~n7925 ;
  assign n7927 = n7924 & n7926 ;
  assign n7928 = ~x2 & n2138 ;
  assign n7929 = n2405 ^ n1264 ;
  assign n7930 = n7929 ^ n2405 ;
  assign n7931 = n2405 ^ x7 ;
  assign n7932 = n7930 & ~n7931 ;
  assign n7933 = n7932 ^ n2405 ;
  assign n7934 = ~n7928 & ~n7933 ;
  assign n7935 = n7927 & n7934 ;
  assign n7936 = n20 & n1340 ;
  assign n7937 = ~n1551 & n7936 ;
  assign n7938 = ~n7935 & ~n7937 ;
  assign n7939 = n1698 & ~n4691 ;
  assign n7940 = ~n7938 & n7939 ;
  assign n7941 = ~n7922 & ~n7940 ;
  assign n7942 = n357 & ~n7941 ;
  assign n7943 = ~n7915 & ~n7942 ;
  assign n7944 = ~n2225 & ~n2445 ;
  assign n7945 = x0 & n98 ;
  assign n7946 = ~n7944 & n7945 ;
  assign n7947 = n250 & n1733 ;
  assign n7948 = n2386 & n7947 ;
  assign n7949 = ~n7946 & ~n7948 ;
  assign n7950 = n1298 & ~n7949 ;
  assign n7951 = x6 & ~n1230 ;
  assign n7952 = ~x10 & ~n2197 ;
  assign n7953 = ~n7925 & ~n7952 ;
  assign n7954 = n7951 & ~n7953 ;
  assign n7955 = x7 & ~x10 ;
  assign n7956 = n394 & ~n7955 ;
  assign n7957 = n6302 & n7956 ;
  assign n7958 = ~n7595 & ~n7957 ;
  assign n7959 = ~n7954 & n7958 ;
  assign n7960 = ~x12 & ~n7959 ;
  assign n7961 = ~x6 & n1256 ;
  assign n7962 = n7605 & n7961 ;
  assign n7963 = n18 & n1273 ;
  assign n7964 = ~n7879 & ~n7963 ;
  assign n7965 = ~n7962 & n7964 ;
  assign n7966 = n7965 ^ x4 ;
  assign n7967 = n7966 ^ n7965 ;
  assign n7968 = n7967 ^ n7960 ;
  assign n7969 = n7960 ^ n7749 ;
  assign n7970 = x7 & n7969 ;
  assign n7971 = n7970 ^ n7965 ;
  assign n7972 = ~n7968 & ~n7971 ;
  assign n7973 = n7972 ^ n7970 ;
  assign n7974 = n7960 & n7973 ;
  assign n7975 = n7974 ^ n7970 ;
  assign n7976 = n7975 ^ n7972 ;
  assign n7977 = n7976 ^ n7960 ;
  assign n7978 = n357 & n7977 ;
  assign n7979 = n167 & n3294 ;
  assign n7980 = x0 & ~n4737 ;
  assign n7981 = n591 & n7980 ;
  assign n7982 = ~n7979 & ~n7981 ;
  assign n7985 = n7982 ^ x0 ;
  assign n7986 = n7985 ^ n7982 ;
  assign n7983 = n7982 ^ n890 ;
  assign n7984 = n7983 ^ n7982 ;
  assign n7987 = n7986 ^ n7984 ;
  assign n7988 = ~x4 & ~x9 ;
  assign n7989 = n7988 ^ n7982 ;
  assign n7990 = n7989 ^ n7982 ;
  assign n7991 = n7990 ^ n7986 ;
  assign n7992 = ~n7986 & ~n7991 ;
  assign n7993 = n7992 ^ n7986 ;
  assign n7994 = ~n7987 & ~n7993 ;
  assign n7995 = n7994 ^ n7992 ;
  assign n7996 = n7995 ^ n7982 ;
  assign n7997 = n7996 ^ n7986 ;
  assign n7998 = ~x10 & n7997 ;
  assign n7999 = n7998 ^ n7982 ;
  assign n8000 = n1503 & ~n7999 ;
  assign n8001 = n206 & ~n1020 ;
  assign n8002 = n2208 & ~n2565 ;
  assign n8003 = n1365 & ~n8002 ;
  assign n8004 = n8001 & n8003 ;
  assign n8005 = ~n8000 & ~n8004 ;
  assign n8006 = ~n7978 & n8005 ;
  assign n8007 = ~n7950 & n8006 ;
  assign n8008 = n221 & ~n8007 ;
  assign n8009 = ~x0 & n2660 ;
  assign n8010 = n3068 & n8009 ;
  assign n8011 = n7963 & n8010 ;
  assign n8012 = n1298 & n2075 ;
  assign n8013 = n570 & n2257 ;
  assign n8014 = ~n8012 & ~n8013 ;
  assign n8015 = n7824 & ~n8014 ;
  assign n8016 = n98 & n8015 ;
  assign n8017 = ~n8011 & ~n8016 ;
  assign n8018 = n1420 & n1669 ;
  assign n8019 = n1779 & n8018 ;
  assign n8020 = n1283 & n2304 ;
  assign n8021 = n2138 & ~n2988 ;
  assign n8022 = ~n1489 & ~n2535 ;
  assign n8023 = ~x8 & n8022 ;
  assign n8024 = ~n8021 & ~n8023 ;
  assign n8025 = ~n8020 & n8024 ;
  assign n8026 = n532 & ~n8025 ;
  assign n8027 = ~n8019 & ~n8026 ;
  assign n8028 = n3671 & ~n8027 ;
  assign n8029 = n8017 & ~n8028 ;
  assign n8030 = ~n8008 & n8029 ;
  assign n8031 = n7943 & n8030 ;
  assign n8032 = ~n7797 & n8031 ;
  assign n8033 = n149 & ~n8032 ;
  assign n8034 = n7734 & ~n8033 ;
  assign n8035 = ~n7643 & n8034 ;
  assign n8036 = x13 & ~n8035 ;
  assign n8037 = n1020 ^ n308 ;
  assign n8038 = ~n284 & n3865 ;
  assign n8039 = n6814 & n8038 ;
  assign n8040 = n49 & n1562 ;
  assign n8041 = ~n6680 & ~n8040 ;
  assign n8042 = n5345 & ~n8041 ;
  assign n8043 = ~n8039 & ~n8042 ;
  assign n8044 = ~x5 & ~n8043 ;
  assign n8045 = n17 & n4592 ;
  assign n8046 = n6814 & n8045 ;
  assign n8047 = ~n38 & ~n86 ;
  assign n8048 = ~x10 & n8047 ;
  assign n8049 = n6264 & n8048 ;
  assign n8050 = ~n8046 & ~n8049 ;
  assign n8051 = ~n8044 & n8050 ;
  assign n8052 = n8051 ^ n8037 ;
  assign n8053 = n1482 ^ n354 ;
  assign n8054 = n1482 ^ n308 ;
  assign n8055 = n8054 ^ n1482 ;
  assign n8056 = n8053 & ~n8055 ;
  assign n8057 = n8056 ^ n1482 ;
  assign n8058 = n8057 ^ n8037 ;
  assign n8059 = ~n8052 & ~n8058 ;
  assign n8060 = n8059 ^ n8056 ;
  assign n8061 = n8060 ^ n1482 ;
  assign n8062 = n8061 ^ n8051 ;
  assign n8063 = n8037 & n8062 ;
  assign n8064 = n8063 ^ n8037 ;
  assign n8065 = ~n8036 & ~n8064 ;
  assign n8066 = ~n7537 & n8065 ;
  assign n8067 = ~n308 & ~n2342 ;
  assign n8068 = n5961 & n8038 ;
  assign n8069 = n5940 & ~n8041 ;
  assign n8070 = ~n8068 & ~n8069 ;
  assign n8071 = ~x7 & ~n8070 ;
  assign n8072 = n1440 & n2752 ;
  assign n8073 = ~x0 & n8072 ;
  assign n8074 = n8047 & n8073 ;
  assign n8075 = n5961 & n8045 ;
  assign n8076 = ~n8074 & ~n8075 ;
  assign n8077 = ~n8071 & n8076 ;
  assign n8078 = ~n355 & ~n5465 ;
  assign n8079 = ~n8077 & ~n8078 ;
  assign n8080 = ~n8067 & n8079 ;
  assign n8081 = n355 ^ x13 ;
  assign n8082 = n210 & n7541 ;
  assign n8083 = n1702 & n7538 ;
  assign n8084 = ~n8082 & ~n8083 ;
  assign n8085 = n257 & ~n8084 ;
  assign n8086 = n8085 ^ n8081 ;
  assign n8087 = n8086 ^ n355 ;
  assign n8088 = n8087 ^ n8086 ;
  assign n8089 = n742 & n3018 ;
  assign n8090 = n3296 & n8089 ;
  assign n8091 = x8 & ~n2021 ;
  assign n8092 = x6 & ~n1732 ;
  assign n8093 = ~n8091 & n8092 ;
  assign n8094 = ~n24 & n1551 ;
  assign n8095 = ~n409 & ~n8094 ;
  assign n8096 = ~n532 & n3643 ;
  assign n8097 = ~n1438 & ~n1581 ;
  assign n8098 = ~n8096 & ~n8097 ;
  assign n8099 = ~n8095 & n8098 ;
  assign n8100 = n8093 & n8099 ;
  assign n8101 = n2331 & n6868 ;
  assign n8102 = ~n78 & n426 ;
  assign n8103 = n1560 & n8102 ;
  assign n8104 = ~n1259 & n8103 ;
  assign n8105 = n1506 & n7961 ;
  assign n8106 = n185 & n8105 ;
  assign n8107 = ~n8104 & ~n8106 ;
  assign n8108 = ~n8101 & n8107 ;
  assign n8109 = ~n8100 & n8108 ;
  assign n8110 = ~x3 & ~n8109 ;
  assign n8111 = n1330 & n2988 ;
  assign n8112 = ~x8 & n8111 ;
  assign n8113 = n21 & n8112 ;
  assign n8114 = ~n4746 & n5510 ;
  assign n8115 = ~n2225 & ~n2710 ;
  assign n8116 = n8115 ^ x0 ;
  assign n8117 = n8116 ^ n8115 ;
  assign n8118 = n8115 ^ n18 ;
  assign n8119 = n8118 ^ n8115 ;
  assign n8120 = ~n8117 & ~n8119 ;
  assign n8121 = n8120 ^ n8115 ;
  assign n8122 = x12 & n8121 ;
  assign n8123 = n8122 ^ n8115 ;
  assign n8124 = n8114 & n8123 ;
  assign n8125 = n1652 & n1969 ;
  assign n8126 = n3296 & n6781 ;
  assign n8127 = ~n8125 & ~n8126 ;
  assign n8128 = n3421 & ~n8127 ;
  assign n8129 = ~n8124 & ~n8128 ;
  assign n8130 = ~n8113 & n8129 ;
  assign n8131 = ~x7 & ~n8130 ;
  assign n8132 = ~n8110 & ~n8131 ;
  assign n8133 = ~n8090 & n8132 ;
  assign n8134 = n286 & ~n8133 ;
  assign n8135 = x10 ^ x6 ;
  assign n8136 = n1073 ^ x10 ;
  assign n8137 = n8136 ^ n1073 ;
  assign n8138 = n5650 ^ n1073 ;
  assign n8139 = n8137 & n8138 ;
  assign n8140 = n8139 ^ n1073 ;
  assign n8141 = ~n8135 & ~n8140 ;
  assign n8142 = n556 & n8141 ;
  assign n8143 = ~n50 & ~n2977 ;
  assign n8144 = n403 & ~n1733 ;
  assign n8145 = ~n8143 & n8144 ;
  assign n8146 = ~n8142 & ~n8145 ;
  assign n8147 = n85 & n404 ;
  assign n8148 = n1530 & n8147 ;
  assign n8149 = ~x1 & ~n8148 ;
  assign n8150 = ~n8146 & ~n8149 ;
  assign n8151 = n354 & ~n1970 ;
  assign n8152 = n1433 & n8151 ;
  assign n8153 = x1 & ~n1772 ;
  assign n8154 = ~n1747 & n8153 ;
  assign n8155 = n8154 ^ n41 ;
  assign n8156 = n1733 ^ x0 ;
  assign n8157 = n8154 ^ x0 ;
  assign n8158 = n8157 ^ x0 ;
  assign n8159 = n8156 & ~n8158 ;
  assign n8160 = n8159 ^ x0 ;
  assign n8161 = n8155 ^ n450 ;
  assign n8162 = n8160 & n8161 ;
  assign n8163 = n8162 ^ n450 ;
  assign n8164 = n8155 & n8163 ;
  assign n8165 = n8164 ^ n8154 ;
  assign n8166 = n8165 ^ n8155 ;
  assign n8167 = ~n8152 & ~n8166 ;
  assign n8168 = n277 & ~n8167 ;
  assign n8169 = ~n8150 & ~n8168 ;
  assign n8170 = n2386 & ~n8169 ;
  assign n8171 = x12 & n1285 ;
  assign n8172 = ~x6 & n1619 ;
  assign n8173 = ~n8171 & ~n8172 ;
  assign n8174 = n8153 & ~n8173 ;
  assign n8175 = ~n8112 & ~n8174 ;
  assign n8176 = n1137 & ~n8175 ;
  assign n8177 = n1551 & n1670 ;
  assign n8178 = n2037 & n8177 ;
  assign n8179 = n793 & n7630 ;
  assign n8180 = n3437 & n7083 ;
  assign n8181 = ~n8179 & ~n8180 ;
  assign n8182 = ~x3 & ~n8181 ;
  assign n8183 = n333 & n7558 ;
  assign n8184 = n6063 & n8183 ;
  assign n8185 = ~n8182 & ~n8184 ;
  assign n8186 = ~x12 & n1503 ;
  assign n8187 = n2977 & n8186 ;
  assign n8188 = ~n8105 & ~n8187 ;
  assign n8189 = n6099 & ~n8188 ;
  assign n8190 = n8185 & ~n8189 ;
  assign n8191 = ~n8178 & n8190 ;
  assign n8192 = ~n8176 & n8191 ;
  assign n8193 = ~n8170 & n8192 ;
  assign n8194 = n2548 & ~n8193 ;
  assign n8195 = ~x8 & n1733 ;
  assign n8196 = n337 & n466 ;
  assign n8197 = n8195 & n8196 ;
  assign n8198 = n5408 & n8197 ;
  assign n8199 = n943 & n5726 ;
  assign n8200 = n6824 & n8199 ;
  assign n8201 = ~n8198 & ~n8200 ;
  assign n8202 = ~n8194 & n8201 ;
  assign n8203 = n235 & n3865 ;
  assign n8204 = ~n4756 & ~n8203 ;
  assign n8205 = n2351 & ~n8204 ;
  assign n8206 = n655 & ~n1404 ;
  assign n8207 = n3708 & n8206 ;
  assign n8208 = n394 & n8207 ;
  assign n8209 = ~x0 & n1551 ;
  assign n8210 = n3701 & n8209 ;
  assign n8211 = ~x2 & ~n8210 ;
  assign n8212 = ~n8208 & n8211 ;
  assign n8213 = ~n8205 & n8212 ;
  assign n8214 = ~n1671 & ~n2157 ;
  assign n8215 = ~n2410 & ~n8214 ;
  assign n8216 = n1234 & n8215 ;
  assign n8217 = ~n8177 & ~n8216 ;
  assign n8218 = n50 & ~n8217 ;
  assign n8219 = ~n1404 & n6124 ;
  assign n8220 = ~n861 & ~n2156 ;
  assign n8221 = x4 & ~n8220 ;
  assign n8222 = ~n2458 & n8221 ;
  assign n8223 = ~n8219 & ~n8222 ;
  assign n8224 = n7961 & ~n8223 ;
  assign n8225 = n307 & n8187 ;
  assign n8226 = x2 & ~n8225 ;
  assign n8227 = ~n8224 & n8226 ;
  assign n8228 = ~n8218 & n8227 ;
  assign n8229 = n185 & ~n8228 ;
  assign n8230 = ~n8213 & n8229 ;
  assign n8231 = n5545 & n7646 ;
  assign n8232 = x4 & n396 ;
  assign n8233 = n7961 & n8232 ;
  assign n8234 = ~n8231 & ~n8233 ;
  assign n8235 = x0 & n2678 ;
  assign n8236 = ~n8234 & n8235 ;
  assign n8237 = ~n8230 & ~n8236 ;
  assign n8238 = n8202 & n8237 ;
  assign n8239 = ~n8134 & n8238 ;
  assign n8240 = n8239 ^ n8086 ;
  assign n8241 = n8240 ^ n8081 ;
  assign n8242 = n8088 & n8241 ;
  assign n8243 = n8242 ^ n8239 ;
  assign n8244 = ~n1703 & ~n6958 ;
  assign n8245 = n2271 & n3249 ;
  assign n8246 = n8244 & ~n8245 ;
  assign n8247 = x8 & n3796 ;
  assign n8248 = ~n8246 & n8247 ;
  assign n8249 = n2931 & n3896 ;
  assign n8250 = ~n8248 & ~n8249 ;
  assign n8251 = n18 & n62 ;
  assign n8252 = n5961 & n8251 ;
  assign n8253 = n1669 & n1953 ;
  assign n8254 = n4132 & n8253 ;
  assign n8255 = ~n8252 & ~n8254 ;
  assign n8256 = n8255 ^ x9 ;
  assign n8257 = n8256 ^ n8255 ;
  assign n8258 = n8257 ^ n8250 ;
  assign n8259 = n5564 & n7853 ;
  assign n8260 = n210 & ~n7853 ;
  assign n8261 = ~n394 & n8260 ;
  assign n8262 = n1264 & n3981 ;
  assign n8263 = n1702 & n8262 ;
  assign n8264 = ~n8261 & ~n8263 ;
  assign n8265 = ~x8 & ~n8264 ;
  assign n8266 = ~n8259 & ~n8265 ;
  assign n8267 = n8266 ^ x12 ;
  assign n8268 = ~x12 & n8267 ;
  assign n8269 = n8268 ^ n8255 ;
  assign n8270 = n8269 ^ x12 ;
  assign n8271 = n8258 & n8270 ;
  assign n8272 = n8271 ^ n8268 ;
  assign n8273 = n8272 ^ x12 ;
  assign n8274 = n8250 & ~n8273 ;
  assign n8275 = n8274 ^ n8250 ;
  assign n8276 = ~x7 & ~n8275 ;
  assign n8277 = ~n1758 & ~n2445 ;
  assign n8278 = n1234 & n8277 ;
  assign n8279 = x8 & ~n1708 ;
  assign n8280 = n6958 & ~n8279 ;
  assign n8281 = n8278 & n8280 ;
  assign n8282 = n205 & n2445 ;
  assign n8283 = n266 & n4775 ;
  assign n8284 = n8282 & n8283 ;
  assign n8285 = ~n8281 & ~n8284 ;
  assign n8286 = ~n8276 & n8285 ;
  assign n8287 = n8239 & n8286 ;
  assign n8288 = n8287 ^ n8081 ;
  assign n8289 = n8243 & ~n8288 ;
  assign n8290 = n8289 ^ n8287 ;
  assign n8291 = ~n8081 & n8290 ;
  assign n8292 = n8291 ^ n8242 ;
  assign n8293 = n8292 ^ x13 ;
  assign n8294 = n8293 ^ n8239 ;
  assign n8295 = ~n247 & n450 ;
  assign n8296 = n1438 & n6421 ;
  assign n8297 = ~x8 & n3369 ;
  assign n8298 = ~n8296 & ~n8297 ;
  assign n8299 = n816 ^ x2 ;
  assign n8300 = n8299 ^ x2 ;
  assign n8301 = n8300 ^ n469 ;
  assign n8302 = n450 ^ n207 ;
  assign n8303 = ~n450 & n8302 ;
  assign n8304 = n8303 ^ x2 ;
  assign n8305 = n8304 ^ n450 ;
  assign n8306 = ~n8301 & n8305 ;
  assign n8307 = n8306 ^ n8303 ;
  assign n8308 = n8307 ^ n450 ;
  assign n8309 = n469 & ~n8308 ;
  assign n8310 = n8309 ^ n469 ;
  assign n8311 = ~n8298 & n8310 ;
  assign n8312 = ~n8295 & n8311 ;
  assign n8313 = n2410 & n7409 ;
  assign n8314 = n8313 ^ n1702 ;
  assign n8315 = n8314 ^ n8313 ;
  assign n8316 = n8313 ^ n7540 ;
  assign n8317 = n8316 ^ n8313 ;
  assign n8318 = n8315 & n8317 ;
  assign n8319 = n8318 ^ n8313 ;
  assign n8320 = x4 & n8319 ;
  assign n8321 = n8320 ^ n8313 ;
  assign n8322 = ~n558 & n8321 ;
  assign n8323 = ~n8312 & ~n8322 ;
  assign n8324 = x4 & n4592 ;
  assign n8325 = n8324 ^ n49 ;
  assign n8326 = n5650 & n8325 ;
  assign n8327 = n8253 & n8326 ;
  assign n8328 = n528 & n1438 ;
  assign n8329 = n1747 & n8328 ;
  assign n8330 = n77 & n1542 ;
  assign n8331 = n8330 ^ x10 ;
  assign n8332 = n8331 ^ n8330 ;
  assign n8333 = n8332 ^ n8329 ;
  assign n8334 = n8047 ^ n278 ;
  assign n8335 = n8047 & n8334 ;
  assign n8336 = n8335 ^ n8330 ;
  assign n8337 = n8336 ^ n8047 ;
  assign n8338 = n8333 & n8337 ;
  assign n8339 = n8338 ^ n8335 ;
  assign n8340 = n8339 ^ n8047 ;
  assign n8341 = ~n8329 & n8340 ;
  assign n8342 = n8341 ^ n8329 ;
  assign n8343 = n1669 & n8342 ;
  assign n8344 = ~n1503 & ~n1581 ;
  assign n8345 = n6773 & ~n8344 ;
  assign n8346 = x13 & n8345 ;
  assign n8347 = n120 & n1440 ;
  assign n8348 = n2704 & n8347 ;
  assign n8349 = ~n8346 & ~n8348 ;
  assign n8350 = ~n8343 & n8349 ;
  assign n8351 = n1786 & ~n8350 ;
  assign n8352 = ~n1330 & ~n1420 ;
  assign n8353 = n1303 & n8352 ;
  assign n8354 = n2223 & n8353 ;
  assign n8355 = ~n278 & n8354 ;
  assign n8356 = ~n38 & ~n907 ;
  assign n8357 = n3296 & ~n8356 ;
  assign n8358 = ~n3839 & ~n8357 ;
  assign n8359 = n2410 & ~n8358 ;
  assign n8360 = n1733 & n8328 ;
  assign n8361 = ~x6 & n8360 ;
  assign n8362 = n1559 & n5817 ;
  assign n8363 = ~n8361 & ~n8362 ;
  assign n8364 = ~n8359 & n8363 ;
  assign n8365 = ~n8355 & n8364 ;
  assign n8366 = n2277 & ~n8365 ;
  assign n8367 = ~n8351 & ~n8366 ;
  assign n8368 = ~n8327 & n8367 ;
  assign n8369 = n2041 & ~n8368 ;
  assign n8370 = n8323 & ~n8369 ;
  assign n8371 = x10 ^ x0 ;
  assign n8372 = ~n1078 & n4505 ;
  assign n8373 = ~n235 & n8372 ;
  assign n8374 = ~n32 & ~n8373 ;
  assign n8375 = n8374 ^ x10 ;
  assign n8376 = n8375 ^ n8374 ;
  assign n8377 = n8376 ^ n8371 ;
  assign n8378 = ~n1433 & n3282 ;
  assign n8379 = ~n1234 & ~n8378 ;
  assign n8380 = n8379 ^ n41 ;
  assign n8381 = ~n41 & n8380 ;
  assign n8382 = n8381 ^ n8374 ;
  assign n8383 = n8382 ^ n41 ;
  assign n8384 = ~n8377 & n8383 ;
  assign n8385 = n8384 ^ n8381 ;
  assign n8386 = n8385 ^ n41 ;
  assign n8387 = n8371 & ~n8386 ;
  assign n8388 = n817 & n8387 ;
  assign n8389 = n1551 & n6647 ;
  assign n8390 = n8389 ^ n4869 ;
  assign n8391 = n8390 ^ n8389 ;
  assign n8392 = n8389 ^ n1256 ;
  assign n8393 = n8392 ^ n8389 ;
  assign n8394 = n8391 & n8393 ;
  assign n8395 = n8394 ^ n8389 ;
  assign n8396 = ~x14 & n8395 ;
  assign n8397 = n8396 ^ n8389 ;
  assign n8398 = n372 & n8397 ;
  assign n8399 = n229 & n2331 ;
  assign n8400 = n1435 & n2929 ;
  assign n8401 = ~n8399 & ~n8400 ;
  assign n8402 = n469 & ~n8401 ;
  assign n8403 = ~n8398 & ~n8402 ;
  assign n8404 = ~n8388 & n8403 ;
  assign n8405 = x9 & ~n8404 ;
  assign n8406 = ~n457 & n8397 ;
  assign n8407 = n1330 & n1706 ;
  assign n8408 = n503 & n7853 ;
  assign n8409 = ~n8407 & ~n8408 ;
  assign n8410 = n73 & ~n8409 ;
  assign n8411 = ~n1716 & n8410 ;
  assign n8412 = ~n8406 & ~n8411 ;
  assign n8413 = n1084 & ~n8412 ;
  assign n8414 = n503 & ~n2169 ;
  assign n8415 = ~n3068 & ~n8414 ;
  assign n8416 = n7853 & ~n8415 ;
  assign n8417 = n2168 & n8407 ;
  assign n8418 = ~n8416 & ~n8417 ;
  assign n8419 = ~n1943 & ~n8418 ;
  assign n8420 = ~n1330 & ~n4152 ;
  assign n8421 = ~n3545 & ~n8353 ;
  assign n8422 = n365 & ~n8421 ;
  assign n8423 = ~n8420 & n8422 ;
  assign n8424 = ~n8419 & ~n8423 ;
  assign n8425 = ~n8413 & n8424 ;
  assign n8426 = ~n8405 & n8425 ;
  assign n8427 = n1672 & ~n8426 ;
  assign n8428 = n3848 & n6680 ;
  assign n8429 = n3043 & n3865 ;
  assign n8430 = x14 & n8429 ;
  assign n8431 = ~n8428 & ~n8430 ;
  assign n8432 = n318 ^ x3 ;
  assign n8433 = n8432 ^ n318 ;
  assign n8434 = n1085 ^ n318 ;
  assign n8435 = ~n8433 & ~n8434 ;
  assign n8436 = n8435 ^ n318 ;
  assign n8437 = ~n8431 & n8436 ;
  assign n8438 = ~n8427 & ~n8437 ;
  assign n8439 = n8370 & n8438 ;
  assign n8440 = n228 & ~n3453 ;
  assign n8441 = ~n38 & ~n2586 ;
  assign n8442 = ~n134 & ~n8441 ;
  assign n8443 = n2660 & n8442 ;
  assign n8444 = ~n8440 & ~n8443 ;
  assign n8445 = n17 & ~n8444 ;
  assign n8446 = ~n207 & ~n2877 ;
  assign n8447 = n2320 & ~n8446 ;
  assign n8448 = ~n2075 & n8447 ;
  assign n8449 = ~n8445 & ~n8448 ;
  assign n8450 = n205 & ~n8449 ;
  assign n8451 = n38 & n3172 ;
  assign n8452 = n4842 & n8451 ;
  assign n8453 = ~n8450 & ~n8452 ;
  assign n8454 = ~n49 & ~n4593 ;
  assign n8455 = n49 & n2225 ;
  assign n8456 = ~n1719 & ~n8455 ;
  assign n8457 = n798 & ~n8456 ;
  assign n8458 = ~n8454 & n8457 ;
  assign n8459 = n119 & n2330 ;
  assign n8460 = n2331 & n4052 ;
  assign n8461 = ~n1608 & n2977 ;
  assign n8462 = ~n891 & n8461 ;
  assign n8463 = ~n8460 & ~n8462 ;
  assign n8464 = ~n8459 & n8463 ;
  assign n8465 = n1715 & ~n8464 ;
  assign n8466 = ~n8458 & ~n8465 ;
  assign n8467 = ~x6 & ~n8466 ;
  assign n8468 = ~n1530 & n3552 ;
  assign n8469 = x0 & ~n8468 ;
  assign n8470 = n6772 & ~n8469 ;
  assign n8471 = x13 & n1256 ;
  assign n8472 = x10 & n1059 ;
  assign n8473 = ~n8471 & ~n8472 ;
  assign n8474 = ~n8470 & n8473 ;
  assign n8475 = n2277 & ~n8474 ;
  assign n8476 = n1733 & n2387 ;
  assign n8477 = ~n1598 & n8476 ;
  assign n8478 = ~n8475 & ~n8477 ;
  assign n8479 = n5403 & ~n8478 ;
  assign n8480 = ~n8467 & ~n8479 ;
  assign n8481 = n1365 & n7030 ;
  assign n8482 = n1309 & n8481 ;
  assign n8483 = n8480 & ~n8482 ;
  assign n8484 = n8453 & n8483 ;
  assign n8485 = n384 & ~n8484 ;
  assign n8486 = n8439 & ~n8485 ;
  assign n8487 = n1559 & n7280 ;
  assign n8488 = n503 & n1415 ;
  assign n8489 = ~n1309 & ~n8488 ;
  assign n8490 = x1 & ~n8489 ;
  assign n8491 = n3143 & ~n6396 ;
  assign n8492 = ~n8490 & ~n8491 ;
  assign n8493 = n1671 & ~n8492 ;
  assign n8494 = x6 & n3658 ;
  assign n8495 = ~n3154 & ~n3172 ;
  assign n8496 = n8494 & ~n8495 ;
  assign n8497 = ~n8493 & ~n8496 ;
  assign n8498 = ~n8487 & n8497 ;
  assign n8499 = ~n248 & ~n8498 ;
  assign n8500 = n2257 & n8407 ;
  assign n8501 = n3196 & n4134 ;
  assign n8502 = ~n8500 & ~n8501 ;
  assign n8503 = ~x13 & ~n8502 ;
  assign n8504 = ~n1530 & n2988 ;
  assign n8505 = ~x4 & n4506 ;
  assign n8506 = n8504 & n8505 ;
  assign n8507 = n1234 & n2239 ;
  assign n8508 = n1285 ^ x12 ;
  assign n8509 = n8508 ^ n1285 ;
  assign n8510 = n8509 ^ n119 ;
  assign n8511 = n1952 ^ n119 ;
  assign n8512 = ~n269 & ~n8511 ;
  assign n8513 = n8512 ^ n1285 ;
  assign n8514 = ~n8510 & n8513 ;
  assign n8515 = n8514 ^ n8512 ;
  assign n8516 = ~n119 & n8515 ;
  assign n8517 = n8516 ^ n8512 ;
  assign n8518 = n8517 ^ n8514 ;
  assign n8519 = ~n8507 & ~n8518 ;
  assign n8520 = ~n8506 & n8519 ;
  assign n8521 = ~n8503 & n8520 ;
  assign n8522 = n2640 & ~n8521 ;
  assign n8523 = x1 & n17 ;
  assign n8524 = ~x2 & n1484 ;
  assign n8525 = ~n4134 & ~n8524 ;
  assign n8526 = n8525 ^ x13 ;
  assign n8527 = n8526 ^ n8525 ;
  assign n8528 = ~n2600 & ~n3728 ;
  assign n8529 = n8528 ^ n8525 ;
  assign n8530 = n8529 ^ n8525 ;
  assign n8531 = n8527 & ~n8530 ;
  assign n8532 = n8531 ^ n8525 ;
  assign n8533 = x12 & ~n8532 ;
  assign n8534 = n8533 ^ n8525 ;
  assign n8535 = n8523 & ~n8534 ;
  assign n8536 = n1954 & ~n3448 ;
  assign n8537 = n2761 & n8536 ;
  assign n8538 = ~n4780 & n8537 ;
  assign n8539 = ~n8535 & ~n8538 ;
  assign n8540 = ~n8522 & n8539 ;
  assign n8541 = n18 & n7316 ;
  assign n8542 = ~n1534 & ~n8541 ;
  assign n8543 = n266 & ~n8542 ;
  assign n8544 = ~n753 & n5277 ;
  assign n8545 = ~n1598 & ~n4114 ;
  assign n8546 = ~n133 & n5545 ;
  assign n8547 = ~n8545 & n8546 ;
  assign n8548 = ~n8544 & ~n8547 ;
  assign n8549 = n3172 & ~n8548 ;
  assign n8550 = ~n8543 & ~n8549 ;
  assign n8551 = n8540 & n8550 ;
  assign n8552 = ~n8499 & n8551 ;
  assign n8553 = n85 & ~n8552 ;
  assign n8554 = ~n3096 & ~n8251 ;
  assign n8555 = n3728 & ~n8554 ;
  assign n8556 = n799 & n8555 ;
  assign n8557 = n3172 & n4690 ;
  assign n8558 = x6 ^ x1 ;
  assign n8559 = n8558 ^ x6 ;
  assign n8560 = n8559 ^ n318 ;
  assign n8561 = n8468 ^ x10 ;
  assign n8562 = ~x6 & ~n8561 ;
  assign n8563 = n8562 ^ n8468 ;
  assign n8564 = ~n8560 & n8563 ;
  assign n8565 = n8564 ^ n8562 ;
  assign n8566 = n8565 ^ n8468 ;
  assign n8567 = n8566 ^ x6 ;
  assign n8568 = ~n318 & ~n8567 ;
  assign n8569 = n1365 & n8568 ;
  assign n8570 = ~n8557 & ~n8569 ;
  assign n8571 = n2691 & ~n8570 ;
  assign n8572 = n7280 & n8471 ;
  assign n8573 = n1440 & n1598 ;
  assign n8574 = ~n1390 & ~n8573 ;
  assign n8575 = n2038 & ~n8574 ;
  assign n8576 = n1669 & ~n3453 ;
  assign n8577 = n284 & n1598 ;
  assign n8578 = ~n1511 & ~n8577 ;
  assign n8579 = n2906 & ~n8578 ;
  assign n8580 = ~n8576 & ~n8579 ;
  assign n8581 = n1719 & ~n8580 ;
  assign n8582 = ~n8575 & ~n8581 ;
  assign n8583 = ~n8572 & n8582 ;
  assign n8584 = x4 & ~n8583 ;
  assign n8585 = n1303 & ~n1322 ;
  assign n8586 = n5636 & n8585 ;
  assign n8587 = ~n2424 & ~n2906 ;
  assign n8588 = n4592 & n8587 ;
  assign n8589 = ~n267 & n3143 ;
  assign n8590 = ~n8588 & ~n8589 ;
  assign n8591 = n7853 & ~n8590 ;
  assign n8592 = x6 & n6368 ;
  assign n8593 = ~n1484 & ~n8592 ;
  assign n8594 = n532 & ~n8593 ;
  assign n8595 = ~n8591 & ~n8594 ;
  assign n8596 = ~n8586 & n8595 ;
  assign n8597 = n2276 & ~n8596 ;
  assign n8598 = n17 & n49 ;
  assign n8599 = x1 & n291 ;
  assign n8600 = n8598 & n8599 ;
  assign n8601 = ~n8597 & ~n8600 ;
  assign n8602 = ~n8584 & n8601 ;
  assign n8603 = ~n8571 & n8602 ;
  assign n8604 = ~n8556 & n8603 ;
  assign n8605 = n50 & ~n8604 ;
  assign n8606 = ~n8553 & ~n8605 ;
  assign n8607 = n1669 & n3903 ;
  assign n8608 = x4 & n8607 ;
  assign n8609 = n1394 & ~n1489 ;
  assign n8610 = n2567 & n8609 ;
  assign n8611 = n252 & n8251 ;
  assign n8612 = n1435 & n1668 ;
  assign n8613 = ~n8611 & ~n8612 ;
  assign n8614 = ~x1 & ~n1716 ;
  assign n8615 = ~n8613 & n8614 ;
  assign n8616 = ~n8610 & ~n8615 ;
  assign n8617 = ~n3438 & n8616 ;
  assign n8618 = ~x3 & ~n8617 ;
  assign n8619 = n2704 & n3508 ;
  assign n8620 = n1703 & n6813 ;
  assign n8621 = ~x0 & ~n1718 ;
  assign n8622 = n7738 & n8621 ;
  assign n8623 = ~n2278 & n8622 ;
  assign n8624 = ~n8620 & ~n8623 ;
  assign n8625 = ~n8619 & n8624 ;
  assign n8626 = n5505 & ~n8625 ;
  assign n8627 = n8626 ^ x1 ;
  assign n8628 = n8627 ^ n8626 ;
  assign n8629 = n1623 & n2606 ;
  assign n8630 = n2601 & n3439 ;
  assign n8631 = ~n8629 & ~n8630 ;
  assign n8632 = x0 & ~n8631 ;
  assign n8633 = ~n7634 & ~n8632 ;
  assign n8634 = n8633 ^ n8626 ;
  assign n8635 = ~n8628 & ~n8634 ;
  assign n8636 = n8635 ^ n8626 ;
  assign n8637 = ~n8618 & ~n8636 ;
  assign n8638 = ~n8608 & n8637 ;
  assign n8639 = x13 & ~n8638 ;
  assign n8640 = n8251 ^ n6492 ;
  assign n8641 = n8640 ^ n8251 ;
  assign n8642 = n8251 ^ x8 ;
  assign n8643 = n8642 ^ n8251 ;
  assign n8644 = n8641 & n8643 ;
  assign n8645 = n8644 ^ n8251 ;
  assign n8646 = ~x2 & n8645 ;
  assign n8647 = n8646 ^ n8251 ;
  assign n8648 = n425 & n8647 ;
  assign n8649 = ~n1528 & ~n3453 ;
  assign n8650 = n1283 & n2405 ;
  assign n8651 = n8649 & n8650 ;
  assign n8652 = ~n8555 & ~n8651 ;
  assign n8653 = ~n8648 & n8652 ;
  assign n8654 = n117 & ~n8653 ;
  assign n8655 = n1248 & ~n8542 ;
  assign n8656 = x6 & ~n3154 ;
  assign n8657 = x12 & n6396 ;
  assign n8658 = ~n8656 & ~n8657 ;
  assign n8659 = n5935 & n8658 ;
  assign n8660 = n469 & n8659 ;
  assign n8661 = ~n8655 & ~n8660 ;
  assign n8662 = ~n8654 & n8661 ;
  assign n8663 = n2660 & ~n8662 ;
  assign n8664 = ~n8639 & ~n8663 ;
  assign n8665 = n8606 & n8664 ;
  assign n8666 = n249 & n2038 ;
  assign n8667 = n8598 & n8666 ;
  assign n8668 = n8667 ^ n792 ;
  assign n8669 = n8668 ^ x3 ;
  assign n8689 = n8669 ^ n8668 ;
  assign n8670 = n1952 & n3658 ;
  assign n8671 = ~x3 & n8670 ;
  assign n8672 = ~x8 & n1952 ;
  assign n8673 = n890 & n8672 ;
  assign n8674 = n1125 & n8673 ;
  assign n8675 = x2 & n890 ;
  assign n8676 = ~n1823 & n3661 ;
  assign n8677 = ~n8675 & n8676 ;
  assign n8678 = ~x13 & n6678 ;
  assign n8679 = ~n8677 & ~n8678 ;
  assign n8680 = ~n8674 & n8679 ;
  assign n8681 = ~n8671 & n8680 ;
  assign n8682 = n2351 & ~n8681 ;
  assign n8683 = n8682 ^ n8669 ;
  assign n8684 = n8683 ^ n8668 ;
  assign n8685 = n8669 ^ n8667 ;
  assign n8686 = n8685 ^ n8682 ;
  assign n8687 = n8686 ^ n8684 ;
  assign n8688 = ~n8684 & ~n8687 ;
  assign n8690 = n8689 ^ n8688 ;
  assign n8691 = n8690 ^ n8684 ;
  assign n8692 = n1551 & n2549 ;
  assign n8693 = ~n1256 & ~n8692 ;
  assign n8694 = n2277 & ~n8693 ;
  assign n8695 = ~n6396 & n8619 ;
  assign n8696 = ~n8694 & ~n8695 ;
  assign n8697 = n425 & ~n8696 ;
  assign n8698 = n8697 ^ n8668 ;
  assign n8699 = n8688 ^ n8684 ;
  assign n8700 = ~n8698 & ~n8699 ;
  assign n8701 = n8700 ^ n8668 ;
  assign n8702 = ~n8691 & n8701 ;
  assign n8703 = n8702 ^ n8668 ;
  assign n8704 = n8703 ^ n792 ;
  assign n8705 = n8704 ^ n8668 ;
  assign n8706 = n8665 & ~n8705 ;
  assign n8707 = n8706 ^ x9 ;
  assign n8708 = n8707 ^ n8706 ;
  assign n8709 = n550 & n5598 ;
  assign n8710 = n817 & n3421 ;
  assign n8711 = ~n8709 & ~n8710 ;
  assign n8712 = n1733 & ~n8711 ;
  assign n8713 = n85 & n1562 ;
  assign n8714 = n3809 & n8713 ;
  assign n8715 = ~n8712 & ~n8714 ;
  assign n8716 = ~x12 & ~n8715 ;
  assign n8717 = ~n49 & ~n8577 ;
  assign n8718 = n2037 & ~n8717 ;
  assign n8719 = n1283 & n8718 ;
  assign n8720 = ~n8716 & ~n8719 ;
  assign n8721 = n2691 & ~n8720 ;
  assign n8722 = n17 & n252 ;
  assign n8723 = n6991 & n8722 ;
  assign n8724 = ~x8 & n1629 ;
  assign n8725 = ~n2932 & ~n8724 ;
  assign n8726 = ~n6396 & ~n6398 ;
  assign n8727 = n8725 & ~n8726 ;
  assign n8728 = ~n1716 & ~n8727 ;
  assign n8729 = n1528 & n3649 ;
  assign n8730 = ~n207 & n2360 ;
  assign n8731 = ~n8729 & ~n8730 ;
  assign n8732 = ~n6429 & ~n8731 ;
  assign n8733 = ~n2928 & ~n2931 ;
  assign n8734 = ~x0 & n3228 ;
  assign n8735 = ~n6989 & ~n8734 ;
  assign n8736 = ~n8733 & ~n8735 ;
  assign n8737 = ~n8732 & ~n8736 ;
  assign n8738 = ~n8728 & n8737 ;
  assign n8739 = x13 & ~n8738 ;
  assign n8740 = ~x13 & ~n3592 ;
  assign n8741 = n1435 & n1665 ;
  assign n8742 = ~n8740 & ~n8741 ;
  assign n8743 = ~n4688 & n8742 ;
  assign n8744 = ~n1716 & ~n8743 ;
  assign n8745 = x6 & n253 ;
  assign n8746 = n17 & n8745 ;
  assign n8747 = ~n3717 & ~n8746 ;
  assign n8748 = x2 & n244 ;
  assign n8749 = ~n8747 & n8748 ;
  assign n8750 = n3840 & n7547 ;
  assign n8751 = ~n8749 & ~n8750 ;
  assign n8752 = ~n8744 & n8751 ;
  assign n8753 = ~n8739 & n8752 ;
  assign n8754 = ~n8723 & n8753 ;
  assign n8755 = n354 & ~n8754 ;
  assign n8756 = ~n8721 & ~n8755 ;
  assign n8757 = n8756 ^ n8706 ;
  assign n8758 = n8708 & n8757 ;
  assign n8759 = n8758 ^ n8706 ;
  assign n8760 = n8486 & n8759 ;
  assign n8761 = n8760 ^ x7 ;
  assign n8762 = n8761 ^ n8760 ;
  assign n8763 = n8762 ^ n8294 ;
  assign n8764 = n1435 & n1669 ;
  assign n8765 = n3896 & n8764 ;
  assign n8766 = n3821 & n6499 ;
  assign n8767 = ~n7538 & ~n7541 ;
  assign n8768 = ~n1716 & ~n8767 ;
  assign n8769 = ~n8766 & ~n8768 ;
  assign n8770 = ~n8765 & n8769 ;
  assign n8771 = n308 & ~n8770 ;
  assign n8772 = n1941 & n8187 ;
  assign n8773 = n6113 & n6824 ;
  assign n8774 = ~n8772 & ~n8773 ;
  assign n8775 = ~n8771 & n8774 ;
  assign n8776 = n8775 ^ x9 ;
  assign n8777 = x9 & ~n8776 ;
  assign n8778 = n8777 ^ n8760 ;
  assign n8779 = n8778 ^ x9 ;
  assign n8780 = n8763 & ~n8779 ;
  assign n8781 = n8780 ^ n8777 ;
  assign n8782 = n8781 ^ x9 ;
  assign n8783 = ~n8294 & n8782 ;
  assign n8784 = n8783 ^ n8294 ;
  assign n8785 = n8784 ^ x5 ;
  assign n8786 = n8785 ^ n8784 ;
  assign n8787 = n8786 ^ n8080 ;
  assign n8788 = n2421 & n7569 ;
  assign n8789 = n1670 & n2331 ;
  assign n8790 = n1435 & n8172 ;
  assign n8791 = ~n8789 & ~n8790 ;
  assign n8792 = n1814 & ~n8791 ;
  assign n8793 = n98 & n3728 ;
  assign n8794 = n3095 & n8793 ;
  assign n8795 = ~x12 & n2991 ;
  assign n8796 = n249 & n3107 ;
  assign n8797 = ~n8795 & ~n8796 ;
  assign n8798 = n2398 & ~n8797 ;
  assign n8799 = ~n8794 & ~n8798 ;
  assign n8800 = ~n8792 & n8799 ;
  assign n8801 = x1 & ~n8800 ;
  assign n8802 = ~n8788 & ~n8801 ;
  assign n8803 = n50 & ~n8802 ;
  assign n8804 = n2282 ^ n2278 ;
  assign n8805 = ~x1 & ~n8804 ;
  assign n8806 = n8805 ^ n2278 ;
  assign n8807 = n404 & ~n8806 ;
  assign n8808 = n1619 & n8012 ;
  assign n8809 = ~n8807 & ~n8808 ;
  assign n8810 = n7955 & ~n8809 ;
  assign n8811 = ~x7 & n2952 ;
  assign n8812 = n1376 & n4691 ;
  assign n8813 = n8811 & n8812 ;
  assign n8814 = ~x12 & n8745 ;
  assign n8815 = ~n2942 & ~n8814 ;
  assign n8816 = n2391 & ~n8815 ;
  assign n8817 = n1528 & n8793 ;
  assign n8818 = ~n8816 & ~n8817 ;
  assign n8819 = n6670 & ~n8818 ;
  assign n8820 = ~n8813 & ~n8819 ;
  assign n8821 = ~n8810 & n8820 ;
  assign n8822 = n85 & ~n8821 ;
  assign n8823 = ~x0 & ~n1954 ;
  assign n8824 = n7569 & n8823 ;
  assign n8825 = n1702 & n2225 ;
  assign n8826 = n404 & n8825 ;
  assign n8827 = ~n8824 & ~n8826 ;
  assign n8828 = n338 & ~n8827 ;
  assign n8829 = x1 & n8828 ;
  assign n8830 = ~n8822 & ~n8829 ;
  assign n8831 = ~n8803 & n8830 ;
  assign n8832 = n8831 ^ x9 ;
  assign n8833 = x9 & ~n8832 ;
  assign n8834 = n8833 ^ n8784 ;
  assign n8835 = n8834 ^ x9 ;
  assign n8836 = n8787 & n8835 ;
  assign n8837 = n8836 ^ n8833 ;
  assign n8838 = n8837 ^ x9 ;
  assign n8839 = ~n8080 & n8838 ;
  assign n8840 = n8839 ^ n8080 ;
  assign n8841 = n8066 & ~n8840 ;
  assign n8842 = n8841 ^ x11 ;
  assign n8843 = n8842 ^ n8841 ;
  assign n8844 = x6 & n1991 ;
  assign n8845 = n2938 & n8844 ;
  assign n8846 = n396 & n2410 ;
  assign n8847 = n4561 & n8846 ;
  assign n8848 = ~n8845 & ~n8847 ;
  assign n8849 = n2704 & ~n8848 ;
  assign n8850 = n25 & n8849 ;
  assign n8851 = n257 & n263 ;
  assign n8852 = ~n862 & ~n8851 ;
  assign n8853 = ~n38 & ~n2331 ;
  assign n8854 = ~n1706 & n8853 ;
  assign n8855 = ~x0 & n3227 ;
  assign n8856 = ~n8854 & n8855 ;
  assign n8857 = ~n3453 & n8722 ;
  assign n8858 = n1715 & n8857 ;
  assign n8859 = ~n8856 & ~n8858 ;
  assign n8860 = ~n8852 & ~n8859 ;
  assign n8861 = ~n8850 & ~n8860 ;
  assign n8862 = n2042 ^ x13 ;
  assign n8863 = n295 & n7963 ;
  assign n8864 = n3294 & n8863 ;
  assign n8865 = n8864 ^ n8862 ;
  assign n8866 = n8865 ^ n2042 ;
  assign n8867 = n8866 ^ n8865 ;
  assign n8868 = n1256 & n2397 ;
  assign n8869 = n1391 & n8868 ;
  assign n8870 = n24 & n8869 ;
  assign n8871 = n23 & n8296 ;
  assign n8872 = x2 & n8871 ;
  assign n8873 = ~n8870 & ~n8872 ;
  assign n8874 = n98 & n2424 ;
  assign n8875 = n7386 & n8874 ;
  assign n8876 = n1990 ^ n1376 ;
  assign n8877 = n8876 ^ n1990 ;
  assign n8878 = n1990 ^ n25 ;
  assign n8879 = n8878 ^ n1990 ;
  assign n8880 = n8877 & n8879 ;
  assign n8881 = n8880 ^ n1990 ;
  assign n8882 = ~x1 & n8881 ;
  assign n8883 = n8882 ^ n1990 ;
  assign n8884 = n3282 & n8883 ;
  assign n8885 = ~n8875 & ~n8884 ;
  assign n8886 = n7824 & ~n8885 ;
  assign n8887 = n824 & n2661 ;
  assign n8888 = n1953 & n2256 ;
  assign n8889 = n8887 & n8888 ;
  assign n8890 = x8 ^ x0 ;
  assign n8891 = n532 & n1597 ;
  assign n8892 = n1815 & n8891 ;
  assign n8893 = n189 & n1275 ;
  assign n8894 = n2600 & n8893 ;
  assign n8895 = n1456 & ~n2452 ;
  assign n8896 = ~n1291 & ~n8895 ;
  assign n8897 = n880 & n1953 ;
  assign n8898 = ~n8896 & n8897 ;
  assign n8899 = ~n8894 & ~n8898 ;
  assign n8900 = ~n8892 & n8899 ;
  assign n8901 = n8900 ^ x8 ;
  assign n8902 = n8901 ^ n8900 ;
  assign n8903 = n1387 & n2075 ;
  assign n8904 = n1256 & n8903 ;
  assign n8905 = n8904 ^ n8900 ;
  assign n8906 = n8902 & ~n8905 ;
  assign n8907 = n8906 ^ n8900 ;
  assign n8908 = n8890 & ~n8907 ;
  assign n8909 = ~n8889 & ~n8908 ;
  assign n8910 = ~n8886 & n8909 ;
  assign n8911 = n8910 ^ x9 ;
  assign n8912 = n8911 ^ n8910 ;
  assign n8913 = n8912 ^ n8873 ;
  assign n8914 = x5 ^ x4 ;
  assign n8915 = n1623 & n6958 ;
  assign n8916 = n8915 ^ n8607 ;
  assign n8917 = ~n8914 & n8916 ;
  assign n8918 = n8917 ^ n8607 ;
  assign n8919 = ~x7 & n8918 ;
  assign n8920 = ~x5 & n1340 ;
  assign n8921 = n1623 & n2352 ;
  assign n8922 = n8920 & n8921 ;
  assign n8923 = ~n8919 & ~n8922 ;
  assign n8924 = n8187 ^ x2 ;
  assign n8925 = n8924 ^ n8187 ;
  assign n8926 = n8925 ^ n132 ;
  assign n8927 = n394 ^ n132 ;
  assign n8928 = n7650 & ~n8927 ;
  assign n8929 = n8928 ^ n8187 ;
  assign n8930 = ~n8926 & n8929 ;
  assign n8931 = n8930 ^ n8928 ;
  assign n8932 = ~n132 & n8931 ;
  assign n8933 = n8932 ^ n8928 ;
  assign n8934 = n8933 ^ n8930 ;
  assign n8935 = n8923 & ~n8934 ;
  assign n8936 = n8935 ^ x1 ;
  assign n8937 = ~n8935 & n8936 ;
  assign n8938 = n8937 ^ n8910 ;
  assign n8939 = n8938 ^ n8935 ;
  assign n8940 = n8913 & n8939 ;
  assign n8941 = n8940 ^ n8937 ;
  assign n8942 = n8941 ^ n8935 ;
  assign n8943 = n8873 & ~n8942 ;
  assign n8944 = n8943 ^ n8873 ;
  assign n8945 = n8944 ^ n8865 ;
  assign n8946 = n8945 ^ n8862 ;
  assign n8947 = ~n8867 & n8946 ;
  assign n8948 = n8947 ^ n8944 ;
  assign n8949 = x6 & ~n409 ;
  assign n8950 = n207 & n6734 ;
  assign n8951 = x0 & n8950 ;
  assign n8952 = ~n8949 & n8951 ;
  assign n8953 = ~x0 & n8673 ;
  assign n8954 = n1255 & n8953 ;
  assign n8955 = n222 & n6866 ;
  assign n8956 = n7666 & n8955 ;
  assign n8957 = ~n8954 & ~n8956 ;
  assign n8958 = ~n8952 & n8957 ;
  assign n8959 = n8944 & n8958 ;
  assign n8960 = n8959 ^ n8862 ;
  assign n8961 = n8948 & n8960 ;
  assign n8962 = n8961 ^ n8959 ;
  assign n8963 = n8862 & n8962 ;
  assign n8964 = n8963 ^ n8947 ;
  assign n8965 = n8964 ^ x13 ;
  assign n8966 = n8965 ^ n8944 ;
  assign n8967 = n8861 & ~n8966 ;
  assign n8968 = ~n3441 & ~n5851 ;
  assign n8969 = ~x8 & n2168 ;
  assign n8970 = ~n2707 & ~n8969 ;
  assign n8971 = ~n1582 & ~n8970 ;
  assign n8972 = ~n1322 & n8971 ;
  assign n8973 = ~x9 & n38 ;
  assign n8974 = n1642 & n8973 ;
  assign n8975 = ~n8972 & ~n8974 ;
  assign n8976 = ~n43 & ~n8975 ;
  assign n8977 = n1365 & n2483 ;
  assign n8978 = n1260 & n5919 ;
  assign n8979 = ~n8977 & ~n8978 ;
  assign n8980 = n585 & ~n8979 ;
  assign n8981 = ~x12 & n2422 ;
  assign n8982 = ~n8980 & ~n8981 ;
  assign n8983 = n529 & n2904 ;
  assign n8984 = x13 & n603 ;
  assign n8985 = ~n8983 & ~n8984 ;
  assign n8986 = n1671 & ~n8985 ;
  assign n8987 = n1252 & n4713 ;
  assign n8988 = ~n8986 & ~n8987 ;
  assign n8989 = n8982 & n8988 ;
  assign n8990 = ~n8976 & n8989 ;
  assign n8991 = n1320 & ~n8990 ;
  assign n8992 = n49 & n98 ;
  assign n8993 = n1404 & n8992 ;
  assign n8994 = ~n133 & n1252 ;
  assign n8995 = n1608 & n2904 ;
  assign n8996 = n86 & n8995 ;
  assign n8997 = ~n8994 & ~n8996 ;
  assign n8998 = ~n1386 & n8997 ;
  assign n8999 = n1312 & ~n8998 ;
  assign n9000 = ~n1528 & ~n2739 ;
  assign n9001 = n1267 & n9000 ;
  assign n9002 = ~n6866 & ~n9001 ;
  assign n9003 = n8983 & ~n9002 ;
  assign n9004 = n1503 & n8973 ;
  assign n9005 = ~n9003 & ~n9004 ;
  assign n9006 = ~n8999 & n9005 ;
  assign n9007 = ~x4 & ~n9006 ;
  assign n9008 = n98 & n4536 ;
  assign n9009 = ~x12 & n9008 ;
  assign n9010 = ~n9007 & ~n9009 ;
  assign n9011 = ~n8993 & n9010 ;
  assign n9012 = ~n8991 & n9011 ;
  assign n9013 = n132 & ~n9012 ;
  assign n9014 = n1492 & n2156 ;
  assign n9015 = n8992 & n9014 ;
  assign n9016 = n153 & n5681 ;
  assign n9017 = n71 & n9016 ;
  assign n9018 = n222 & n4690 ;
  assign n9019 = ~x13 & n190 ;
  assign n9020 = ~n1322 & n9019 ;
  assign n9021 = n1581 & n9020 ;
  assign n9022 = ~n9018 & ~n9021 ;
  assign n9023 = ~n9017 & n9022 ;
  assign n9024 = n257 & ~n9023 ;
  assign n9025 = n49 & n1669 ;
  assign n9026 = ~n395 & ~n9025 ;
  assign n9027 = n264 & ~n9026 ;
  assign n9028 = n167 & n7595 ;
  assign n9029 = x7 & n2483 ;
  assign n9030 = ~n2197 & n9029 ;
  assign n9031 = n1376 & n2500 ;
  assign n9032 = ~n9030 & ~n9031 ;
  assign n9033 = ~n9028 & n9032 ;
  assign n9034 = ~n9027 & n9033 ;
  assign n9035 = n104 & ~n9034 ;
  assign n9036 = ~n9024 & ~n9035 ;
  assign n9037 = ~n9015 & n9036 ;
  assign n9038 = ~n9013 & n9037 ;
  assign n9039 = n1952 & ~n9038 ;
  assign n9040 = n655 & n1671 ;
  assign n9041 = n58 & n1669 ;
  assign n9042 = ~n9040 & ~n9041 ;
  assign n9043 = n264 & ~n9042 ;
  assign n9044 = n6481 & n9043 ;
  assign n9045 = ~x13 & ~n919 ;
  assign n9046 = n1630 & n9045 ;
  assign n9047 = ~n1511 & ~n5344 ;
  assign n9048 = ~n133 & ~n2233 ;
  assign n9049 = ~n9047 & n9048 ;
  assign n9050 = ~n9046 & ~n9049 ;
  assign n9051 = n20 & n307 ;
  assign n9052 = ~x10 & n9051 ;
  assign n9053 = ~n9050 & n9052 ;
  assign n9054 = n38 & n104 ;
  assign n9055 = n17 & n2483 ;
  assign n9056 = n9054 & n9055 ;
  assign n9057 = n6358 & n6824 ;
  assign n9058 = n280 & n1991 ;
  assign n9059 = n1642 & n9058 ;
  assign n9060 = ~n9057 & ~n9059 ;
  assign n9061 = x0 & ~n9060 ;
  assign n9062 = ~n9056 & ~n9061 ;
  assign n9063 = ~n9053 & n9062 ;
  assign n9064 = n98 & ~n9063 ;
  assign n9065 = x1 & ~n9064 ;
  assign n9066 = ~n9044 & n9065 ;
  assign n9067 = ~x5 & n1758 ;
  assign n9068 = n6248 & n9067 ;
  assign n9069 = n160 & n9068 ;
  assign n9070 = n22 & n140 ;
  assign n9071 = n86 & n9070 ;
  assign n9072 = ~n25 & ~n9071 ;
  assign n9073 = n2483 & ~n9072 ;
  assign n9074 = n9073 ^ x8 ;
  assign n9075 = ~n409 & ~n470 ;
  assign n9076 = ~x13 & n9075 ;
  assign n9077 = ~x12 & ~n9076 ;
  assign n9078 = n2181 & ~n9077 ;
  assign n9079 = ~n257 & ~n9078 ;
  assign n9080 = n9079 ^ x5 ;
  assign n9081 = n9080 ^ n9079 ;
  assign n9082 = n2105 & ~n9077 ;
  assign n9083 = n135 ^ x13 ;
  assign n9084 = n9083 ^ n135 ;
  assign n9085 = n9075 ^ n135 ;
  assign n9086 = n9085 ^ n135 ;
  assign n9087 = n9084 & n9086 ;
  assign n9088 = n9087 ^ n135 ;
  assign n9089 = ~x12 & n9088 ;
  assign n9090 = n9089 ^ n135 ;
  assign n9091 = n2181 & n9090 ;
  assign n9092 = n277 & ~n470 ;
  assign n9093 = ~n528 & ~n2233 ;
  assign n9094 = ~x12 & n9093 ;
  assign n9095 = ~n9092 & ~n9094 ;
  assign n9096 = n257 & ~n9095 ;
  assign n9097 = ~n9091 & ~n9096 ;
  assign n9098 = ~n9082 & n9097 ;
  assign n9099 = n9098 ^ n9079 ;
  assign n9100 = ~n9081 & n9099 ;
  assign n9101 = n9100 ^ n9079 ;
  assign n9102 = n9101 ^ n9073 ;
  assign n9103 = n9074 & n9102 ;
  assign n9104 = n9103 ^ n9100 ;
  assign n9105 = n9104 ^ n9079 ;
  assign n9106 = n9105 ^ x8 ;
  assign n9107 = ~n9073 & n9106 ;
  assign n9108 = n9107 ^ n9073 ;
  assign n9109 = n9108 ^ n9073 ;
  assign n9110 = ~x10 & ~n9109 ;
  assign n9111 = n425 & n1231 ;
  assign n9112 = ~x5 & n2904 ;
  assign n9113 = ~n503 & ~n6930 ;
  assign n9114 = n9112 & ~n9113 ;
  assign n9115 = ~x12 & n281 ;
  assign n9116 = n1254 & n9115 ;
  assign n9117 = ~n2439 & n5299 ;
  assign n9118 = ~n9116 & ~n9117 ;
  assign n9119 = ~n9114 & n9118 ;
  assign n9120 = n9119 ^ x7 ;
  assign n9121 = n9120 ^ n9119 ;
  assign n9122 = n9121 ^ n9111 ;
  assign n9123 = n2483 ^ x5 ;
  assign n9124 = ~n2483 & ~n9123 ;
  assign n9125 = n9124 ^ n9119 ;
  assign n9126 = n9125 ^ n2483 ;
  assign n9127 = ~n9122 & n9126 ;
  assign n9128 = n9127 ^ n9124 ;
  assign n9129 = n9128 ^ n2483 ;
  assign n9130 = ~n9111 & ~n9129 ;
  assign n9131 = n9130 ^ n9111 ;
  assign n9132 = n2225 & n9131 ;
  assign n9133 = n475 & n551 ;
  assign n9134 = ~n399 & ~n7955 ;
  assign n9135 = n9133 & n9134 ;
  assign n9136 = ~n135 & ~n5465 ;
  assign n9137 = x13 & ~n257 ;
  assign n9138 = ~n9136 & n9137 ;
  assign n9139 = ~n9135 & ~n9138 ;
  assign n9140 = n8186 & ~n9139 ;
  assign n9141 = n1138 & n1598 ;
  assign n9142 = ~x15 & ~n674 ;
  assign n9143 = n9141 & ~n9142 ;
  assign n9144 = n8002 & n9143 ;
  assign n9145 = n1415 & n2174 ;
  assign n9146 = n343 & n9145 ;
  assign n9147 = ~n9144 & ~n9146 ;
  assign n9148 = x6 & ~n9147 ;
  assign n9149 = ~n9140 & ~n9148 ;
  assign n9150 = ~n9132 & n9149 ;
  assign n9151 = ~n9110 & n9150 ;
  assign n9152 = ~n9069 & n9151 ;
  assign n9153 = n3896 & ~n9152 ;
  assign n9154 = n9066 & ~n9153 ;
  assign n9458 = n434 & n2659 ;
  assign n9459 = n1303 & n9458 ;
  assign n9460 = x15 & n3565 ;
  assign n9461 = ~x10 & ~n9460 ;
  assign n9155 = ~x13 & n1588 ;
  assign n9462 = ~n49 & ~n9155 ;
  assign n9463 = n551 & ~n9462 ;
  assign n9464 = ~n9461 & n9463 ;
  assign n9291 = n167 & n475 ;
  assign n9465 = n701 & n9291 ;
  assign n9466 = ~x9 & ~n8854 ;
  assign n9467 = ~n9067 & ~n9466 ;
  assign n9468 = ~n9465 & n9467 ;
  assign n9469 = ~n9464 & n9468 ;
  assign n9470 = n3643 & ~n9469 ;
  assign n9471 = ~n504 & n5353 ;
  assign n9472 = n1231 ^ x10 ;
  assign n9473 = n9472 ^ n9471 ;
  assign n9474 = n431 ^ x13 ;
  assign n9475 = ~n1231 & n9474 ;
  assign n9476 = n9475 ^ x13 ;
  assign n9477 = n9473 & ~n9476 ;
  assign n9478 = n9477 ^ n9475 ;
  assign n9479 = n9478 ^ x13 ;
  assign n9480 = n9479 ^ n1231 ;
  assign n9481 = ~n9471 & n9480 ;
  assign n9482 = x8 & ~n9481 ;
  assign n9483 = n200 & n1708 ;
  assign n9484 = n2904 & n9483 ;
  assign n9485 = n43 ^ x10 ;
  assign n9486 = n43 ^ x13 ;
  assign n9487 = n9486 ^ x13 ;
  assign n9488 = ~x5 & ~n2169 ;
  assign n9489 = n9488 ^ x13 ;
  assign n9490 = ~n9487 & ~n9489 ;
  assign n9491 = n9490 ^ x13 ;
  assign n9492 = n9485 & ~n9491 ;
  assign n9493 = n9492 ^ x10 ;
  assign n9494 = ~n9484 & n9493 ;
  assign n9495 = n1394 & ~n9494 ;
  assign n9496 = ~n2342 & ~n9495 ;
  assign n9497 = ~n9482 & n9496 ;
  assign n9498 = ~n1562 & ~n9497 ;
  assign n9499 = ~n2256 & n9498 ;
  assign n9500 = ~n9470 & ~n9499 ;
  assign n9501 = n9500 ^ x7 ;
  assign n9502 = n9501 ^ n9500 ;
  assign n9503 = ~x13 & n1394 ;
  assign n9504 = n294 & n3969 ;
  assign n9505 = ~n9503 & ~n9504 ;
  assign n9506 = n1502 & ~n9505 ;
  assign n9507 = ~n1257 & n7886 ;
  assign n9508 = n1138 & ~n9507 ;
  assign n9509 = n529 & n9000 ;
  assign n9510 = n1332 & n9509 ;
  assign n9511 = ~n9508 & ~n9510 ;
  assign n9512 = ~x0 & ~n9511 ;
  assign n9513 = ~n9506 & ~n9512 ;
  assign n9514 = n2904 & ~n9513 ;
  assign n9515 = n1551 & n3406 ;
  assign n9516 = ~n3865 & ~n9515 ;
  assign n9517 = n768 & ~n9516 ;
  assign n9518 = x14 & ~n3658 ;
  assign n9519 = n19 & n9518 ;
  assign n9520 = ~x14 & n3095 ;
  assign n9521 = n1394 ^ n434 ;
  assign n9522 = x10 & n9521 ;
  assign n9523 = n9522 ^ n1394 ;
  assign n9524 = ~n9520 & ~n9523 ;
  assign n9525 = ~n9519 & n9524 ;
  assign n9526 = n470 & n8853 ;
  assign n9527 = ~n190 & n1415 ;
  assign n9528 = x8 & ~n200 ;
  assign n9529 = ~n9527 & ~n9528 ;
  assign n9530 = ~n9526 & n9529 ;
  assign n9531 = n692 & n9530 ;
  assign n9532 = n9525 & n9531 ;
  assign n9533 = n475 & n2331 ;
  assign n9534 = n642 & n9533 ;
  assign n9535 = x8 & n9534 ;
  assign n9536 = ~n9532 & ~n9535 ;
  assign n9537 = ~n9517 & n9536 ;
  assign n9538 = ~n9514 & n9537 ;
  assign n9539 = n9538 ^ n9500 ;
  assign n9540 = ~n9502 & n9539 ;
  assign n9541 = n9540 ^ n9500 ;
  assign n9542 = ~n9459 & n9541 ;
  assign n9543 = ~x6 & ~n9542 ;
  assign n9544 = n429 & n3065 ;
  assign n9545 = n1290 & n9544 ;
  assign n9546 = x12 & n1252 ;
  assign n9547 = n3552 & n9546 ;
  assign n9548 = ~n2158 & ~n9547 ;
  assign n9549 = ~n43 & ~n9548 ;
  assign n9550 = x10 & x15 ;
  assign n9551 = ~n603 & ~n2708 ;
  assign n9552 = n9550 & n9551 ;
  assign n9553 = ~n9549 & ~n9552 ;
  assign n9554 = n429 & ~n9553 ;
  assign n9555 = ~x10 & n1366 ;
  assign n9556 = n3969 & n9555 ;
  assign n9557 = ~n1708 & ~n2677 ;
  assign n9558 = n2168 & n9557 ;
  assign n9559 = ~n3046 & ~n9558 ;
  assign n9560 = n1657 & ~n9559 ;
  assign n9561 = ~n1394 & n8983 ;
  assign n9562 = ~n8994 & ~n9561 ;
  assign n9563 = n1733 & ~n9562 ;
  assign n9564 = ~n9560 & ~n9563 ;
  assign n9565 = ~x7 & ~n9564 ;
  assign n9566 = ~n9556 & ~n9565 ;
  assign n9567 = ~n9554 & n9566 ;
  assign n9568 = n1583 & ~n9567 ;
  assign n9569 = n1758 & n2139 ;
  assign n9570 = n132 & n9569 ;
  assign n9571 = ~n9568 & ~n9570 ;
  assign n9572 = ~n9545 & n9571 ;
  assign n9573 = ~n9543 & n9572 ;
  assign n9574 = x4 & ~n9573 ;
  assign n9575 = n18 & n2219 ;
  assign n9576 = n549 & n9575 ;
  assign n9160 = ~x13 & n343 ;
  assign n9577 = n1332 & n9160 ;
  assign n9578 = n291 & n6169 ;
  assign n9579 = n9577 & n9578 ;
  assign n9580 = n475 & n570 ;
  assign n9581 = n9580 ^ x4 ;
  assign n9582 = n9581 ^ x6 ;
  assign n9588 = n9582 ^ n9581 ;
  assign n9583 = n9582 ^ n9580 ;
  assign n9584 = n9583 ^ n4713 ;
  assign n9585 = n9582 ^ n4713 ;
  assign n9586 = n9585 ^ n9581 ;
  assign n9587 = n9584 & n9586 ;
  assign n9589 = n9588 ^ n9587 ;
  assign n9590 = ~n43 & ~n2169 ;
  assign n9199 = ~x9 & n475 ;
  assign n9591 = ~x14 & n9199 ;
  assign n9592 = ~n9590 & ~n9591 ;
  assign n9593 = x12 & ~n9592 ;
  assign n9594 = n9593 ^ n9582 ;
  assign n9595 = ~n9588 & n9594 ;
  assign n9596 = n9595 ^ n9593 ;
  assign n9597 = ~n9589 & n9596 ;
  assign n9598 = n9597 ^ n9587 ;
  assign n9599 = n9598 ^ n9582 ;
  assign n9600 = n9599 ^ x4 ;
  assign n9601 = n9600 ^ n9581 ;
  assign n9602 = n429 & n9601 ;
  assign n9603 = n1597 & n9602 ;
  assign n9604 = ~n9579 & ~n9603 ;
  assign n9605 = x8 & ~n9604 ;
  assign n9606 = n5092 & n7042 ;
  assign n9156 = ~x7 & n9155 ;
  assign n9607 = n267 & n9156 ;
  assign n9608 = ~n153 & n1273 ;
  assign n9609 = ~n9607 & ~n9608 ;
  assign n9610 = ~n9606 & n9609 ;
  assign n9611 = n642 & ~n9610 ;
  assign n9612 = n2469 & n6169 ;
  assign n9613 = ~n269 & n721 ;
  assign n9614 = n9613 ^ x12 ;
  assign n9615 = n9614 ^ n9112 ;
  assign n9616 = n6564 ^ x6 ;
  assign n9617 = n9616 ^ n9614 ;
  assign n9618 = ~n9613 & ~n9617 ;
  assign n9619 = n9618 ^ x6 ;
  assign n9620 = n9619 ^ n9613 ;
  assign n9621 = n9620 ^ n9614 ;
  assign n9622 = n9621 ^ n9112 ;
  assign n9623 = n9615 & n9622 ;
  assign n9624 = n9623 ^ n9618 ;
  assign n9625 = n9624 ^ x6 ;
  assign n9626 = n9625 ^ n9614 ;
  assign n9627 = n9112 & ~n9626 ;
  assign n9628 = n9627 ^ n9112 ;
  assign n9629 = n9628 ^ n9112 ;
  assign n9630 = ~n9612 & ~n9629 ;
  assign n9631 = ~n9611 & n9630 ;
  assign n9632 = n3294 & ~n9631 ;
  assign n9359 = ~x5 & n1276 ;
  assign n9633 = n603 & n768 ;
  assign n9634 = n9359 & n9633 ;
  assign n9397 = ~n2105 & ~n2483 ;
  assign n9635 = ~x13 & ~n2126 ;
  assign n9636 = ~n504 & n9635 ;
  assign n9637 = n9397 & ~n9636 ;
  assign n9638 = n3294 & ~n9637 ;
  assign n9639 = ~n2182 & n7980 ;
  assign n9640 = ~n9638 & ~n9639 ;
  assign n9641 = n25 & ~n9640 ;
  assign n9642 = ~n9634 & ~n9641 ;
  assign n9643 = ~n9632 & n9642 ;
  assign n9644 = n17 & ~n9643 ;
  assign n9645 = ~n9605 & ~n9644 ;
  assign n9646 = ~n9576 & n9645 ;
  assign n9647 = ~n9574 & n9646 ;
  assign n9157 = ~n121 & ~n9156 ;
  assign n9158 = n9157 ^ x7 ;
  assign n9159 = n9158 ^ n9157 ;
  assign n9161 = n9160 ^ n9157 ;
  assign n9162 = n9161 ^ n9157 ;
  assign n9163 = ~n9159 & n9162 ;
  assign n9164 = n9163 ^ n9157 ;
  assign n9165 = ~x4 & ~n9164 ;
  assign n9166 = n9165 ^ n9157 ;
  assign n9167 = n2516 & ~n9166 ;
  assign n9168 = ~x6 & n61 ;
  assign n9169 = ~n588 & n1124 ;
  assign n9170 = n9168 & n9169 ;
  assign n9171 = ~x7 & n3068 ;
  assign n9172 = n5054 & n9171 ;
  assign n9173 = n475 & n9172 ;
  assign n9174 = ~n9170 & ~n9173 ;
  assign n9175 = n1073 & n6204 ;
  assign n9176 = n334 & n9175 ;
  assign n9177 = n9174 & ~n9176 ;
  assign n9178 = ~n9167 & n9177 ;
  assign n9179 = n9178 ^ x10 ;
  assign n9180 = n42 & n167 ;
  assign n9181 = ~n561 & ~n9180 ;
  assign n9182 = n684 & ~n9181 ;
  assign n9184 = n160 & n7177 ;
  assign n9185 = ~n166 & ~n9184 ;
  assign n9183 = n62 & n592 ;
  assign n9186 = n9185 ^ n9183 ;
  assign n9187 = n9186 ^ n9185 ;
  assign n9188 = n9185 ^ x13 ;
  assign n9189 = n9188 ^ n9185 ;
  assign n9190 = n9187 & n9189 ;
  assign n9191 = n9190 ^ n9185 ;
  assign n9192 = ~x9 & ~n9191 ;
  assign n9193 = n9192 ^ n9185 ;
  assign n9194 = ~n9182 & n9193 ;
  assign n9195 = n252 & ~n9194 ;
  assign n9196 = n431 & n9168 ;
  assign n9197 = n591 & n9196 ;
  assign n9198 = ~n9195 & ~n9197 ;
  assign n9200 = ~x0 & n1290 ;
  assign n9201 = n9199 & n9200 ;
  assign n9202 = n608 & n9201 ;
  assign n9203 = n9202 ^ n9198 ;
  assign n9204 = ~x13 & n731 ;
  assign n9205 = ~n865 & ~n9204 ;
  assign n9206 = n101 & ~n9205 ;
  assign n9207 = n429 & n8984 ;
  assign n9208 = ~n9206 & ~n9207 ;
  assign n9209 = ~x6 & n752 ;
  assign n9210 = ~n9208 & n9209 ;
  assign n9211 = n549 & n5299 ;
  assign n9212 = n153 & n9211 ;
  assign n9213 = ~n9210 & ~n9212 ;
  assign n9214 = ~n470 & ~n9213 ;
  assign n9215 = n49 & n718 ;
  assign n9216 = n190 ^ x0 ;
  assign n9217 = n190 ^ x12 ;
  assign n9218 = n9217 ^ x12 ;
  assign n9219 = x5 & ~n504 ;
  assign n9220 = n9219 ^ x12 ;
  assign n9221 = ~n9218 & n9220 ;
  assign n9222 = n9221 ^ x12 ;
  assign n9223 = ~n9216 & ~n9222 ;
  assign n9224 = n9223 ^ x0 ;
  assign n9225 = n721 & ~n9224 ;
  assign n9226 = ~n476 & n1175 ;
  assign n9227 = n684 & n1454 ;
  assign n9228 = ~n9054 & ~n9227 ;
  assign n9229 = ~n166 & n9228 ;
  assign n9230 = ~n9226 & n9229 ;
  assign n9231 = ~n9225 & n9230 ;
  assign n9232 = ~x9 & ~n9231 ;
  assign n9233 = x7 & n2342 ;
  assign n9234 = ~n320 & n642 ;
  assign n9235 = ~n61 & ~n9234 ;
  assign n9236 = n586 & ~n9235 ;
  assign n9237 = ~n9233 & ~n9236 ;
  assign n9238 = ~n9232 & n9237 ;
  assign n9239 = ~n9215 & n9238 ;
  assign n9240 = n9239 ^ x6 ;
  assign n9241 = n9240 ^ n9239 ;
  assign n9242 = n9241 ^ n9214 ;
  assign n9243 = n166 & ~n476 ;
  assign n9244 = n5149 & n7177 ;
  assign n9245 = ~n9243 & ~n9244 ;
  assign n9246 = n9245 ^ n570 ;
  assign n9247 = ~n9245 & ~n9246 ;
  assign n9248 = n9247 ^ n9239 ;
  assign n9249 = n9248 ^ n9245 ;
  assign n9250 = n9242 & n9249 ;
  assign n9251 = n9250 ^ n9247 ;
  assign n9252 = n9251 ^ n9245 ;
  assign n9253 = ~n9214 & ~n9252 ;
  assign n9254 = n9253 ^ n9214 ;
  assign n9255 = n9254 ^ x4 ;
  assign n9256 = n9255 ^ n9254 ;
  assign n9257 = ~n284 & n2904 ;
  assign n9258 = ~n49 & ~n9257 ;
  assign n9259 = n684 & ~n9258 ;
  assign n9260 = n1154 & n9204 ;
  assign n9261 = ~n1886 & ~n9260 ;
  assign n9262 = n2904 & ~n9261 ;
  assign n9263 = n1138 & ~n6616 ;
  assign n9264 = ~n5843 & ~n9263 ;
  assign n9265 = ~n504 & ~n9264 ;
  assign n9266 = n4845 & n6554 ;
  assign n9267 = ~n9265 & ~n9266 ;
  assign n9268 = ~n1208 & n9267 ;
  assign n9269 = ~n9262 & n9268 ;
  assign n9270 = n9269 ^ n2235 ;
  assign n9271 = n9270 ^ x0 ;
  assign n9278 = n9271 ^ n9270 ;
  assign n9272 = n9271 ^ n9233 ;
  assign n9273 = n9272 ^ n9270 ;
  assign n9274 = n9271 ^ n9269 ;
  assign n9275 = n9274 ^ n9233 ;
  assign n9276 = n9275 ^ n9273 ;
  assign n9277 = n9273 & n9276 ;
  assign n9279 = n9278 ^ n9277 ;
  assign n9280 = n9279 ^ n9273 ;
  assign n9281 = n9270 ^ n551 ;
  assign n9282 = n9277 ^ n9273 ;
  assign n9283 = ~n9281 & n9282 ;
  assign n9284 = n9283 ^ n9270 ;
  assign n9285 = ~n9280 & n9284 ;
  assign n9286 = n9285 ^ n9270 ;
  assign n9287 = n9286 ^ n2235 ;
  assign n9288 = n9287 ^ n9270 ;
  assign n9289 = ~n9259 & n9288 ;
  assign n9290 = ~x6 & ~n9289 ;
  assign n9292 = n718 & n9291 ;
  assign n9293 = ~n9290 & ~n9292 ;
  assign n9294 = n9293 ^ n9254 ;
  assign n9295 = n9256 & ~n9294 ;
  assign n9296 = n9295 ^ n9254 ;
  assign n9297 = n9296 ^ n9198 ;
  assign n9298 = ~n9203 & ~n9297 ;
  assign n9299 = n9298 ^ n9295 ;
  assign n9300 = n9299 ^ n9254 ;
  assign n9301 = n9300 ^ n9202 ;
  assign n9302 = n9198 & n9301 ;
  assign n9303 = n9302 ^ n9198 ;
  assign n9304 = n9303 ^ x8 ;
  assign n9305 = n9304 ^ n9303 ;
  assign n9306 = n1583 & n2904 ;
  assign n9307 = n7293 & n9306 ;
  assign n9308 = n133 & n9307 ;
  assign n9309 = n1397 ^ n42 ;
  assign n9310 = n9309 ^ n1366 ;
  assign n9311 = n9310 ^ n1397 ;
  assign n9312 = n9311 ^ n9310 ;
  assign n9313 = ~n2169 & n5124 ;
  assign n9314 = n9313 ^ n9310 ;
  assign n9315 = n9314 ^ n9309 ;
  assign n9316 = n9312 & ~n9315 ;
  assign n9317 = n9316 ^ n9313 ;
  assign n9318 = ~n1902 & ~n9313 ;
  assign n9319 = n9318 ^ n9309 ;
  assign n9320 = ~n9317 & ~n9319 ;
  assign n9321 = n9320 ^ n9318 ;
  assign n9322 = ~n9309 & n9321 ;
  assign n9323 = n9322 ^ n9316 ;
  assign n9324 = n9323 ^ n42 ;
  assign n9325 = n9324 ^ n9313 ;
  assign n9326 = n586 & ~n9325 ;
  assign n9327 = ~x4 & n2105 ;
  assign n9328 = n640 & n9327 ;
  assign n9329 = n52 & ~n1434 ;
  assign n9330 = n217 & n5408 ;
  assign n9331 = ~n9329 & ~n9330 ;
  assign n9332 = ~n9328 & n9331 ;
  assign n9333 = n9160 & ~n9332 ;
  assign n9334 = x6 ^ x5 ;
  assign n9335 = n2904 ^ x6 ;
  assign n9336 = n9335 ^ n2904 ;
  assign n9337 = ~x9 & n343 ;
  assign n9338 = ~n3068 & ~n9337 ;
  assign n9339 = n9338 ^ n2904 ;
  assign n9340 = n9336 & ~n9339 ;
  assign n9341 = n9340 ^ n2904 ;
  assign n9342 = ~n9334 & n9341 ;
  assign n9343 = n721 & n9342 ;
  assign n9344 = n867 & n2483 ;
  assign n9345 = n277 & n6358 ;
  assign n9346 = ~n9344 & ~n9345 ;
  assign n9347 = ~n9343 & n9346 ;
  assign n9348 = ~x4 & ~n9347 ;
  assign n9349 = n5156 & n7826 ;
  assign n9350 = ~n4645 & ~n9171 ;
  assign n9351 = n1123 & ~n1267 ;
  assign n9352 = ~n9350 & n9351 ;
  assign n9353 = ~n9349 & ~n9352 ;
  assign n9354 = n252 & n3068 ;
  assign n9355 = n22 & n9354 ;
  assign n9356 = n42 & n9355 ;
  assign n9357 = n9353 & ~n9356 ;
  assign n9358 = ~n476 & ~n9357 ;
  assign n9360 = n119 & n9359 ;
  assign n9361 = ~n9338 & n9360 ;
  assign n9362 = n2585 ^ n25 ;
  assign n9363 = x13 & n9183 ;
  assign n9364 = n9363 ^ n2585 ;
  assign n9365 = n9364 ^ n9363 ;
  assign n9366 = n9365 ^ n9362 ;
  assign n9367 = n6923 ^ x9 ;
  assign n9368 = ~x9 & ~n9367 ;
  assign n9369 = n9368 ^ n9363 ;
  assign n9370 = n9369 ^ x9 ;
  assign n9371 = ~n9366 & n9370 ;
  assign n9372 = n9371 ^ n9368 ;
  assign n9373 = n9372 ^ x9 ;
  assign n9374 = n9362 & ~n9373 ;
  assign n9375 = n9374 ^ n2585 ;
  assign n9376 = ~n9361 & ~n9375 ;
  assign n9377 = ~n9358 & n9376 ;
  assign n9378 = ~n9348 & n9377 ;
  assign n9379 = ~n9333 & n9378 ;
  assign n9380 = n9379 ^ x0 ;
  assign n9381 = n9380 ^ n9379 ;
  assign n9382 = ~n284 & n608 ;
  assign n9383 = n190 & n9382 ;
  assign n9384 = n25 & n9160 ;
  assign n9385 = ~n865 & ~n9384 ;
  assign n9386 = ~n9383 & n9385 ;
  assign n9387 = n4327 & ~n9386 ;
  assign n9388 = n62 & ~n214 ;
  assign n9389 = ~x9 & ~n49 ;
  assign n9390 = ~n1230 & ~n1254 ;
  assign n9391 = ~n249 & ~n9390 ;
  assign n9392 = ~n9389 & n9391 ;
  assign n9393 = ~n9388 & n9392 ;
  assign n9394 = ~n9387 & ~n9393 ;
  assign n9395 = x12 & ~n2169 ;
  assign n9396 = n2118 & n9395 ;
  assign n9398 = n608 & ~n9397 ;
  assign n9399 = ~n9396 & ~n9398 ;
  assign n9400 = n963 & ~n9399 ;
  assign n9401 = n25 & n2181 ;
  assign n9402 = ~x13 & n1492 ;
  assign n9403 = n570 & n9402 ;
  assign n9404 = ~x14 & n9403 ;
  assign n9405 = ~n9401 & ~n9404 ;
  assign n9406 = ~x13 & ~n42 ;
  assign n9407 = n591 & ~n9406 ;
  assign n9408 = ~n257 & ~n570 ;
  assign n9409 = ~n9407 & ~n9408 ;
  assign n9410 = n1492 & ~n9409 ;
  assign n9411 = n2174 & n2469 ;
  assign n9412 = ~x14 & n2174 ;
  assign n9413 = n1260 & n9412 ;
  assign n9414 = ~n9411 & ~n9413 ;
  assign n9415 = ~n9410 & n9414 ;
  assign n9416 = n9405 & n9415 ;
  assign n9417 = ~n9400 & n9416 ;
  assign n9418 = n9417 ^ x4 ;
  assign n9419 = n9418 ^ n9417 ;
  assign n9420 = n9419 ^ n9394 ;
  assign n9421 = x5 & ~n2169 ;
  assign n9422 = ~x7 & n1607 ;
  assign n9423 = n9421 & n9422 ;
  assign n9424 = n264 & ~n3453 ;
  assign n9425 = n167 & n592 ;
  assign n9426 = x14 & n9425 ;
  assign n9427 = ~n9424 & ~n9426 ;
  assign n9428 = n434 & n1454 ;
  assign n9429 = x7 & n9428 ;
  assign n9430 = ~n9233 & ~n9429 ;
  assign n9431 = n9427 & n9430 ;
  assign n9432 = ~n9423 & n9431 ;
  assign n9433 = n9432 ^ x6 ;
  assign n9434 = ~n9432 & ~n9433 ;
  assign n9435 = n9434 ^ n9417 ;
  assign n9436 = n9435 ^ n9432 ;
  assign n9437 = ~n9420 & n9436 ;
  assign n9438 = n9437 ^ n9434 ;
  assign n9439 = n9438 ^ n9432 ;
  assign n9440 = n9394 & ~n9439 ;
  assign n9441 = n9440 ^ n9394 ;
  assign n9442 = n9441 ^ n9379 ;
  assign n9443 = n9381 & n9442 ;
  assign n9444 = n9443 ^ n9379 ;
  assign n9445 = ~n9326 & n9444 ;
  assign n9446 = ~n9308 & n9445 ;
  assign n9447 = n9446 ^ n9303 ;
  assign n9448 = n9305 & n9447 ;
  assign n9449 = n9448 ^ n9303 ;
  assign n9450 = n9449 ^ n9178 ;
  assign n9451 = n9179 & n9450 ;
  assign n9452 = n9451 ^ n9448 ;
  assign n9453 = n9452 ^ n9303 ;
  assign n9454 = n9453 ^ x10 ;
  assign n9455 = n9178 & n9454 ;
  assign n9456 = n9455 ^ n9178 ;
  assign n9457 = n9456 ^ x10 ;
  assign n9648 = n9647 ^ n9457 ;
  assign n9649 = n9648 ^ n9647 ;
  assign n9650 = ~n1365 & ~n1667 ;
  assign n9651 = n1886 & n9650 ;
  assign n9652 = n5344 & n7045 ;
  assign n9653 = ~n9651 & ~n9652 ;
  assign n9654 = n1376 & ~n9653 ;
  assign n9655 = n86 & n1669 ;
  assign n9656 = ~n1547 & ~n9655 ;
  assign n9657 = n1886 & ~n9656 ;
  assign n9658 = n1698 & n6564 ;
  assign n9659 = n6362 & n9658 ;
  assign n9660 = n1945 & n9503 ;
  assign n9661 = ~n9659 & ~n9660 ;
  assign n9662 = ~n9657 & n9661 ;
  assign n9663 = n9662 ^ n399 ;
  assign n9664 = n9663 ^ n9662 ;
  assign n9665 = n1214 & n2103 ;
  assign n9666 = ~n1529 & n9402 ;
  assign n9667 = ~n9665 & ~n9666 ;
  assign n9668 = n9667 ^ n9662 ;
  assign n9669 = n9668 ^ n9662 ;
  assign n9670 = n9664 & ~n9669 ;
  assign n9671 = n9670 ^ n9662 ;
  assign n9672 = x4 & ~n9671 ;
  assign n9673 = n9672 ^ n9662 ;
  assign n9674 = ~n9654 & n9673 ;
  assign n9675 = n2904 & ~n9674 ;
  assign n9676 = ~n8172 & ~n9327 ;
  assign n9677 = n1208 & ~n9676 ;
  assign n9678 = ~n1352 & n8577 ;
  assign n9679 = ~n1078 & ~n4052 ;
  assign n9680 = ~n2309 & n9679 ;
  assign n9681 = n4713 & n9680 ;
  assign n9682 = ~n9678 & ~n9681 ;
  assign n9683 = n2174 & ~n9682 ;
  assign n9684 = x15 & n9683 ;
  assign n9685 = ~n9677 & ~n9684 ;
  assign n9686 = x5 & ~n9397 ;
  assign n9687 = ~n2227 & ~n9686 ;
  assign n9688 = n4052 & ~n9687 ;
  assign n9689 = n551 & n1644 ;
  assign n9690 = n1642 & n4737 ;
  assign n9691 = n865 & n9690 ;
  assign n9692 = ~n9689 & ~n9691 ;
  assign n9693 = ~n9688 & n9692 ;
  assign n9694 = x7 & ~n9693 ;
  assign n9695 = n291 & ~n738 ;
  assign n9696 = n394 & n646 ;
  assign n9697 = ~n1292 & ~n9696 ;
  assign n9698 = ~n9695 & n9697 ;
  assign n9699 = n1252 & ~n9698 ;
  assign n9700 = n394 & ~n2565 ;
  assign n9701 = ~n1261 & ~n9700 ;
  assign n9702 = ~x7 & ~n431 ;
  assign n9703 = n1550 & n9702 ;
  assign n9704 = ~n9701 & n9703 ;
  assign n9705 = x13 & n9008 ;
  assign n9706 = n250 & n4922 ;
  assign n9707 = n1902 & n9706 ;
  assign n9708 = ~n9705 & ~n9707 ;
  assign n9709 = ~n9704 & n9708 ;
  assign n9710 = ~n9699 & n9709 ;
  assign n9711 = ~x12 & ~n9710 ;
  assign n9712 = ~n9694 & ~n9711 ;
  assign n9713 = ~n52 & ~n9412 ;
  assign n9714 = n1581 & ~n9713 ;
  assign n9715 = n9714 ^ x8 ;
  assign n9716 = n1123 ^ x9 ;
  assign n9717 = n9716 ^ n1123 ;
  assign n9718 = ~n1266 & n1320 ;
  assign n9719 = ~n8920 & ~n9718 ;
  assign n9720 = n9719 ^ n1123 ;
  assign n9721 = n9717 & ~n9720 ;
  assign n9722 = n9721 ^ n1123 ;
  assign n9723 = n9722 ^ n9714 ;
  assign n9724 = n9715 & ~n9723 ;
  assign n9725 = n9724 ^ n9721 ;
  assign n9726 = n9725 ^ n1123 ;
  assign n9727 = n9726 ^ x8 ;
  assign n9728 = ~n9714 & ~n9727 ;
  assign n9729 = n9728 ^ n9714 ;
  assign n9730 = n9729 ^ n9714 ;
  assign n9731 = n4713 & ~n9730 ;
  assign n9732 = n9712 & ~n9731 ;
  assign n9733 = n9685 & n9732 ;
  assign n9734 = ~n9675 & n9733 ;
  assign n9735 = n1747 & ~n9734 ;
  assign n9736 = n549 & n4536 ;
  assign n9737 = n1123 & n9736 ;
  assign n9738 = x0 & ~n8352 ;
  assign n9739 = ~n4132 & ~n9738 ;
  assign n9740 = n2168 & ~n9739 ;
  assign n9741 = n294 & n7979 ;
  assign n9742 = ~n9740 & ~n9741 ;
  assign n9743 = n2308 & ~n9742 ;
  assign n9744 = n167 & n6564 ;
  assign n9745 = n5221 & n9744 ;
  assign n9746 = n244 & n1312 ;
  assign n9747 = n5465 & n9746 ;
  assign n9748 = n1457 & n9747 ;
  assign n9749 = ~n9745 & ~n9748 ;
  assign n9750 = ~n9743 & n9749 ;
  assign n9751 = n1633 & ~n9750 ;
  assign n9752 = n25 & n6139 ;
  assign n9753 = n1551 & n9752 ;
  assign n9754 = x9 & n9141 ;
  assign n9755 = x9 ^ x8 ;
  assign n9756 = n9755 ^ x8 ;
  assign n9757 = n9756 ^ n1502 ;
  assign n9758 = x12 & ~n475 ;
  assign n9759 = n4762 & ~n9758 ;
  assign n9760 = n9759 ^ n4753 ;
  assign n9761 = ~n9759 & n9760 ;
  assign n9762 = n9761 ^ x8 ;
  assign n9763 = n9762 ^ n9759 ;
  assign n9764 = ~n9757 & ~n9763 ;
  assign n9765 = n9764 ^ n9761 ;
  assign n9766 = n9765 ^ n9759 ;
  assign n9767 = n1502 & ~n9766 ;
  assign n9768 = n9767 ^ n1502 ;
  assign n9769 = ~n9754 & ~n9768 ;
  assign n9770 = n98 & ~n9769 ;
  assign n9771 = n22 & n1365 ;
  assign n9772 = n1548 & n9771 ;
  assign n9773 = x15 & n6013 ;
  assign n9774 = n9773 ^ n4573 ;
  assign n9775 = n9772 & n9774 ;
  assign n9776 = ~n9770 & ~n9775 ;
  assign n9777 = ~n9753 & n9776 ;
  assign n9778 = ~n3462 & ~n9777 ;
  assign n9779 = n551 & n6923 ;
  assign n9780 = n1073 & n2304 ;
  assign n9781 = n9779 & n9780 ;
  assign n9782 = ~n9778 & ~n9781 ;
  assign n9783 = ~n9751 & n9782 ;
  assign n9784 = ~n9737 & n9783 ;
  assign n9785 = ~n9735 & n9784 ;
  assign n9786 = n9785 ^ n9647 ;
  assign n9787 = n9786 ^ n9647 ;
  assign n9788 = ~n9649 & n9787 ;
  assign n9789 = n9788 ^ n9647 ;
  assign n9790 = x2 & n9789 ;
  assign n9791 = n9790 ^ n9647 ;
  assign n9792 = n9154 & n9791 ;
  assign n9793 = ~n9039 & n9792 ;
  assign n9794 = n3065 & n4941 ;
  assign n9795 = ~n167 & n4619 ;
  assign n9796 = n3018 & n9795 ;
  assign n9797 = ~n2006 & n9796 ;
  assign n9798 = ~n9794 & ~n9797 ;
  assign n9799 = n165 & ~n9798 ;
  assign n9800 = ~n717 & ~n1123 ;
  assign n9801 = ~n1622 & ~n9800 ;
  assign n9802 = n3454 & n9801 ;
  assign n9803 = x12 & n6481 ;
  assign n9804 = ~x14 & n9803 ;
  assign n9805 = ~n9802 & ~n9804 ;
  assign n9806 = ~n1716 & ~n9805 ;
  assign n9807 = x13 & n7387 ;
  assign n9808 = n9807 ^ n649 ;
  assign n9809 = n8389 & n9808 ;
  assign n9810 = ~n9806 & ~n9809 ;
  assign n9811 = n1503 & ~n9810 ;
  assign n9812 = ~n161 & ~n434 ;
  assign n9813 = n1520 & ~n9812 ;
  assign n9814 = n5345 & n9813 ;
  assign n9815 = x13 & n7726 ;
  assign n9816 = ~n9814 & ~n9815 ;
  assign n9817 = n210 & n1123 ;
  assign n9818 = n1534 & n9817 ;
  assign n9819 = ~n77 & n8598 ;
  assign n9820 = ~n104 & ~n3264 ;
  assign n9821 = n291 & n9820 ;
  assign n9822 = n9819 & n9821 ;
  assign n9823 = n38 & n3283 ;
  assign n9824 = n1332 & n5277 ;
  assign n9825 = n9823 & n9824 ;
  assign n9826 = ~n9822 & ~n9825 ;
  assign n9827 = ~n9818 & n9826 ;
  assign n9828 = n9816 & n9827 ;
  assign n9829 = ~n9811 & n9828 ;
  assign n9830 = n257 & ~n9829 ;
  assign n9831 = ~n9799 & ~n9830 ;
  assign n9832 = ~x9 & n4312 ;
  assign n9833 = ~n8188 & n9832 ;
  assign n9834 = ~x8 & n4561 ;
  assign n9835 = n20 & n2331 ;
  assign n9836 = n9834 & n9835 ;
  assign n9837 = n2387 & n8177 ;
  assign n9838 = ~n9836 & ~n9837 ;
  assign n9839 = ~n9833 & n9838 ;
  assign n9840 = n104 & ~n9839 ;
  assign n9841 = n3437 & n5940 ;
  assign n9842 = n3439 & n5961 ;
  assign n9843 = ~n9841 & ~n9842 ;
  assign n9844 = ~n6358 & ~n9421 ;
  assign n9845 = ~n9843 & ~n9844 ;
  assign n9846 = ~x1 & ~n9845 ;
  assign n9847 = n768 & n7884 ;
  assign n9848 = n2724 & n9847 ;
  assign n9849 = ~x4 & n6358 ;
  assign n9850 = n2556 & n9849 ;
  assign n9851 = n1256 & n9850 ;
  assign n9852 = ~n9848 & ~n9851 ;
  assign n9853 = n9846 & n9852 ;
  assign n9854 = ~n9840 & n9853 ;
  assign n9855 = n6401 & n6814 ;
  assign n9856 = n3981 & n4756 ;
  assign n9857 = n1670 & n3217 ;
  assign n9858 = ~n9856 & ~n9857 ;
  assign n9859 = ~n1716 & ~n9858 ;
  assign n9860 = n3267 & n5345 ;
  assign n9861 = ~n9859 & ~n9860 ;
  assign n9862 = ~n9855 & n9861 ;
  assign n9863 = n551 & n721 ;
  assign n9864 = ~n9862 & n9863 ;
  assign n9865 = n9854 & ~n9864 ;
  assign n9988 = n133 & n222 ;
  assign n9989 = ~n6093 & ~n9988 ;
  assign n9990 = ~n1716 & ~n9989 ;
  assign n9991 = n194 & n1702 ;
  assign n9992 = n210 & n6092 ;
  assign n9993 = ~n9991 & ~n9992 ;
  assign n9994 = n1330 & ~n9993 ;
  assign n9995 = ~n9990 & ~n9994 ;
  assign n9996 = n2422 & ~n9995 ;
  assign n9997 = n2309 & n2399 ;
  assign n9998 = n9817 & n9997 ;
  assign n9999 = ~n9996 & ~n9998 ;
  assign n10000 = n529 & n2397 ;
  assign n10001 = ~n609 & n5992 ;
  assign n10002 = ~n10000 & ~n10001 ;
  assign n10003 = x0 & ~n10002 ;
  assign n10004 = n1310 & n3452 ;
  assign n10005 = ~n292 & n3643 ;
  assign n10006 = ~n3508 & n10005 ;
  assign n10007 = n529 & n10006 ;
  assign n10008 = ~n10004 & ~n10007 ;
  assign n10009 = ~n10003 & n10008 ;
  assign n10010 = x9 & ~n10009 ;
  assign n10011 = ~x9 & ~n210 ;
  assign n10012 = ~n5564 & ~n10011 ;
  assign n10013 = n717 & ~n10012 ;
  assign n10014 = ~n3452 & n10013 ;
  assign n10015 = ~n10010 & ~n10014 ;
  assign n10016 = n5124 & ~n10015 ;
  assign n10047 = n228 & n4107 ;
  assign n10048 = ~n294 & n3060 ;
  assign n10049 = ~n8047 & n10048 ;
  assign n10050 = n4122 & n10000 ;
  assign n10051 = ~n10049 & ~n10050 ;
  assign n10052 = n291 & ~n10051 ;
  assign n10053 = ~n10047 & ~n10052 ;
  assign n10054 = n291 & n852 ;
  assign n10055 = ~n6909 & ~n10054 ;
  assign n10056 = ~n2278 & ~n10055 ;
  assign n10057 = n10053 & ~n10056 ;
  assign n10017 = ~n1511 & ~n9546 ;
  assign n10018 = n1826 & ~n10017 ;
  assign n10019 = n3068 & ~n6110 ;
  assign n10020 = n8745 & n10019 ;
  assign n10021 = x9 & n1698 ;
  assign n10022 = n3557 & n10021 ;
  assign n10023 = ~n10020 & ~n10022 ;
  assign n10024 = ~n10018 & n10023 ;
  assign n10025 = ~n1716 & ~n10024 ;
  assign n10026 = n529 & n1252 ;
  assign n10027 = ~n3808 & ~n10026 ;
  assign n10028 = ~n2916 & ~n10027 ;
  assign n10029 = ~n3848 & ~n3896 ;
  assign n10030 = n717 & n1252 ;
  assign n10031 = ~n10029 & n10030 ;
  assign n10032 = ~n10028 & ~n10031 ;
  assign n10033 = ~n10025 & n10032 ;
  assign n10058 = n10057 ^ n10033 ;
  assign n10034 = n1598 & n3980 ;
  assign n10035 = x8 & ~n1322 ;
  assign n10036 = ~n10034 & ~n10035 ;
  assign n10037 = ~n1716 & ~n10036 ;
  assign n10038 = ~n6815 & ~n10037 ;
  assign n10039 = ~x13 & ~n10038 ;
  assign n10040 = ~n134 & n394 ;
  assign n10041 = ~n7001 & ~n10040 ;
  assign n10042 = n2309 & ~n10041 ;
  assign n10043 = ~n1684 & ~n10042 ;
  assign n10044 = n210 & ~n10043 ;
  assign n10045 = ~n10039 & ~n10044 ;
  assign n10046 = n10045 ^ n10033 ;
  assign n10059 = n10058 ^ n10046 ;
  assign n10060 = n10046 ^ x9 ;
  assign n10061 = n10060 ^ n10046 ;
  assign n10062 = n10059 & ~n10061 ;
  assign n10063 = n10062 ^ n10046 ;
  assign n10064 = x5 & n10063 ;
  assign n10065 = n10064 ^ n10033 ;
  assign n10066 = ~n10016 & n10065 ;
  assign n10067 = n10066 ^ x10 ;
  assign n10068 = n10067 ^ n10066 ;
  assign n10069 = n10068 ^ n9999 ;
  assign n10070 = ~n249 & ~n1581 ;
  assign n10071 = ~n5919 & ~n10070 ;
  assign n10072 = ~n2585 & ~n10071 ;
  assign n10073 = n1248 & ~n10072 ;
  assign n10074 = ~n394 & ~n2710 ;
  assign n10075 = ~x2 & n9397 ;
  assign n10076 = n10074 & n10075 ;
  assign n10077 = ~n4327 & ~n4632 ;
  assign n10078 = n1702 & ~n10077 ;
  assign n10079 = ~n10076 & ~n10078 ;
  assign n10080 = n307 & n1673 ;
  assign n10081 = n9397 ^ n2156 ;
  assign n10082 = x4 & ~n10081 ;
  assign n10083 = n10082 ^ n2156 ;
  assign n10084 = n1715 & n10083 ;
  assign n10085 = ~n10080 & ~n10084 ;
  assign n10086 = n10079 & n10085 ;
  assign n10087 = ~n10073 & n10086 ;
  assign n10088 = n161 & ~n10087 ;
  assign n10089 = n2743 ^ n2282 ;
  assign n10090 = n10089 ^ n2282 ;
  assign n10091 = n2282 ^ x2 ;
  assign n10092 = n10091 ^ n2282 ;
  assign n10093 = n10090 & ~n10092 ;
  assign n10094 = n10093 ^ n2282 ;
  assign n10095 = x12 & n10094 ;
  assign n10096 = n10095 ^ n2282 ;
  assign n10097 = n692 & n10096 ;
  assign n10098 = n62 & n5949 ;
  assign n10099 = ~n1365 & ~n3264 ;
  assign n10100 = n357 & ~n10099 ;
  assign n10101 = ~n3282 & n10100 ;
  assign n10102 = ~n10098 & ~n10101 ;
  assign n10103 = ~n10097 & n10102 ;
  assign n10104 = n2162 & ~n10103 ;
  assign n10105 = ~n768 & ~n1352 ;
  assign n10106 = n3068 & n3264 ;
  assign n10107 = x8 & n10106 ;
  assign n10108 = n10105 & n10107 ;
  assign n10109 = n214 & n8619 ;
  assign n10110 = n252 & n10109 ;
  assign n10111 = ~n10108 & ~n10110 ;
  assign n10112 = ~x5 & n10111 ;
  assign n10113 = ~n10104 & n10112 ;
  assign n10114 = n1404 & ~n2877 ;
  assign n10115 = x2 ^ x0 ;
  assign n10116 = n10115 ^ x2 ;
  assign n10117 = ~n1438 & ~n2387 ;
  assign n10118 = ~n1298 & n10117 ;
  assign n10119 = n10118 ^ x2 ;
  assign n10120 = ~n10116 & ~n10119 ;
  assign n10121 = n10120 ^ x2 ;
  assign n10122 = n10114 & ~n10121 ;
  assign n10123 = ~n1582 & ~n3824 ;
  assign n10124 = n10123 ^ n10122 ;
  assign n10125 = n4341 ^ n210 ;
  assign n10126 = n10125 ^ n4341 ;
  assign n10127 = n4341 ^ n249 ;
  assign n10128 = n10126 & n10127 ;
  assign n10129 = n10128 ^ n4341 ;
  assign n10130 = n10129 ^ n10122 ;
  assign n10131 = n10124 & ~n10130 ;
  assign n10132 = n10131 ^ n10128 ;
  assign n10133 = n10132 ^ n4341 ;
  assign n10134 = n10133 ^ n10123 ;
  assign n10135 = n10122 & ~n10134 ;
  assign n10136 = n10135 ^ n10122 ;
  assign n10137 = x14 & n10136 ;
  assign n10138 = n10113 & ~n10137 ;
  assign n10139 = ~n10088 & n10138 ;
  assign n10140 = n291 & n4116 ;
  assign n10141 = n2598 & n5973 ;
  assign n10142 = ~n8524 & ~n10141 ;
  assign n10143 = n2709 & ~n10142 ;
  assign n10144 = ~n5960 & ~n10143 ;
  assign n10145 = ~n10140 & n10144 ;
  assign n10146 = ~x9 & ~n10145 ;
  assign n10147 = n1902 & n4869 ;
  assign n10148 = n1073 & n4312 ;
  assign n10149 = ~n7054 & ~n10148 ;
  assign n10150 = ~n9397 & ~n10149 ;
  assign n10151 = ~n10147 & ~n10150 ;
  assign n10152 = n2558 & ~n10151 ;
  assign n10153 = n2168 & n3896 ;
  assign n10154 = n4312 & ~n4737 ;
  assign n10155 = ~n2565 & n2709 ;
  assign n10156 = n10154 & n10155 ;
  assign n10157 = ~n10153 & ~n10156 ;
  assign n10158 = x6 & ~n10157 ;
  assign n10159 = x8 & ~n2169 ;
  assign n10164 = n5174 ^ x2 ;
  assign n10161 = n267 ^ x2 ;
  assign n10160 = n5174 ^ x0 ;
  assign n10162 = n10161 ^ n10160 ;
  assign n10163 = n10162 ^ x2 ;
  assign n10165 = n10164 ^ n10163 ;
  assign n10166 = n10161 ^ n5174 ;
  assign n10167 = n10166 ^ x2 ;
  assign n10168 = n10167 ^ x2 ;
  assign n10169 = n10162 & ~n10168 ;
  assign n10170 = n10169 ^ n10162 ;
  assign n10171 = ~n10167 & n10170 ;
  assign n10172 = n10171 ^ x2 ;
  assign n10173 = ~n10165 & n10172 ;
  assign n10174 = n10173 ^ n10169 ;
  assign n10175 = n10174 ^ x2 ;
  assign n10176 = n10175 ^ x0 ;
  assign n10177 = n10176 ^ n10164 ;
  assign n10178 = n10159 & n10177 ;
  assign n10179 = n609 & ~n1667 ;
  assign n10180 = ~x9 & n394 ;
  assign n10181 = n10179 & n10180 ;
  assign n9971 = n214 & n250 ;
  assign n10182 = n1503 & n9971 ;
  assign n10183 = ~n10181 & ~n10182 ;
  assign n10184 = ~n1716 & ~n10183 ;
  assign n10185 = ~n10178 & ~n10184 ;
  assign n10186 = ~n10158 & n10185 ;
  assign n10187 = ~n10152 & n10186 ;
  assign n10188 = n10187 ^ x12 ;
  assign n10189 = n10188 ^ n10187 ;
  assign n10190 = n394 & n2156 ;
  assign n10191 = ~n284 & n10190 ;
  assign n10192 = ~x13 & n9327 ;
  assign n10193 = ~n10191 & ~n10192 ;
  assign n10194 = ~n1716 & ~n10193 ;
  assign n10195 = n675 & n1670 ;
  assign n10196 = n394 & n2707 ;
  assign n10197 = ~n10195 & ~n10196 ;
  assign n10198 = n1702 & ~n10197 ;
  assign n10199 = ~n10194 & ~n10198 ;
  assign n10200 = n10199 ^ n10187 ;
  assign n10201 = ~n10189 & n10200 ;
  assign n10202 = n10201 ^ n10187 ;
  assign n10203 = ~n10146 & n10202 ;
  assign n10204 = x5 & n10203 ;
  assign n10205 = n10204 ^ n10139 ;
  assign n10206 = ~n10139 & n10205 ;
  assign n10207 = n10206 ^ n10066 ;
  assign n10208 = n10207 ^ n10139 ;
  assign n10209 = n10069 & n10208 ;
  assign n10210 = n10209 ^ n10206 ;
  assign n10211 = n10210 ^ n10139 ;
  assign n10212 = n9999 & ~n10211 ;
  assign n10213 = n10212 ^ n9999 ;
  assign n10214 = x15 & ~n10213 ;
  assign n9866 = ~n1123 & ~n1630 ;
  assign n9867 = ~n1529 & ~n9866 ;
  assign n9868 = n1261 & ~n1528 ;
  assign n9869 = ~n9867 & ~n9868 ;
  assign n9870 = n528 & ~n9869 ;
  assign n9871 = n1231 & n1494 ;
  assign n9872 = ~n9870 & ~n9871 ;
  assign n9873 = n2904 & ~n9872 ;
  assign n9874 = ~n153 & n1404 ;
  assign n9875 = n1261 & n9874 ;
  assign n9876 = ~n9873 & ~n9875 ;
  assign n9877 = n1285 & ~n9876 ;
  assign n9878 = x4 & ~n9559 ;
  assign n9879 = n1542 & n4801 ;
  assign n9880 = ~n9878 & ~n9879 ;
  assign n9881 = n1518 & ~n9880 ;
  assign n9882 = x15 & n9881 ;
  assign n9883 = ~n9877 & ~n9882 ;
  assign n9894 = n18 & n222 ;
  assign n9961 = n604 & n9894 ;
  assign n9962 = n343 & n1261 ;
  assign n9963 = n8969 & n9962 ;
  assign n9964 = ~n9961 & ~n9963 ;
  assign n9884 = ~x8 & n1456 ;
  assign n9885 = n3552 & n9884 ;
  assign n9886 = ~n6477 & ~n9885 ;
  assign n9887 = ~n43 & ~n9886 ;
  assign n9888 = n1390 & n1456 ;
  assign n9889 = ~n9887 & ~n9888 ;
  assign n9890 = x12 & ~n9889 ;
  assign n9891 = n1415 & n1588 ;
  assign n9892 = ~n1623 & ~n9891 ;
  assign n9893 = n1456 & ~n9892 ;
  assign n9895 = x9 & ~n9894 ;
  assign n9896 = ~n9893 & n9895 ;
  assign n9897 = ~n9890 & n9896 ;
  assign n9898 = n9803 ^ x15 ;
  assign n9899 = n9898 ^ x9 ;
  assign n9900 = ~x13 & n1528 ;
  assign n9901 = n9900 ^ x4 ;
  assign n9902 = n9901 ^ n1700 ;
  assign n9904 = n9900 ^ n1078 ;
  assign n9903 = n9902 ^ n9503 ;
  assign n9905 = n9904 ^ n9903 ;
  assign n9906 = n9903 ^ n1078 ;
  assign n9907 = n9906 ^ n9902 ;
  assign n9908 = n9905 & ~n9907 ;
  assign n9909 = n9908 ^ n1078 ;
  assign n9910 = ~n1078 & n1700 ;
  assign n9911 = n9910 ^ n9902 ;
  assign n9912 = ~n9909 & ~n9911 ;
  assign n9913 = n9912 ^ n9910 ;
  assign n9914 = ~n9902 & n9913 ;
  assign n9915 = n9914 ^ n9908 ;
  assign n9916 = n9915 ^ n9900 ;
  assign n9917 = n9916 ^ n1078 ;
  assign n9918 = x5 & ~n9917 ;
  assign n9919 = ~n609 & n3865 ;
  assign n9920 = n18 & n529 ;
  assign n9921 = ~x8 & n1303 ;
  assign n9922 = ~n9920 & ~n9921 ;
  assign n9923 = ~n9919 & n9922 ;
  assign n9924 = n1456 & ~n9923 ;
  assign n9925 = ~n9918 & ~n9924 ;
  assign n9926 = n9925 ^ n2743 ;
  assign n9927 = ~x15 & n9926 ;
  assign n9928 = n9927 ^ n9925 ;
  assign n9929 = ~n9899 & n9928 ;
  assign n9930 = n9929 ^ n9927 ;
  assign n9931 = n9930 ^ n9925 ;
  assign n9932 = n9931 ^ x15 ;
  assign n9933 = ~x9 & ~n9932 ;
  assign n9934 = ~n9897 & ~n9933 ;
  assign n9935 = x8 & ~n701 ;
  assign n9936 = n120 & ~n9935 ;
  assign n9937 = ~n1493 & n9650 ;
  assign n9938 = n1123 & ~n9937 ;
  assign n9939 = ~n9936 & ~n9938 ;
  assign n9940 = n1760 & ~n9939 ;
  assign n9941 = n1511 & n6476 ;
  assign n9942 = ~n9940 & ~n9941 ;
  assign n9943 = ~n9934 & n9942 ;
  assign n9965 = n9964 ^ n9943 ;
  assign n9966 = n9965 ^ n9943 ;
  assign n9944 = n1581 & n2565 ;
  assign n9945 = n1433 & ~n5919 ;
  assign n9946 = ~n9944 & ~n9945 ;
  assign n9947 = n1521 & ~n9946 ;
  assign n9948 = n222 & n3069 ;
  assign n9949 = ~n5355 & ~n9948 ;
  assign n9950 = ~x12 & ~n6110 ;
  assign n9951 = ~n9949 & n9950 ;
  assign n9952 = n1261 & n2886 ;
  assign n9953 = n167 & n6360 ;
  assign n9954 = ~n1490 & n9953 ;
  assign n9955 = ~n9952 & ~n9954 ;
  assign n9956 = ~n9951 & n9955 ;
  assign n9957 = ~n9947 & n9956 ;
  assign n9958 = n1467 & ~n9957 ;
  assign n9959 = n9958 ^ n9943 ;
  assign n9960 = n9959 ^ n9943 ;
  assign n9967 = n9966 ^ n9960 ;
  assign n9968 = x14 & n8969 ;
  assign n9969 = ~n5365 & ~n9968 ;
  assign n9970 = n222 & ~n9969 ;
  assign n9972 = n1518 & n9971 ;
  assign n9973 = ~n9970 & ~n9972 ;
  assign n9974 = n1551 & ~n9973 ;
  assign n9975 = n9974 ^ n9943 ;
  assign n9976 = n9975 ^ n9943 ;
  assign n9977 = n9976 ^ n9966 ;
  assign n9978 = n9966 & ~n9977 ;
  assign n9979 = n9978 ^ n9966 ;
  assign n9980 = ~n9967 & n9979 ;
  assign n9981 = n9980 ^ n9978 ;
  assign n9982 = n9981 ^ n9943 ;
  assign n9983 = n9982 ^ n9966 ;
  assign n9984 = x6 & n9983 ;
  assign n9985 = n9984 ^ n9943 ;
  assign n9986 = n9883 & n9985 ;
  assign n9987 = ~n1716 & ~n9986 ;
  assign n10215 = n10214 ^ n9987 ;
  assign n10216 = n10215 ^ n10214 ;
  assign n10217 = n7159 ^ n2182 ;
  assign n10218 = n10217 ^ n7159 ;
  assign n10219 = n7159 ^ x4 ;
  assign n10220 = n10219 ^ n7159 ;
  assign n10221 = ~n10218 & ~n10220 ;
  assign n10222 = n10221 ^ n7159 ;
  assign n10223 = x8 & n10222 ;
  assign n10224 = n10223 ^ n7159 ;
  assign n10225 = n4506 & n10224 ;
  assign n10226 = x0 & ~n10225 ;
  assign n10227 = ~n1747 & ~n10226 ;
  assign n10228 = ~n3453 & n9327 ;
  assign n10229 = n294 & n403 ;
  assign n10230 = ~n963 & ~n10229 ;
  assign n10231 = ~n133 & ~n1298 ;
  assign n10232 = n7988 & n10231 ;
  assign n10233 = ~n10230 & n10232 ;
  assign n10234 = ~n10228 & ~n10233 ;
  assign n10235 = x8 & ~n10234 ;
  assign n10236 = x15 & ~n5297 ;
  assign n10237 = ~n2105 & n10236 ;
  assign n10238 = ~n291 & ~n10237 ;
  assign n10239 = n9141 & ~n10238 ;
  assign n10240 = n4196 ^ n133 ;
  assign n10241 = x4 & n10240 ;
  assign n10242 = n10241 ^ n133 ;
  assign n10243 = n1404 & n10242 ;
  assign n10244 = n963 & n10243 ;
  assign n10245 = ~n10239 & ~n10244 ;
  assign n10246 = ~n10235 & n10245 ;
  assign n10247 = n1719 & ~n10246 ;
  assign n10248 = n2904 & n4117 ;
  assign n10249 = ~n4530 & ~n10248 ;
  assign n10250 = ~n1404 & ~n4593 ;
  assign n10251 = ~n960 & n10250 ;
  assign n10252 = n10249 & n10251 ;
  assign n10253 = n1285 & ~n10252 ;
  assign n10254 = n1607 & n3018 ;
  assign n10255 = ~n1468 & ~n3217 ;
  assign n10256 = ~n2289 & ~n10255 ;
  assign n10257 = ~n10254 & ~n10256 ;
  assign n10258 = ~n2169 & ~n10257 ;
  assign n10259 = ~n10253 & ~n10258 ;
  assign n10260 = n2904 & n9900 ;
  assign n10261 = ~n214 & ~n10260 ;
  assign n10262 = ~n17 & ~n10261 ;
  assign n10263 = ~n7705 & ~n10262 ;
  assign n10264 = n10263 ^ x6 ;
  assign n10265 = n10264 ^ n10263 ;
  assign n10266 = n10265 ^ n10259 ;
  assign n10267 = n1367 ^ x15 ;
  assign n10276 = n10267 ^ n1367 ;
  assign n10268 = n1367 ^ x8 ;
  assign n10269 = n10268 ^ n10267 ;
  assign n10270 = n10269 ^ n10267 ;
  assign n10271 = n10270 ^ n1367 ;
  assign n10272 = n10269 ^ n4481 ;
  assign n10273 = n10272 ^ n10269 ;
  assign n10274 = n10273 ^ n10271 ;
  assign n10275 = ~n10271 & n10274 ;
  assign n10277 = n10276 ^ n10275 ;
  assign n10278 = n10277 ^ n10271 ;
  assign n10279 = n1367 ^ x13 ;
  assign n10280 = n10275 ^ n10271 ;
  assign n10281 = ~n10279 & ~n10280 ;
  assign n10282 = n10281 ^ n1367 ;
  assign n10283 = ~n10278 & ~n10282 ;
  assign n10284 = n10283 ^ n1367 ;
  assign n10285 = n10284 ^ x15 ;
  assign n10286 = n10285 ^ n1367 ;
  assign n10287 = n10286 ^ x10 ;
  assign n10288 = n10286 & ~n10287 ;
  assign n10289 = n10288 ^ n10263 ;
  assign n10290 = n10289 ^ n10286 ;
  assign n10291 = n10266 & ~n10290 ;
  assign n10292 = n10291 ^ n10288 ;
  assign n10293 = n10292 ^ n10286 ;
  assign n10294 = n10259 & n10293 ;
  assign n10295 = n10294 ^ n10259 ;
  assign n10296 = n228 & ~n10295 ;
  assign n10297 = n1671 & n6448 ;
  assign n10298 = n1953 & n2503 ;
  assign n10299 = ~n10297 & ~n10298 ;
  assign n10300 = x4 & ~n10299 ;
  assign n10301 = n585 & n1256 ;
  assign n10302 = ~n1551 & ~n10301 ;
  assign n10303 = ~x6 & ~n10302 ;
  assign n10304 = ~n9891 & ~n10303 ;
  assign n10305 = n2445 & ~n10304 ;
  assign n10306 = ~n42 & ~n1618 ;
  assign n10307 = n1483 & ~n10306 ;
  assign n10308 = ~n2169 & n10307 ;
  assign n10309 = ~n8733 & n9590 ;
  assign n10310 = ~n10308 & ~n10309 ;
  assign n10311 = x10 & n1669 ;
  assign n10312 = n42 & n153 ;
  assign n10313 = n10311 & n10312 ;
  assign n10314 = ~x9 & n10313 ;
  assign n10315 = n10310 & ~n10314 ;
  assign n10316 = ~n10305 & n10315 ;
  assign n10317 = n247 & ~n10316 ;
  assign n10318 = n2258 & n2724 ;
  assign n10319 = ~n10317 & ~n10318 ;
  assign n10320 = ~n10300 & n10319 ;
  assign n10321 = ~n1528 & n1582 ;
  assign n10322 = x10 & n10321 ;
  assign n10323 = n18 & ~n403 ;
  assign n10324 = ~n8455 & ~n10323 ;
  assign n10325 = ~n4690 & n10324 ;
  assign n10326 = ~n10322 & n10325 ;
  assign n10327 = n4561 & ~n10326 ;
  assign n10330 = n10327 ^ n6471 ;
  assign n10331 = n10330 ^ n10327 ;
  assign n10328 = n10327 ^ n2289 ;
  assign n10329 = n10328 ^ n10327 ;
  assign n10332 = n10331 ^ n10329 ;
  assign n10333 = n10327 ^ x9 ;
  assign n10334 = n10333 ^ n10327 ;
  assign n10335 = n10334 ^ n10331 ;
  assign n10336 = n10331 & n10335 ;
  assign n10337 = n10336 ^ n10331 ;
  assign n10338 = n10332 & n10337 ;
  assign n10339 = n10338 ^ n10336 ;
  assign n10340 = n10339 ^ n10327 ;
  assign n10341 = n10340 ^ n10331 ;
  assign n10342 = ~x2 & n10341 ;
  assign n10343 = n10342 ^ n10327 ;
  assign n10344 = n10320 & ~n10343 ;
  assign n10345 = ~n10296 & n10344 ;
  assign n10346 = n10345 ^ x5 ;
  assign n10347 = n10346 ^ n10345 ;
  assign n10348 = n10347 ^ n10247 ;
  assign n10349 = n475 & n3068 ;
  assign n10350 = n1504 & n10349 ;
  assign n10351 = n254 & n9155 ;
  assign n10352 = ~n2197 & n10351 ;
  assign n10353 = ~n2904 & ~n10352 ;
  assign n10354 = ~n609 & n7569 ;
  assign n10355 = n1484 & n9650 ;
  assign n10356 = ~n10354 & ~n10355 ;
  assign n10357 = ~x9 & n10356 ;
  assign n10358 = ~n10353 & ~n10357 ;
  assign n10359 = x14 & ~n214 ;
  assign n10360 = ~n1902 & n7569 ;
  assign n10361 = ~n10359 & n10360 ;
  assign n10362 = ~n10358 & ~n10361 ;
  assign n10363 = ~x10 & ~n10362 ;
  assign n10364 = ~n10350 & ~n10363 ;
  assign n10365 = n10364 ^ x2 ;
  assign n10366 = x2 & ~n10365 ;
  assign n10367 = n10366 ^ n10345 ;
  assign n10368 = n10367 ^ x2 ;
  assign n10369 = n10348 & ~n10368 ;
  assign n10370 = n10369 ^ n10366 ;
  assign n10371 = n10370 ^ x2 ;
  assign n10372 = ~n10247 & n10371 ;
  assign n10373 = n10372 ^ n10247 ;
  assign n10374 = ~n10227 & ~n10373 ;
  assign n10375 = n1368 ^ n291 ;
  assign n10376 = n10375 ^ n1506 ;
  assign n10377 = n10376 ^ n1368 ;
  assign n10378 = n10377 ^ n10376 ;
  assign n10379 = x14 ^ x9 ;
  assign n10380 = n9755 & ~n10379 ;
  assign n10381 = n10380 ^ x9 ;
  assign n10382 = n38 & n10381 ;
  assign n10383 = n10382 ^ n10376 ;
  assign n10384 = n10383 ^ n10375 ;
  assign n10385 = n10378 & ~n10384 ;
  assign n10386 = n10385 ^ n10382 ;
  assign n10387 = ~n2309 & ~n10382 ;
  assign n10388 = n10387 ^ n10375 ;
  assign n10389 = ~n10386 & ~n10388 ;
  assign n10390 = n10389 ^ n10387 ;
  assign n10391 = ~n10375 & n10390 ;
  assign n10392 = n10391 ^ n10385 ;
  assign n10393 = n10392 ^ n291 ;
  assign n10394 = n10393 ^ n10382 ;
  assign n10395 = n190 & ~n10394 ;
  assign n10396 = n2422 & n9093 ;
  assign n10397 = n1231 & n10396 ;
  assign n10398 = n33 & n1214 ;
  assign n10399 = ~n9115 & ~n10398 ;
  assign n10400 = n2445 & ~n10399 ;
  assign n10401 = n1518 & n8983 ;
  assign n10402 = n1252 & n8047 ;
  assign n10403 = ~n10401 & ~n10402 ;
  assign n10404 = ~n1511 & n10403 ;
  assign n10405 = ~n10400 & n10404 ;
  assign n10406 = n394 & ~n10405 ;
  assign n10407 = ~n10397 & ~n10406 ;
  assign n10408 = ~n10395 & n10407 ;
  assign n10409 = n1718 & ~n10408 ;
  assign n10410 = n38 & n2445 ;
  assign n10411 = n71 & n269 ;
  assign n10412 = n10410 & n10411 ;
  assign n10413 = n1303 & n1420 ;
  assign n10414 = n2506 & n10413 ;
  assign n10415 = ~n1368 & ~n2886 ;
  assign n10416 = n394 & ~n10415 ;
  assign n10417 = n1902 & n6583 ;
  assign n10418 = ~n10416 & ~n10417 ;
  assign n10419 = n9550 & ~n10418 ;
  assign n10420 = ~n10414 & ~n10419 ;
  assign n10421 = ~n10412 & n10420 ;
  assign n10422 = n1834 & ~n10421 ;
  assign n10423 = ~n10409 & ~n10422 ;
  assign n10424 = x12 & ~n2708 ;
  assign n10425 = ~n470 & n10424 ;
  assign n10426 = ~n9874 & ~n10425 ;
  assign n10427 = n394 & ~n10426 ;
  assign n10428 = n570 & n2761 ;
  assign n10429 = n8970 ^ n2904 ;
  assign n10430 = n10429 ^ n2506 ;
  assign n10431 = n5065 ^ n1608 ;
  assign n10432 = n8970 & ~n10431 ;
  assign n10433 = n10432 ^ n5065 ;
  assign n10434 = n10430 & ~n10433 ;
  assign n10435 = n10434 ^ n10432 ;
  assign n10436 = n10435 ^ n5065 ;
  assign n10437 = n10436 ^ n8970 ;
  assign n10438 = ~n2506 & ~n10437 ;
  assign n10439 = n10438 ^ x12 ;
  assign n10440 = n10439 ^ n10438 ;
  assign n10441 = n1550 & n2565 ;
  assign n10442 = ~n6449 & ~n10441 ;
  assign n10443 = n1618 & ~n10442 ;
  assign n10444 = ~n5397 & ~n10443 ;
  assign n10445 = n10444 ^ n10438 ;
  assign n10446 = ~n10440 & n10445 ;
  assign n10447 = n10446 ^ n10438 ;
  assign n10448 = ~x4 & ~n10447 ;
  assign n10449 = ~n10428 & ~n10448 ;
  assign n10450 = ~n10427 & n10449 ;
  assign n10451 = n1953 & ~n10450 ;
  assign n10452 = n4713 & n9834 ;
  assign n10453 = n5408 & n5994 ;
  assign n10454 = ~n10452 & ~n10453 ;
  assign n10455 = ~x2 & ~n10454 ;
  assign n10456 = n1511 & n4561 ;
  assign n10457 = n1506 & n9580 ;
  assign n10458 = ~n10456 & ~n10457 ;
  assign n10459 = n3728 & ~n10458 ;
  assign n10460 = ~n10455 & ~n10459 ;
  assign n10461 = n249 & n1395 ;
  assign n10462 = ~n3227 & ~n10461 ;
  assign n10463 = ~n2761 & n10462 ;
  assign n10464 = n1758 & ~n10463 ;
  assign n10465 = n6966 & ~n8970 ;
  assign n10466 = n570 & n1608 ;
  assign n10467 = ~n10465 & ~n10466 ;
  assign n10468 = n20 & n1467 ;
  assign n10469 = ~n10467 & n10468 ;
  assign n10470 = ~n10464 & ~n10469 ;
  assign n10471 = n10460 & n10470 ;
  assign n10472 = ~x2 & ~n1252 ;
  assign n10473 = ~n2444 & ~n10472 ;
  assign n10474 = n2005 & ~n2233 ;
  assign n10475 = n7507 & n10474 ;
  assign n10476 = ~x15 & ~n2558 ;
  assign n10477 = n153 & n2548 ;
  assign n10478 = ~n10476 & n10477 ;
  assign n10479 = ~n10475 & ~n10478 ;
  assign n10480 = ~n10473 & n10479 ;
  assign n10481 = n1797 & ~n10480 ;
  assign n10482 = n3508 & ~n8970 ;
  assign n10483 = ~n2752 & ~n10482 ;
  assign n10484 = n33 & ~n10483 ;
  assign n10485 = ~n470 & n1608 ;
  assign n10486 = ~n6737 & ~n8973 ;
  assign n10487 = ~n10485 & n10486 ;
  assign n10488 = n266 & ~n10487 ;
  assign n10489 = ~n9834 & ~n10488 ;
  assign n10490 = ~n10484 & n10489 ;
  assign n10491 = n2410 & ~n10490 ;
  assign n10492 = ~n10481 & ~n10491 ;
  assign n10493 = n10471 & n10492 ;
  assign n10494 = ~n10451 & n10493 ;
  assign n10495 = x5 & ~n10494 ;
  assign n10496 = n214 & n2192 ;
  assign n10497 = n2282 & n10496 ;
  assign n10498 = ~x0 & ~n10497 ;
  assign n10499 = ~n10495 & n10498 ;
  assign n10500 = n10423 & n10499 ;
  assign n10501 = ~n10374 & ~n10500 ;
  assign n10502 = n10501 ^ n10214 ;
  assign n10503 = n10502 ^ n10214 ;
  assign n10504 = ~n10216 & ~n10503 ;
  assign n10505 = n10504 ^ n10214 ;
  assign n10506 = x7 & ~n10505 ;
  assign n10507 = n10506 ^ n10214 ;
  assign n10508 = n9865 & ~n10507 ;
  assign n10509 = n9831 & n10508 ;
  assign n10510 = ~n9793 & ~n10509 ;
  assign n10511 = x8 & n9180 ;
  assign n10512 = ~n2124 & ~n10511 ;
  assign n10513 = n1597 & ~n10512 ;
  assign n10514 = n1630 & n9555 ;
  assign n10515 = n1607 & n10514 ;
  assign n10516 = ~n10513 & ~n10515 ;
  assign n10517 = n3821 & ~n10516 ;
  assign n10518 = ~x1 & n10517 ;
  assign n10519 = n5647 & n7884 ;
  assign n10520 = n33 & n1457 ;
  assign n10521 = x2 & n450 ;
  assign n10522 = n10520 & n10521 ;
  assign n10523 = n10519 & n10522 ;
  assign n10524 = ~n450 & ~n1716 ;
  assign n10525 = ~n2042 & n10524 ;
  assign n10526 = ~x8 & n9093 ;
  assign n10527 = ~n200 & n10526 ;
  assign n10528 = n10525 & n10527 ;
  assign n10529 = n310 & n6708 ;
  assign n10530 = n2659 & n10529 ;
  assign n10531 = ~n10528 & ~n10530 ;
  assign n10532 = n1265 & ~n10531 ;
  assign n10533 = ~n10523 & ~n10532 ;
  assign n10534 = ~n10518 & n10533 ;
  assign n10535 = n2452 & ~n10534 ;
  assign n10536 = n1267 & n1404 ;
  assign n10537 = ~n6646 & ~n10536 ;
  assign n10538 = n24 & n1454 ;
  assign n10539 = ~n3507 & ~n5633 ;
  assign n10540 = ~n10538 & n10539 ;
  assign n10541 = n434 & ~n10540 ;
  assign n10542 = ~n319 & ~n880 ;
  assign n10543 = n10542 ^ n792 ;
  assign n10544 = n10543 ^ n792 ;
  assign n10545 = n1073 ^ n792 ;
  assign n10546 = n10545 ^ n792 ;
  assign n10547 = ~n10544 & n10546 ;
  assign n10548 = n10547 ^ n792 ;
  assign n10549 = ~x5 & n10548 ;
  assign n10550 = n10549 ^ n792 ;
  assign n10551 = ~n10541 & ~n10550 ;
  assign n10552 = x10 & ~n10551 ;
  assign n10553 = n450 & n1261 ;
  assign n10554 = ~n1106 & ~n10553 ;
  assign n10555 = ~x12 & ~n3552 ;
  assign n10556 = ~n10554 & n10555 ;
  assign n10557 = n3839 & n4746 ;
  assign n10558 = n1138 & n10557 ;
  assign n10559 = ~n10556 & ~n10558 ;
  assign n10560 = ~n470 & ~n10559 ;
  assign n10561 = n107 & n1303 ;
  assign n10562 = n475 & ~n1700 ;
  assign n10563 = n132 & n10562 ;
  assign n10564 = ~n10561 & ~n10563 ;
  assign n10565 = n1438 & ~n10564 ;
  assign n10566 = n10565 ^ x1 ;
  assign n10567 = n10566 ^ n10565 ;
  assign n10568 = n10567 ^ n10560 ;
  assign n10569 = x13 ^ x10 ;
  assign n10570 = x13 ^ x5 ;
  assign n10571 = n10570 ^ x5 ;
  assign n10572 = n1261 ^ x5 ;
  assign n10573 = n10571 & n10572 ;
  assign n10574 = n10573 ^ x5 ;
  assign n10575 = ~n10569 & n10574 ;
  assign n10576 = n3652 & n10575 ;
  assign n10577 = n222 & n3545 ;
  assign n10578 = ~n10576 & ~n10577 ;
  assign n10579 = n10578 ^ x12 ;
  assign n10580 = ~x12 & n10579 ;
  assign n10581 = n10580 ^ n10565 ;
  assign n10582 = n10581 ^ x12 ;
  assign n10583 = n10568 & ~n10582 ;
  assign n10584 = n10583 ^ n10580 ;
  assign n10585 = n10584 ^ x12 ;
  assign n10586 = ~n10560 & ~n10585 ;
  assign n10587 = n10586 ^ n10560 ;
  assign n10588 = ~n10552 & ~n10587 ;
  assign n10589 = x2 & ~n10588 ;
  assign n10590 = n5669 & n8471 ;
  assign n10591 = ~x1 & n1123 ;
  assign n10592 = n816 & ~n1467 ;
  assign n10593 = ~n10591 & ~n10592 ;
  assign n10594 = ~n450 & ~n2331 ;
  assign n10595 = ~n1438 & ~n1456 ;
  assign n10596 = n10594 & n10595 ;
  assign n10597 = ~x1 & ~n470 ;
  assign n10598 = ~n153 & n1597 ;
  assign n10599 = ~n10597 & ~n10598 ;
  assign n10600 = ~x2 & ~n1552 ;
  assign n10601 = ~n1457 & n10600 ;
  assign n10602 = ~n10599 & n10601 ;
  assign n10603 = n10596 & n10602 ;
  assign n10604 = n10593 & n10603 ;
  assign n10605 = ~n10590 & ~n10604 ;
  assign n10606 = ~n10589 & n10605 ;
  assign n10607 = ~n10537 & ~n10606 ;
  assign n10608 = n3232 & n4951 ;
  assign n10609 = ~x2 & n2555 ;
  assign n10610 = n3865 & n10609 ;
  assign n10611 = n1969 & n3048 ;
  assign n10612 = ~n1672 & n10611 ;
  assign n10613 = ~n10610 & ~n10612 ;
  assign n10614 = n222 & ~n10613 ;
  assign n10615 = n280 & ~n1285 ;
  assign n10616 = n244 & n10615 ;
  assign n10617 = n3290 & n10616 ;
  assign n10618 = ~n10614 & ~n10617 ;
  assign n10619 = ~n10608 & n10618 ;
  assign n10620 = n264 & ~n10619 ;
  assign n10621 = n429 & n2506 ;
  assign n10622 = n7644 & n10621 ;
  assign n10623 = n1622 & n3226 ;
  assign n10624 = ~n25 & n2105 ;
  assign n10625 = n2397 & n10624 ;
  assign n10626 = n10623 & n10625 ;
  assign n10627 = n132 & n3532 ;
  assign n10628 = n2491 & n10627 ;
  assign n10629 = ~n10626 & ~n10628 ;
  assign n10630 = ~n10622 & n10629 ;
  assign n10631 = ~n10620 & n10630 ;
  assign n10632 = x13 & ~n10631 ;
  assign n10633 = n2186 & n3058 ;
  assign n10634 = n71 & n10633 ;
  assign n10635 = n2304 & n4561 ;
  assign n10636 = n3678 & n10635 ;
  assign n10637 = ~n10634 & ~n10636 ;
  assign n10638 = ~x1 & n4304 ;
  assign n10639 = ~n10637 & n10638 ;
  assign n10640 = n2369 & n10521 ;
  assign n10641 = n7916 & n10640 ;
  assign n10642 = n2075 & n3294 ;
  assign n10643 = ~n470 & n10642 ;
  assign n10644 = n7650 & n10643 ;
  assign n10645 = ~n10641 & ~n10644 ;
  assign n10646 = ~n2169 & ~n10645 ;
  assign n10647 = n1404 & n6787 ;
  assign n10648 = n1779 & n10647 ;
  assign n10649 = ~n10646 & ~n10648 ;
  assign n10650 = ~n10639 & n10649 ;
  assign n10651 = ~n2218 & ~n10650 ;
  assign n10662 = n2929 & n6499 ;
  assign n10663 = n229 & n8764 ;
  assign n10664 = ~n10662 & ~n10663 ;
  assign n10652 = n1285 & n4850 ;
  assign n10653 = x4 ^ x2 ;
  assign n10654 = n1969 ^ n1747 ;
  assign n10655 = n1747 ^ x4 ;
  assign n10656 = n10655 ^ n1747 ;
  assign n10657 = n10654 & n10656 ;
  assign n10658 = n10657 ^ n1747 ;
  assign n10659 = ~n10653 & n10658 ;
  assign n10660 = n1672 & n10659 ;
  assign n10661 = ~n10652 & ~n10660 ;
  assign n10665 = n10664 ^ n10661 ;
  assign n10666 = n10664 ^ x9 ;
  assign n10667 = n10666 ^ n10664 ;
  assign n10668 = n10667 ^ n25 ;
  assign n10669 = n10668 ^ x7 ;
  assign n10670 = n10665 & n10669 ;
  assign n10671 = n10670 ^ n10664 ;
  assign n10672 = n25 & n10671 ;
  assign n10673 = n10672 ^ n25 ;
  assign n10674 = ~n10651 & ~n10673 ;
  assign n10675 = ~n10632 & n10674 ;
  assign n10676 = ~n10607 & n10675 ;
  assign n10677 = ~n10535 & n10676 ;
  assign n10678 = ~n10510 & n10677 ;
  assign n10679 = ~n8968 & n10678 ;
  assign n10680 = n10679 ^ x3 ;
  assign n10681 = n10680 ^ n10679 ;
  assign n10682 = n7630 & n10553 ;
  assign n10683 = n1332 & ~n5650 ;
  assign n10684 = n1123 & ~n1747 ;
  assign n10685 = ~n10683 & ~n10684 ;
  assign n10688 = n10685 ^ x5 ;
  assign n10689 = n10688 ^ n10685 ;
  assign n10686 = n10685 ^ n1073 ;
  assign n10687 = n10686 ^ n10685 ;
  assign n10690 = n10689 ^ n10687 ;
  assign n10691 = x4 & n1970 ;
  assign n10692 = n10691 ^ n10685 ;
  assign n10693 = n10692 ^ n10685 ;
  assign n10694 = n10693 ^ n10689 ;
  assign n10695 = ~n10689 & n10694 ;
  assign n10696 = n10695 ^ n10689 ;
  assign n10697 = n10690 & ~n10696 ;
  assign n10698 = n10697 ^ n10695 ;
  assign n10699 = n10698 ^ n10685 ;
  assign n10700 = n10699 ^ n10689 ;
  assign n10701 = x1 & n10700 ;
  assign n10702 = n10701 ^ n10685 ;
  assign n10703 = n8186 & ~n10702 ;
  assign n10704 = ~n10682 & ~n10703 ;
  assign n10705 = n2005 & ~n10704 ;
  assign n10706 = n1073 & ~n4747 ;
  assign n10707 = ~n799 & n1969 ;
  assign n10708 = ~n10706 & ~n10707 ;
  assign n10709 = n7492 & ~n10708 ;
  assign n10710 = n793 & n6824 ;
  assign n10711 = ~n10709 & ~n10710 ;
  assign n10712 = x2 & n431 ;
  assign n10713 = ~n10711 & n10712 ;
  assign n10714 = ~x5 & n2931 ;
  assign n10715 = n10642 & n10714 ;
  assign n10716 = ~n10713 & ~n10715 ;
  assign n10717 = ~n10705 & n10716 ;
  assign n10718 = x13 & ~n10717 ;
  assign n10719 = ~n5353 & ~n9488 ;
  assign n10720 = ~n43 & ~n10719 ;
  assign n10721 = n2565 & n9019 ;
  assign n10722 = ~n10720 & ~n10721 ;
  assign n10723 = x12 & ~n10722 ;
  assign n10724 = ~n1526 & ~n10723 ;
  assign n10725 = n3728 & ~n10724 ;
  assign n10726 = ~n5299 & ~n10725 ;
  assign n10727 = n17 & ~n10726 ;
  assign n10728 = n2005 & ~n9045 ;
  assign n10729 = x5 & ~n10728 ;
  assign n10730 = ~x9 & ~n2439 ;
  assign n10731 = n10730 ^ x6 ;
  assign n10732 = n10731 ^ n2126 ;
  assign n10733 = n4713 ^ x5 ;
  assign n10734 = x6 & ~n10733 ;
  assign n10735 = n10734 ^ x5 ;
  assign n10736 = n10732 & ~n10735 ;
  assign n10737 = n10736 ^ n10734 ;
  assign n10738 = n10737 ^ x5 ;
  assign n10739 = n10738 ^ x6 ;
  assign n10740 = ~n2126 & ~n10739 ;
  assign n10741 = ~n10729 & n10740 ;
  assign n10742 = ~n2182 & n2225 ;
  assign n10743 = ~n2247 & ~n10742 ;
  assign n10744 = ~n1801 & ~n10743 ;
  assign n10745 = ~n10741 & n10744 ;
  assign n10746 = ~n1266 & n1588 ;
  assign n10747 = n6817 ^ x10 ;
  assign n10748 = ~x13 & ~n1706 ;
  assign n10749 = n10748 ^ x10 ;
  assign n10750 = ~n10747 & n10749 ;
  assign n10751 = n10750 ^ x10 ;
  assign n10752 = ~n10746 & n10751 ;
  assign n10753 = n2483 & ~n10752 ;
  assign n10754 = ~x13 & n1469 ;
  assign n10755 = n5299 & ~n10754 ;
  assign n10756 = ~x6 & n9067 ;
  assign n10757 = ~n10755 & ~n10756 ;
  assign n10758 = ~n10753 & n10757 ;
  assign n10759 = n2397 & ~n10758 ;
  assign n10760 = n2410 & n5344 ;
  assign n10761 = x9 & n10760 ;
  assign n10762 = ~n10759 & ~n10761 ;
  assign n10763 = ~n10745 & n10762 ;
  assign n10764 = ~n10727 & n10763 ;
  assign n10765 = x4 & ~n10764 ;
  assign n10766 = ~x8 & n9891 ;
  assign n10767 = x6 & ~n2225 ;
  assign n10768 = ~n10766 & n10767 ;
  assign n10769 = ~n1646 & n10768 ;
  assign n10770 = n1562 & n2483 ;
  assign n10771 = n1123 & ~n7711 ;
  assign n10772 = ~n10770 & n10771 ;
  assign n10773 = ~n10769 & n10772 ;
  assign n10774 = ~n153 & n2105 ;
  assign n10775 = ~n9580 & ~n10774 ;
  assign n10776 = n17 & ~n10775 ;
  assign n10777 = ~n8987 & ~n10776 ;
  assign n10778 = n1261 & ~n10777 ;
  assign n10779 = ~n10773 & ~n10778 ;
  assign n10780 = ~n9575 & n10779 ;
  assign n10781 = ~x2 & ~n10780 ;
  assign n10782 = ~n10765 & ~n10781 ;
  assign n10783 = n816 & ~n10782 ;
  assign n10784 = n1550 & n3048 ;
  assign n10785 = n1261 & n1440 ;
  assign n10786 = n10784 & n10785 ;
  assign n10787 = ~n3377 & ~n3926 ;
  assign n10788 = n295 & ~n10787 ;
  assign n10789 = n1435 & n4883 ;
  assign n10790 = ~n2920 & n2921 ;
  assign n10791 = n280 & n10790 ;
  assign n10792 = ~n10789 & ~n10791 ;
  assign n10793 = ~n10788 & n10792 ;
  assign n10794 = x8 & ~n10793 ;
  assign n10795 = n1286 & n3048 ;
  assign n10796 = n1265 & n3728 ;
  assign n10797 = ~n10795 & ~n10796 ;
  assign n10798 = n5647 & ~n10797 ;
  assign n10799 = ~n10794 & ~n10798 ;
  assign n10801 = ~n249 & ~n3926 ;
  assign n10800 = n1352 ^ x10 ;
  assign n10802 = n10801 ^ n10800 ;
  assign n10803 = n10801 ^ x2 ;
  assign n10804 = n10803 ^ n10801 ;
  assign n10805 = ~n10802 & n10804 ;
  assign n10806 = n10805 ^ n10801 ;
  assign n10807 = n5344 & ~n10806 ;
  assign n10808 = n10799 & ~n10807 ;
  assign n10809 = ~x9 & ~n10808 ;
  assign n10810 = ~n10786 & ~n10809 ;
  assign n10811 = x5 & ~n2602 ;
  assign n10812 = n291 & n7278 ;
  assign n10813 = ~n10811 & ~n10812 ;
  assign n10814 = n1760 & ~n10813 ;
  assign n10815 = ~n253 & n1953 ;
  assign n10816 = n5299 & n10815 ;
  assign n10817 = ~n10814 & ~n10816 ;
  assign n10818 = n343 & ~n10817 ;
  assign n10819 = n1953 & ~n4944 ;
  assign n10820 = x12 ^ x5 ;
  assign n10821 = n4737 ^ x12 ;
  assign n10822 = n10821 ^ n4737 ;
  assign n10823 = n7988 ^ n4737 ;
  assign n10824 = n10822 & n10823 ;
  assign n10825 = n10824 ^ n4737 ;
  assign n10826 = ~n10820 & n10825 ;
  assign n10827 = n10819 & n10826 ;
  assign n10828 = x15 & n295 ;
  assign n10829 = ~n963 & ~n3314 ;
  assign n10830 = x6 & ~n10829 ;
  assign n10831 = ~n10828 & ~n10830 ;
  assign n10832 = n1420 & n1991 ;
  assign n10833 = ~n10831 & n10832 ;
  assign n10834 = ~n10827 & ~n10833 ;
  assign n10835 = ~n10818 & n10834 ;
  assign n10836 = n1608 & ~n10835 ;
  assign n10837 = x8 ^ x2 ;
  assign n10838 = n10837 ^ x10 ;
  assign n10839 = x8 ^ x5 ;
  assign n10840 = n10839 ^ n10838 ;
  assign n10841 = n8471 ^ x10 ;
  assign n10842 = x5 & ~n10841 ;
  assign n10843 = n10842 ^ n8471 ;
  assign n10844 = n10840 & n10843 ;
  assign n10845 = n10844 ^ n10842 ;
  assign n10846 = n10845 ^ n8471 ;
  assign n10847 = n10846 ^ x5 ;
  assign n10848 = ~n10838 & n10847 ;
  assign n10849 = n252 & n10848 ;
  assign n10850 = n1261 & n8253 ;
  assign n10851 = ~n10849 & ~n10850 ;
  assign n10852 = ~n1290 & ~n1630 ;
  assign n10853 = ~n19 & ~n10852 ;
  assign n10854 = n4047 & n10853 ;
  assign n10855 = n10854 ^ x4 ;
  assign n10856 = n10855 ^ n10854 ;
  assign n10857 = n10856 ^ n10851 ;
  assign n10858 = ~n1623 & ~n2124 ;
  assign n10859 = ~n8455 & n10858 ;
  assign n10860 = n1801 & ~n10859 ;
  assign n10861 = ~n18 & ~n38 ;
  assign n10862 = n1834 & ~n10861 ;
  assign n10863 = ~n295 & ~n10862 ;
  assign n10864 = ~n19 & ~n10863 ;
  assign n10865 = ~n10860 & ~n10864 ;
  assign n10866 = n10865 ^ x6 ;
  assign n10867 = ~x6 & n10866 ;
  assign n10868 = n10867 ^ n10854 ;
  assign n10869 = n10868 ^ x6 ;
  assign n10870 = n10857 & ~n10869 ;
  assign n10871 = n10870 ^ n10867 ;
  assign n10872 = n10871 ^ x6 ;
  assign n10873 = n10851 & ~n10872 ;
  assign n10874 = n10873 ^ n10851 ;
  assign n10875 = x9 & ~n10874 ;
  assign n10876 = ~n3010 & n9471 ;
  assign n10877 = n1562 & n10876 ;
  assign n10878 = ~n10875 & ~n10877 ;
  assign n10879 = ~n10836 & n10878 ;
  assign n10880 = n1397 & n1760 ;
  assign n10881 = ~n291 & ~n6476 ;
  assign n10882 = n2181 ^ x9 ;
  assign n10883 = x10 ^ x9 ;
  assign n10884 = n10883 ^ x5 ;
  assign n10885 = n10884 ^ x9 ;
  assign n10886 = n10882 & ~n10885 ;
  assign n10887 = n10886 ^ x9 ;
  assign n10888 = n10881 ^ n2342 ;
  assign n10889 = n10887 & ~n10888 ;
  assign n10890 = n10889 ^ n2342 ;
  assign n10891 = ~n10881 & n10890 ;
  assign n10892 = n10891 ^ n10881 ;
  assign n10893 = ~n10880 & n10892 ;
  assign n10894 = x2 & ~n10893 ;
  assign n10895 = ~x9 & n280 ;
  assign n10896 = n2991 & n10895 ;
  assign n10897 = ~n10894 & ~n10896 ;
  assign n10898 = ~n470 & ~n10897 ;
  assign n10900 = n291 & ~n1700 ;
  assign n10901 = ~n1772 & ~n10900 ;
  assign n10899 = ~x4 & ~n1706 ;
  assign n10902 = n10901 ^ n10899 ;
  assign n10903 = n10902 ^ n10901 ;
  assign n10904 = n10901 ^ n1352 ;
  assign n10905 = n10904 ^ n10901 ;
  assign n10906 = ~n10903 & ~n10905 ;
  assign n10907 = n10906 ^ n10901 ;
  assign n10908 = x2 & ~n10907 ;
  assign n10909 = n10908 ^ n10901 ;
  assign n10910 = n9112 & ~n10909 ;
  assign n10911 = ~n10898 & ~n10910 ;
  assign n10912 = n9900 & ~n10911 ;
  assign n10913 = n207 & ~n504 ;
  assign n10914 = ~n247 & ~n2598 ;
  assign n10915 = ~n1322 & ~n10914 ;
  assign n10916 = ~n4341 & ~n10915 ;
  assign n10917 = ~n10913 & n10916 ;
  assign n10918 = x10 & ~n10917 ;
  assign n10919 = n3627 & n4883 ;
  assign n10920 = ~n10918 & ~n10919 ;
  assign n10921 = n5647 & ~n10920 ;
  assign n10922 = ~n247 & ~n6476 ;
  assign n10923 = ~n1285 & ~n1492 ;
  assign n10924 = ~n10922 & ~n10923 ;
  assign n10925 = ~n249 & n10615 ;
  assign n10926 = ~n10924 & ~n10925 ;
  assign n10927 = n1394 & ~n10926 ;
  assign n10928 = n2397 & n8111 ;
  assign n10929 = ~n10927 & ~n10928 ;
  assign n10930 = n3865 & n10811 ;
  assign n10931 = n1286 & n1834 ;
  assign n10932 = x12 & n10931 ;
  assign n10933 = ~n10930 & ~n10932 ;
  assign n10934 = n10929 & n10933 ;
  assign n10935 = ~n10921 & n10934 ;
  assign n10936 = n1366 & ~n10935 ;
  assign n10937 = ~n10912 & ~n10936 ;
  assign n10938 = n10879 & n10937 ;
  assign n10939 = n10810 & n10938 ;
  assign n10940 = n24 & ~n10939 ;
  assign n10941 = ~n10783 & ~n10940 ;
  assign n10942 = x10 & n2282 ;
  assign n10943 = ~x10 & n2397 ;
  assign n10944 = ~n10942 & ~n10943 ;
  assign n10945 = n5432 & ~n10944 ;
  assign n10946 = ~n1716 & n10945 ;
  assign n10947 = ~n3226 & ~n3232 ;
  assign n10948 = ~n2694 & ~n2872 ;
  assign n10949 = ~n10947 & n10948 ;
  assign n10950 = n1138 & n10949 ;
  assign n10951 = ~n18 & ~n1559 ;
  assign n10952 = ~n1716 & ~n10951 ;
  assign n10953 = n1493 & n1952 ;
  assign n10954 = ~n58 & n10953 ;
  assign n10955 = ~n10952 & ~n10954 ;
  assign n10956 = n5156 & ~n10955 ;
  assign n10957 = ~n1352 & ~n1702 ;
  assign n10958 = ~n210 & ~n3848 ;
  assign n10959 = ~n19 & n10958 ;
  assign n10960 = ~n10957 & n10959 ;
  assign n10961 = n17 & n3009 ;
  assign n10962 = ~n5184 & n8195 ;
  assign n10963 = ~n10961 & ~n10962 ;
  assign n10964 = ~n10960 & n10963 ;
  assign n10965 = n10964 ^ x5 ;
  assign n10966 = n10965 ^ n10964 ;
  assign n10967 = ~n1435 & n8823 ;
  assign n10968 = n9048 & n10967 ;
  assign n10969 = x0 & n10600 ;
  assign n10970 = ~n153 & n10969 ;
  assign n10971 = ~n10968 & ~n10970 ;
  assign n10972 = n4052 & ~n10971 ;
  assign n10973 = n1303 & n8619 ;
  assign n10974 = ~n1719 & ~n1955 ;
  assign n10975 = n1581 & ~n10974 ;
  assign n10976 = ~n10973 & ~n10975 ;
  assign n10977 = ~n10972 & n10976 ;
  assign n10978 = x6 & ~n10977 ;
  assign n10979 = n1551 & n2282 ;
  assign n10980 = ~n2397 & ~n10979 ;
  assign n10981 = n2687 & ~n10980 ;
  assign n10982 = ~n133 & ~n1260 ;
  assign n10983 = n10982 ^ x6 ;
  assign n10984 = n10983 ^ n10982 ;
  assign n10985 = n10982 ^ n9160 ;
  assign n10986 = n10985 ^ n10982 ;
  assign n10987 = ~n10984 & n10986 ;
  assign n10988 = n10987 ^ n10982 ;
  assign n10989 = x2 & n10988 ;
  assign n10990 = n10989 ^ n10982 ;
  assign n10991 = n1506 & n10990 ;
  assign n10992 = ~n2387 & ~n4505 ;
  assign n10993 = ~x2 & x15 ;
  assign n10994 = n153 & ~n10993 ;
  assign n10995 = n10992 & ~n10994 ;
  assign n10996 = n1504 & n10995 ;
  assign n10997 = ~n10991 & ~n10996 ;
  assign n10998 = ~n1970 & ~n10997 ;
  assign n10999 = ~n10981 & ~n10998 ;
  assign n11000 = ~n10978 & n10999 ;
  assign n11001 = n11000 ^ n10964 ;
  assign n11002 = ~n10966 & n11001 ;
  assign n11003 = n11002 ^ n10964 ;
  assign n11004 = ~n10956 & n11003 ;
  assign n11005 = x1 & ~n11004 ;
  assign n11006 = ~n10950 & ~n11005 ;
  assign n11007 = ~n10946 & n11006 ;
  assign n11008 = ~x9 & ~n11007 ;
  assign n11009 = n1290 & n7853 ;
  assign n11010 = ~n1597 & ~n9111 ;
  assign n11011 = x4 & ~n11010 ;
  assign n11012 = ~n1285 & n11011 ;
  assign n11013 = ~n11009 & ~n11012 ;
  assign n11016 = n11013 ^ n2218 ;
  assign n11017 = n11016 ^ n11013 ;
  assign n11014 = n11013 ^ x10 ;
  assign n11015 = n11014 ^ n11013 ;
  assign n11018 = n11017 ^ n11015 ;
  assign n11019 = n11013 ^ x4 ;
  assign n11020 = n11019 ^ n11013 ;
  assign n11021 = n11020 ^ n11017 ;
  assign n11022 = ~n11017 & n11021 ;
  assign n11023 = n11022 ^ n11017 ;
  assign n11024 = ~n11018 & ~n11023 ;
  assign n11025 = n11024 ^ n11022 ;
  assign n11026 = n11025 ^ n11013 ;
  assign n11027 = n11026 ^ n11017 ;
  assign n11028 = x8 & n11027 ;
  assign n11029 = n11028 ^ n11013 ;
  assign n11030 = n286 & ~n11029 ;
  assign n11031 = n1597 & n2548 ;
  assign n11032 = ~n1674 & n11031 ;
  assign n11033 = n1285 & n5949 ;
  assign n11034 = n222 & n11033 ;
  assign n11035 = x9 & n295 ;
  assign n11036 = n133 & n9112 ;
  assign n11037 = ~n11035 & ~n11036 ;
  assign n11038 = n1670 & n1733 ;
  assign n11039 = ~n11037 & n11038 ;
  assign n11040 = ~n11034 & ~n11039 ;
  assign n11041 = ~n11032 & n11040 ;
  assign n11042 = ~n11030 & n11041 ;
  assign n11043 = ~x1 & ~n11042 ;
  assign n11044 = x1 & ~n1073 ;
  assign n11045 = x10 & ~n1352 ;
  assign n11046 = n11044 & n11045 ;
  assign n11047 = n2405 & n11046 ;
  assign n11048 = n3172 & n3294 ;
  assign n11049 = ~n6256 & n11048 ;
  assign n11050 = x0 & n8072 ;
  assign n11051 = n228 & n3018 ;
  assign n11052 = ~n24 & n11051 ;
  assign n11053 = ~n11050 & ~n11052 ;
  assign n11054 = ~n11049 & n11053 ;
  assign n11055 = ~n11047 & n11054 ;
  assign n11056 = n642 & ~n11055 ;
  assign n11057 = ~n11043 & ~n11056 ;
  assign n11058 = x7 & n11057 ;
  assign n11059 = ~n11008 & n11058 ;
  assign n11060 = n10941 & n11059 ;
  assign n11061 = n768 & n1551 ;
  assign n11062 = ~n1747 & ~n2709 ;
  assign n11063 = ~n1529 & n11062 ;
  assign n11064 = n10562 & n11063 ;
  assign n11065 = ~n11061 & ~n11064 ;
  assign n11066 = n3194 & ~n11065 ;
  assign n11067 = n2680 & n8471 ;
  assign n11068 = n426 & n3819 ;
  assign n11069 = n475 & n11068 ;
  assign n11070 = ~n11067 & ~n11069 ;
  assign n11071 = ~x0 & ~n11070 ;
  assign n11072 = n2124 & ~n6013 ;
  assign n11073 = ~n890 & ~n1366 ;
  assign n11074 = n10159 & ~n11073 ;
  assign n11075 = ~n1368 & ~n11074 ;
  assign n11076 = ~n11072 & n11075 ;
  assign n11077 = n9550 & ~n11076 ;
  assign n11078 = n1562 & n6101 ;
  assign n11079 = n1760 & n9509 ;
  assign n11080 = x15 & n11079 ;
  assign n11081 = ~n11078 & ~n11080 ;
  assign n11082 = ~n11077 & n11081 ;
  assign n11083 = n5270 & ~n11082 ;
  assign n11084 = ~n11071 & ~n11083 ;
  assign n11085 = ~n19 & n286 ;
  assign n11086 = ~n2709 & n11085 ;
  assign n11087 = ~n470 & ~n5897 ;
  assign n11088 = n33 & n10466 ;
  assign n11089 = ~n1511 & ~n11088 ;
  assign n11090 = ~n11087 & n11089 ;
  assign n11091 = n11090 ^ n10730 ;
  assign n11092 = n11091 ^ x10 ;
  assign n11100 = n11092 ^ n11091 ;
  assign n11093 = n753 & n1633 ;
  assign n11094 = n11093 ^ n11092 ;
  assign n11095 = n11094 ^ n11091 ;
  assign n11096 = n11092 ^ n11090 ;
  assign n11097 = n11096 ^ n11093 ;
  assign n11098 = n11097 ^ n11095 ;
  assign n11099 = ~n11095 & ~n11098 ;
  assign n11101 = n11100 ^ n11099 ;
  assign n11102 = n11101 ^ n11095 ;
  assign n11103 = n11091 ^ x8 ;
  assign n11104 = n11099 ^ n11095 ;
  assign n11105 = n11103 & ~n11104 ;
  assign n11106 = n11105 ^ n11091 ;
  assign n11107 = ~n11102 & ~n11106 ;
  assign n11108 = n11107 ^ n11091 ;
  assign n11109 = n11108 ^ n10730 ;
  assign n11110 = n11109 ^ n11091 ;
  assign n11111 = n210 & n11110 ;
  assign n11112 = ~n11086 & ~n11111 ;
  assign n11113 = x1 & ~n11112 ;
  assign n11114 = n11084 & ~n11113 ;
  assign n11115 = ~n11066 & n11114 ;
  assign n11116 = ~n1352 & ~n11115 ;
  assign n11117 = n2075 & n9460 ;
  assign n11118 = n2503 & n11117 ;
  assign n11119 = n11118 ^ x6 ;
  assign n11120 = ~x1 & n1718 ;
  assign n11121 = n585 & n11120 ;
  assign n11122 = ~n1394 & n11121 ;
  assign n11123 = x10 & n10784 ;
  assign n11124 = ~x8 & n2075 ;
  assign n11125 = n9550 & n11124 ;
  assign n11126 = ~n1698 & n11120 ;
  assign n11127 = ~n11125 & ~n11126 ;
  assign n11128 = ~n140 & ~n717 ;
  assign n11129 = ~n11127 & ~n11128 ;
  assign n11130 = ~n11123 & ~n11129 ;
  assign n11131 = ~n11122 & n11130 ;
  assign n11132 = n11131 ^ x9 ;
  assign n11133 = n11132 ^ n11131 ;
  assign n11134 = n1588 ^ x2 ;
  assign n11141 = n11134 ^ n1588 ;
  assign n11135 = n11134 ^ x8 ;
  assign n11136 = n11135 ^ n1588 ;
  assign n11137 = x10 ^ x8 ;
  assign n11138 = n11137 ^ x8 ;
  assign n11139 = n11138 ^ n11136 ;
  assign n11140 = ~n11136 & n11139 ;
  assign n11142 = n11141 ^ n11140 ;
  assign n11143 = n11142 ^ n11136 ;
  assign n11144 = n1588 ^ n504 ;
  assign n11145 = n11144 ^ n1588 ;
  assign n11146 = n11140 ^ n11136 ;
  assign n11147 = ~n11145 & ~n11146 ;
  assign n11148 = n11147 ^ n1588 ;
  assign n11149 = ~n11143 & n11148 ;
  assign n11150 = n11149 ^ n1588 ;
  assign n11151 = n11150 ^ n1588 ;
  assign n11152 = n11151 ^ n1588 ;
  assign n11153 = n318 & n11152 ;
  assign n11154 = ~n133 & ~n10944 ;
  assign n11155 = n11154 ^ x1 ;
  assign n11156 = n11154 ^ n10942 ;
  assign n11157 = n11156 ^ n10942 ;
  assign n11158 = ~n320 & n8868 ;
  assign n11159 = n11158 ^ n10942 ;
  assign n11160 = ~n11157 & ~n11159 ;
  assign n11161 = n11160 ^ n10942 ;
  assign n11162 = ~n11155 & n11161 ;
  assign n11163 = n11162 ^ x1 ;
  assign n11164 = ~n11153 & n11163 ;
  assign n11165 = n11164 ^ n11131 ;
  assign n11166 = n11133 & n11165 ;
  assign n11167 = n11166 ^ n11131 ;
  assign n11168 = n11167 ^ n11118 ;
  assign n11169 = ~n11119 & n11168 ;
  assign n11170 = n11169 ^ n11166 ;
  assign n11171 = n11170 ^ n11131 ;
  assign n11172 = n11171 ^ x6 ;
  assign n11173 = ~n11118 & ~n11172 ;
  assign n11174 = n11173 ^ n11118 ;
  assign n11175 = n11174 ^ n11118 ;
  assign n11176 = n278 & ~n11175 ;
  assign n11177 = n792 & n3649 ;
  assign n11178 = ~n17 & n2548 ;
  assign n11179 = ~n11123 & ~n11178 ;
  assign n11180 = n11177 & ~n11179 ;
  assign n11181 = ~n11176 & ~n11180 ;
  assign n11182 = n2257 & n6448 ;
  assign n11183 = ~n86 & n2225 ;
  assign n11184 = n1404 & n9048 ;
  assign n11185 = ~n11183 & ~n11184 ;
  assign n11186 = ~n1467 & ~n1706 ;
  assign n11187 = ~n1640 & n11186 ;
  assign n11188 = ~n890 & ~n11187 ;
  assign n11189 = ~x9 & n11188 ;
  assign n11190 = n11185 & ~n11189 ;
  assign n11191 = ~n3065 & n11190 ;
  assign n11192 = n3728 & ~n11191 ;
  assign n11193 = n3083 & n6721 ;
  assign n11194 = n10943 ^ x9 ;
  assign n11195 = n11194 ^ n10943 ;
  assign n11196 = n11195 ^ n11193 ;
  assign n11197 = n1283 & n1608 ;
  assign n11198 = n11197 ^ n343 ;
  assign n11199 = n343 & n11198 ;
  assign n11200 = n11199 ^ n10943 ;
  assign n11201 = n11200 ^ n343 ;
  assign n11202 = n11196 & n11201 ;
  assign n11203 = n11202 ^ n11199 ;
  assign n11204 = n11203 ^ n343 ;
  assign n11205 = ~n11193 & n11204 ;
  assign n11206 = n11205 ^ n11193 ;
  assign n11207 = ~n11192 & ~n11206 ;
  assign n11208 = ~n11182 & n11207 ;
  assign n11209 = n8009 & ~n11208 ;
  assign n11210 = n2156 & n9533 ;
  assign n11211 = n8666 & n11210 ;
  assign n11212 = ~n11209 & ~n11211 ;
  assign n11213 = ~x14 & n9337 ;
  assign n11214 = ~n9115 & ~n11213 ;
  assign n11215 = n6421 & ~n11214 ;
  assign n11216 = n4801 & n9093 ;
  assign n11217 = n310 & n2181 ;
  assign n11218 = ~n11216 & ~n11217 ;
  assign n11219 = n1528 & ~n11218 ;
  assign n11220 = n1758 & ~n10476 ;
  assign n11221 = n6923 & n11220 ;
  assign n11222 = ~n3808 & ~n9546 ;
  assign n11223 = ~n470 & n2410 ;
  assign n11224 = ~n11222 & n11223 ;
  assign n11225 = ~n11221 & ~n11224 ;
  assign n11226 = ~n11219 & n11225 ;
  assign n11227 = ~n11215 & n11226 ;
  assign n11228 = n10642 & ~n11227 ;
  assign n11229 = n9199 & n9557 ;
  assign n11230 = n2277 & n11229 ;
  assign n11231 = n692 ^ x2 ;
  assign n11232 = n1303 & n7418 ;
  assign n11233 = ~n10943 & ~n11232 ;
  assign n11234 = ~n8455 & n11233 ;
  assign n11235 = n11234 ^ n11231 ;
  assign n11236 = n11235 ^ n692 ;
  assign n11237 = n11236 ^ n11235 ;
  assign n11238 = n1551 & n2705 ;
  assign n11239 = n1454 & n11238 ;
  assign n11240 = n11239 ^ n11235 ;
  assign n11241 = n11240 ^ n11231 ;
  assign n11242 = n11237 & n11241 ;
  assign n11243 = n11242 ^ n11239 ;
  assign n11244 = n10858 & ~n11239 ;
  assign n11245 = n11244 ^ n11231 ;
  assign n11246 = ~n11243 & ~n11245 ;
  assign n11247 = n11246 ^ n11244 ;
  assign n11248 = ~n11231 & n11247 ;
  assign n11249 = n11248 ^ n11242 ;
  assign n11250 = n11249 ^ x2 ;
  assign n11251 = n11250 ^ n11239 ;
  assign n11252 = ~n11230 & n11251 ;
  assign n11253 = x6 & ~n11252 ;
  assign n11254 = ~x2 & ~n10302 ;
  assign n11255 = ~n9891 & ~n11254 ;
  assign n11256 = n8282 & ~n11255 ;
  assign n11257 = ~n11253 & ~n11256 ;
  assign n11258 = n792 & ~n11257 ;
  assign n11259 = ~n11228 & ~n11258 ;
  assign n11260 = n11212 & n11259 ;
  assign n11261 = n11181 & n11260 ;
  assign n11262 = ~n11116 & n11261 ;
  assign n11263 = ~x5 & ~n11262 ;
  assign n11264 = n20 & n5669 ;
  assign n11265 = ~x1 & n1702 ;
  assign n11266 = ~n222 & n11265 ;
  assign n11267 = n107 & n799 ;
  assign n11268 = ~n295 & n816 ;
  assign n11269 = ~n1622 & n11268 ;
  assign n11270 = ~n11267 & ~n11269 ;
  assign n11271 = ~x0 & ~n2691 ;
  assign n11272 = ~n5021 & ~n11271 ;
  assign n11273 = n263 & ~n11272 ;
  assign n11274 = n11270 & ~n11273 ;
  assign n11275 = ~n11266 & n11274 ;
  assign n11276 = n267 & ~n11275 ;
  assign n11277 = n210 & ~n1027 ;
  assign n11278 = ~n2660 & n11277 ;
  assign n11279 = ~n6067 & ~n11278 ;
  assign n11280 = x14 & n1254 ;
  assign n11281 = ~n11279 & n11280 ;
  assign n11282 = n132 & n221 ;
  assign n11283 = n3991 & n11282 ;
  assign n11284 = ~n11281 & ~n11283 ;
  assign n11285 = ~n11276 & n11284 ;
  assign n11286 = ~n11264 & n11285 ;
  assign n11287 = n1483 & ~n11286 ;
  assign n11288 = x1 & n3317 ;
  assign n11289 = n20 & n5636 ;
  assign n11290 = ~n11288 & ~n11289 ;
  assign n11291 = n1518 & ~n11290 ;
  assign n11292 = n3226 & n11291 ;
  assign n11293 = n245 & n6670 ;
  assign n11294 = n24 & n1551 ;
  assign n11295 = ~n11293 & ~n11294 ;
  assign n11296 = n3317 & ~n11295 ;
  assign n11297 = ~n269 & ~n1702 ;
  assign n11298 = ~n2331 & ~n3048 ;
  assign n11299 = ~n7087 & n11298 ;
  assign n11300 = ~n291 & ~n5733 ;
  assign n11301 = ~n1285 & ~n11277 ;
  assign n11302 = n11300 & n11301 ;
  assign n11303 = x1 & ~n1435 ;
  assign n11304 = ~n3249 & n11303 ;
  assign n11305 = ~n533 & ~n11304 ;
  assign n11306 = n11302 & ~n11305 ;
  assign n11307 = n11299 & n11306 ;
  assign n11308 = ~n11297 & n11307 ;
  assign n11309 = ~n11296 & ~n11308 ;
  assign n11310 = n5647 & ~n11309 ;
  assign n11311 = n2687 & n11120 ;
  assign n11312 = n86 & n5344 ;
  assign n11313 = n11311 & n11312 ;
  assign n11314 = ~n11310 & ~n11313 ;
  assign n11315 = ~n11292 & n11314 ;
  assign n11316 = ~n11287 & n11315 ;
  assign n11317 = x15 & ~n11316 ;
  assign n11318 = n266 & n6693 ;
  assign n11319 = n1234 & n10942 ;
  assign n11320 = ~n8868 & ~n10979 ;
  assign n11321 = n792 & ~n11320 ;
  assign n11322 = ~n11319 & ~n11321 ;
  assign n11323 = ~n11318 & n11322 ;
  assign n11324 = n11323 ^ x2 ;
  assign n11325 = n11324 ^ n11323 ;
  assign n11326 = ~x1 & n1394 ;
  assign n11327 = n7853 & n11326 ;
  assign n11328 = n11327 ^ n11323 ;
  assign n11329 = n11328 ^ n11323 ;
  assign n11330 = ~n11325 & n11329 ;
  assign n11331 = n11330 ^ n11323 ;
  assign n11332 = x5 & ~n11331 ;
  assign n11333 = n11332 ^ n11323 ;
  assign n11334 = n205 & ~n11333 ;
  assign n11335 = ~n5222 & ~n11124 ;
  assign n11336 = n1260 & n2102 ;
  assign n11337 = ~n11335 & n11336 ;
  assign n11338 = n2352 & n11327 ;
  assign n11339 = n1483 & n11177 ;
  assign n11340 = n1834 & n11339 ;
  assign n11341 = ~n11338 & ~n11340 ;
  assign n11342 = ~n11337 & n11341 ;
  assign n11343 = ~n11334 & n11342 ;
  assign n11344 = n11343 ^ x14 ;
  assign n11345 = n11344 ^ n11343 ;
  assign n11346 = n11345 ^ n11317 ;
  assign n11347 = n1620 & n5270 ;
  assign n11348 = n1623 & n1715 ;
  assign n11349 = n2405 & n11293 ;
  assign n11350 = ~n11348 & ~n11349 ;
  assign n11351 = n450 & ~n11320 ;
  assign n11352 = n11350 & ~n11351 ;
  assign n11353 = n1261 & ~n11352 ;
  assign n11354 = ~n11347 & ~n11353 ;
  assign n11355 = n11354 ^ x6 ;
  assign n11356 = ~x6 & n11355 ;
  assign n11357 = n11356 ^ n11343 ;
  assign n11358 = n11357 ^ x6 ;
  assign n11359 = ~n11346 & n11358 ;
  assign n11360 = n11359 ^ n11356 ;
  assign n11361 = n11360 ^ x6 ;
  assign n11362 = ~n11317 & ~n11361 ;
  assign n11363 = n11362 ^ n11317 ;
  assign n11364 = ~n2169 & n11363 ;
  assign n11365 = n1658 & n4402 ;
  assign n11366 = n2352 & n11365 ;
  assign n11367 = n2680 & n6067 ;
  assign n11368 = n228 & n2639 ;
  assign n11369 = ~n11367 & ~n11368 ;
  assign n11370 = x15 & n6617 ;
  assign n11371 = ~n11369 & n11370 ;
  assign n11372 = n2445 & n2656 ;
  assign n11373 = n1404 & n2647 ;
  assign n11374 = ~n11372 & ~n11373 ;
  assign n11375 = ~x5 & ~n11374 ;
  assign n11376 = ~x1 & n222 ;
  assign n11377 = n4536 & n11376 ;
  assign n11378 = ~n11375 & ~n11377 ;
  assign n11379 = ~n470 & n8748 ;
  assign n11380 = ~n11378 & n11379 ;
  assign n11381 = ~n11371 & ~n11380 ;
  assign n11382 = ~n11366 & n11381 ;
  assign n11383 = ~n3552 & ~n11382 ;
  assign n11384 = n1597 ^ n692 ;
  assign n11385 = n1502 & ~n3161 ;
  assign n11386 = ~n1027 & n11385 ;
  assign n11387 = n11386 ^ n2075 ;
  assign n11388 = n11386 ^ n5544 ;
  assign n11389 = n11388 ^ n5544 ;
  assign n11390 = n11389 ^ n11387 ;
  assign n11391 = n3659 ^ n394 ;
  assign n11392 = n394 & n11391 ;
  assign n11393 = n11392 ^ n5544 ;
  assign n11394 = n11393 ^ n394 ;
  assign n11395 = ~n11390 & ~n11394 ;
  assign n11396 = n11395 ^ n11392 ;
  assign n11397 = n11396 ^ n394 ;
  assign n11398 = n11387 & n11397 ;
  assign n11399 = n11398 ^ n11386 ;
  assign n11400 = n11399 ^ n11384 ;
  assign n11401 = n11400 ^ n692 ;
  assign n11402 = n11401 ^ n11400 ;
  assign n11403 = n1670 & n1979 ;
  assign n11404 = n291 & n1252 ;
  assign n11405 = ~n10190 & ~n11404 ;
  assign n11406 = n2038 & ~n11405 ;
  assign n11407 = n2503 & n8232 ;
  assign n11408 = ~n11406 & ~n11407 ;
  assign n11409 = ~n11403 & n11408 ;
  assign n11410 = n11409 ^ n11400 ;
  assign n11411 = n11410 ^ n11384 ;
  assign n11412 = n11402 & n11411 ;
  assign n11413 = n11412 ^ n11409 ;
  assign n11414 = ~x1 & n10992 ;
  assign n11415 = n394 & ~n2278 ;
  assign n11416 = ~n11414 & n11415 ;
  assign n11417 = ~n4951 & ~n11416 ;
  assign n11418 = n11409 & n11417 ;
  assign n11419 = n11418 ^ n11384 ;
  assign n11420 = n11413 & ~n11419 ;
  assign n11421 = n11420 ^ n11418 ;
  assign n11422 = ~n11384 & n11421 ;
  assign n11423 = n11422 ^ n11412 ;
  assign n11424 = n11423 ^ n1597 ;
  assign n11425 = n11424 ^ n11409 ;
  assign n11426 = ~n11383 & ~n11425 ;
  assign n11427 = ~x7 & n11426 ;
  assign n11428 = ~n11364 & n11427 ;
  assign n11429 = n11428 ^ n11263 ;
  assign n11430 = n679 & n8666 ;
  assign n11431 = n2156 & n11430 ;
  assign n11460 = ~n1529 & n2565 ;
  assign n11461 = n11460 ^ n7857 ;
  assign n11462 = n11461 ^ n11460 ;
  assign n11463 = ~x9 & n62 ;
  assign n11464 = x8 & n11463 ;
  assign n11465 = n11464 ^ n11460 ;
  assign n11466 = n11465 ^ n11460 ;
  assign n11467 = ~n11462 & ~n11466 ;
  assign n11468 = n11467 ^ n11460 ;
  assign n11469 = x2 & ~n11468 ;
  assign n11470 = n11469 ^ n11460 ;
  assign n11432 = n3246 & n7549 ;
  assign n11433 = ~n4327 & ~n9354 ;
  assign n11434 = n2282 & ~n11433 ;
  assign n11435 = n2005 & n6397 ;
  assign n11436 = ~n11434 & ~n11435 ;
  assign n11437 = ~n11432 & n11436 ;
  assign n11438 = x13 & ~n11437 ;
  assign n11439 = n1368 & n1643 ;
  assign n11440 = n153 & n2586 ;
  assign n11441 = n2776 & n11440 ;
  assign n11442 = ~n11439 & ~n11441 ;
  assign n11443 = ~n603 & n1539 ;
  assign n11444 = n3521 & n11443 ;
  assign n11445 = n11442 & ~n11444 ;
  assign n11446 = n284 & n2005 ;
  assign n11447 = ~n1394 & n11446 ;
  assign n11448 = n281 & n1365 ;
  assign n11449 = ~n8577 & ~n11448 ;
  assign n11450 = n286 & ~n11449 ;
  assign n11451 = n9650 & n9832 ;
  assign n11452 = ~n5896 & ~n11451 ;
  assign n11453 = ~n11450 & n11452 ;
  assign n11454 = ~n11447 & n11453 ;
  assign n11455 = ~n1352 & ~n11454 ;
  assign n11456 = n11445 & ~n11455 ;
  assign n11457 = ~n11438 & n11456 ;
  assign n11471 = n11470 ^ n11457 ;
  assign n11472 = n11471 ^ n11457 ;
  assign n11458 = n11457 ^ n1352 ;
  assign n11459 = n11458 ^ n11457 ;
  assign n11473 = n11472 ^ n11459 ;
  assign n11474 = n11457 ^ x13 ;
  assign n11475 = n11474 ^ n11457 ;
  assign n11476 = n11475 ^ n11472 ;
  assign n11477 = n11472 & ~n11476 ;
  assign n11478 = n11477 ^ n11472 ;
  assign n11479 = ~n11473 & n11478 ;
  assign n11480 = n11479 ^ n11477 ;
  assign n11481 = n11480 ^ n11457 ;
  assign n11482 = n11481 ^ n11472 ;
  assign n11483 = x1 & ~n11482 ;
  assign n11484 = n11483 ^ n11457 ;
  assign n11485 = ~n11431 & n11484 ;
  assign n11486 = x15 & ~n11485 ;
  assign n11487 = x1 & n2257 ;
  assign n11488 = n71 & n11487 ;
  assign n11489 = ~n43 & ~n4376 ;
  assign n11490 = n1376 & n11489 ;
  assign n11491 = ~n11488 & ~n11490 ;
  assign n11492 = ~n1370 & ~n11491 ;
  assign n11493 = ~n533 & ~n880 ;
  assign n11494 = n214 & ~n11493 ;
  assign n11495 = n3233 & n11494 ;
  assign n11496 = ~x5 & ~n11495 ;
  assign n11497 = n2871 & n3508 ;
  assign n11498 = n3068 & ~n5678 ;
  assign n11499 = ~n1979 & ~n4313 ;
  assign n11500 = ~n11498 & n11499 ;
  assign n11501 = ~x8 & ~n11500 ;
  assign n11502 = ~n11497 & ~n11501 ;
  assign n11503 = n1376 & ~n11502 ;
  assign n11504 = n1511 & n4134 ;
  assign n11505 = x1 & ~n5678 ;
  assign n11506 = x13 & ~n3264 ;
  assign n11507 = ~n11505 & ~n11506 ;
  assign n11508 = n3056 & ~n11507 ;
  assign n11509 = ~n4498 & ~n4505 ;
  assign n11510 = n249 & ~n11509 ;
  assign n11511 = ~n11508 & ~n11510 ;
  assign n11512 = n1252 & ~n11511 ;
  assign n11513 = ~n11504 & ~n11512 ;
  assign n11514 = ~n11503 & n11513 ;
  assign n11515 = n11496 & n11514 ;
  assign n11516 = ~n11492 & n11515 ;
  assign n11517 = ~n11486 & n11516 ;
  assign n11518 = n532 & ~n2006 ;
  assign n11519 = ~x12 & n9832 ;
  assign n11520 = ~x2 & ~n2042 ;
  assign n11521 = ~n11519 & ~n11520 ;
  assign n11522 = ~n11518 & n11521 ;
  assign n11523 = n291 & ~n11522 ;
  assign n11524 = n4423 ^ n926 ;
  assign n11525 = n11524 ^ n4423 ;
  assign n11526 = n4423 ^ n475 ;
  assign n11527 = n11526 ^ n4423 ;
  assign n11528 = n11525 & n11527 ;
  assign n11529 = n11528 ^ n4423 ;
  assign n11530 = ~x6 & ~n11529 ;
  assign n11531 = n11530 ^ n4423 ;
  assign n11532 = ~n2006 & ~n11531 ;
  assign n11533 = ~n2233 & n11505 ;
  assign n11534 = n2483 & n4423 ;
  assign n11535 = n11533 & n11534 ;
  assign n11536 = ~n11532 & ~n11535 ;
  assign n11537 = n1330 & ~n11536 ;
  assign n11538 = ~n2387 & ~n3048 ;
  assign n11539 = n943 & ~n11538 ;
  assign n11540 = ~n2548 & ~n4275 ;
  assign n11541 = ~n11539 & n11540 ;
  assign n11542 = n394 & ~n11541 ;
  assign n11543 = ~n11537 & ~n11542 ;
  assign n11544 = ~n11523 & n11543 ;
  assign n11545 = ~x8 & ~n11544 ;
  assign n11546 = n214 & n426 ;
  assign n11547 = ~n228 & ~n2397 ;
  assign n11548 = n11546 & n11547 ;
  assign n11549 = n1581 & ~n11548 ;
  assign n11550 = n2038 & n9580 ;
  assign n11551 = n11550 ^ n11548 ;
  assign n11552 = n167 & n11505 ;
  assign n11553 = n11552 ^ n11549 ;
  assign n11554 = n11551 & n11553 ;
  assign n11555 = n11554 ^ n11552 ;
  assign n11556 = n11549 & n11555 ;
  assign n11557 = n11556 ^ n11548 ;
  assign n11558 = n11557 ^ n1506 ;
  assign n11559 = n11558 ^ n11557 ;
  assign n11560 = ~n334 & n396 ;
  assign n11561 = ~n3967 & ~n8973 ;
  assign n11562 = ~n11560 & ~n11561 ;
  assign n11563 = n11562 ^ n11557 ;
  assign n11564 = n11563 ^ n11557 ;
  assign n11565 = n11559 & n11564 ;
  assign n11566 = n11565 ^ n11557 ;
  assign n11567 = ~x6 & n11566 ;
  assign n11568 = n11567 ^ n11557 ;
  assign n11569 = ~n11545 & ~n11568 ;
  assign n11570 = x5 & n11569 ;
  assign n11571 = ~n11517 & ~n11570 ;
  assign n11572 = n394 & n2075 ;
  assign n11573 = n10410 & n11572 ;
  assign n11574 = n3740 & n5124 ;
  assign n11575 = n396 & n1671 ;
  assign n11576 = n222 & n11575 ;
  assign n11577 = ~n11574 & ~n11576 ;
  assign n11578 = n679 & ~n11577 ;
  assign n11579 = ~n4505 & ~n7407 ;
  assign n11580 = n817 & ~n2276 ;
  assign n11581 = n5124 & n11580 ;
  assign n11582 = ~n11579 & n11581 ;
  assign n11583 = ~n11578 & ~n11582 ;
  assign n11584 = ~n2905 & ~n11583 ;
  assign n11585 = ~n11573 & ~n11584 ;
  assign n11586 = ~n11571 & n11585 ;
  assign n11587 = ~x10 & ~n11586 ;
  assign n11588 = n291 & n9759 ;
  assign n11589 = n394 & ~n9900 ;
  assign n11590 = ~n11588 & ~n11589 ;
  assign n11591 = n10895 & ~n11590 ;
  assign n11592 = ~n7492 & ~n8494 ;
  assign n11593 = ~x9 & ~n11592 ;
  assign n11594 = ~n2503 & ~n11593 ;
  assign n11595 = n247 & ~n11594 ;
  assign n11596 = n1657 & n3453 ;
  assign n11597 = ~n1404 & ~n11596 ;
  assign n11598 = ~n7001 & ~n11597 ;
  assign n11599 = ~n7988 & n11598 ;
  assign n11600 = n3728 & n11599 ;
  assign n11601 = n167 & n1454 ;
  assign n11602 = ~n49 & ~n11601 ;
  assign n11603 = n4878 & ~n11602 ;
  assign n11604 = ~n11600 & ~n11603 ;
  assign n11605 = n2483 & n3658 ;
  assign n11606 = n3673 & n9389 ;
  assign n11607 = n1669 & ~n11606 ;
  assign n11608 = ~n476 & ~n3069 ;
  assign n11609 = n133 & ~n11608 ;
  assign n11610 = n1503 & ~n11609 ;
  assign n11611 = ~n11607 & ~n11610 ;
  assign n11612 = ~n11605 & n11611 ;
  assign n11613 = n228 & ~n11612 ;
  assign n11614 = n2445 & n10312 ;
  assign n11615 = ~n460 & ~n11614 ;
  assign n11616 = n11597 & n11615 ;
  assign n11617 = n5545 & ~n11616 ;
  assign n11618 = ~n11613 & ~n11617 ;
  assign n11619 = n11604 & n11618 ;
  assign n11620 = ~n11595 & n11619 ;
  assign n11621 = ~x5 & ~n11620 ;
  assign n11622 = n3453 & ~n9428 ;
  assign n11623 = n3967 & ~n11622 ;
  assign n11624 = ~n11035 & ~n11623 ;
  assign n11625 = n1670 & ~n11624 ;
  assign n11626 = ~n11621 & ~n11625 ;
  assign n11627 = ~n11591 & n11626 ;
  assign n11628 = n6670 & ~n11627 ;
  assign n11629 = n1138 & n8981 ;
  assign n11630 = n200 & n1618 ;
  assign n11631 = ~n6611 & ~n11630 ;
  assign n11632 = n570 & n4691 ;
  assign n11633 = ~n11631 & n11632 ;
  assign n11634 = ~n11629 & ~n11633 ;
  assign n11635 = n266 & ~n11634 ;
  assign n11636 = n1633 & ~n2483 ;
  assign n11637 = n5465 & n11636 ;
  assign n11638 = n396 & n1457 ;
  assign n11639 = n11637 & n11638 ;
  assign n11640 = ~n1322 & n11639 ;
  assign n11641 = ~n11635 & ~n11640 ;
  assign n11642 = ~n11628 & n11641 ;
  assign n11643 = ~n1394 & ~n9092 ;
  assign n11644 = n1138 & ~n11643 ;
  assign n11645 = ~n1528 & n6611 ;
  assign n11646 = ~n9020 & ~n11645 ;
  assign n11647 = n425 & n5647 ;
  assign n11648 = ~n504 & n11647 ;
  assign n11649 = n11646 & ~n11648 ;
  assign n11650 = ~n11644 & n11649 ;
  assign n11651 = x9 & ~n11650 ;
  assign n11652 = ~n42 & ~n3249 ;
  assign n11653 = n2218 & ~n11652 ;
  assign n11654 = ~n5897 & n11653 ;
  assign n11655 = n190 & n1366 ;
  assign n11656 = ~n2289 & n11655 ;
  assign n11657 = ~n11654 & ~n11656 ;
  assign n11658 = ~n11651 & n11657 ;
  assign n11659 = n266 & ~n11658 ;
  assign n11660 = n2105 & n2282 ;
  assign n11661 = x9 & n3729 ;
  assign n11662 = ~n267 & n2277 ;
  assign n11663 = ~n11661 & ~n11662 ;
  assign n11664 = ~n11660 & n11663 ;
  assign n11665 = n49 & ~n11664 ;
  assign n11666 = n49 & ~n2282 ;
  assign n11667 = ~n3282 & ~n11666 ;
  assign n11668 = n267 & n5919 ;
  assign n11669 = ~n11667 & n11668 ;
  assign n11670 = n425 & n603 ;
  assign n11671 = n2397 & n11670 ;
  assign n11672 = ~n11669 & ~n11671 ;
  assign n11673 = ~n890 & ~n6000 ;
  assign n11674 = n2483 & ~n11673 ;
  assign n11675 = n11674 ^ x2 ;
  assign n11676 = n11675 ^ n11674 ;
  assign n11677 = n11676 ^ n11672 ;
  assign n11678 = n49 & n2739 ;
  assign n11679 = ~n9551 & ~n11678 ;
  assign n11680 = n11679 ^ x6 ;
  assign n11681 = ~n11679 & n11680 ;
  assign n11682 = n11681 ^ n11674 ;
  assign n11683 = n11682 ^ n11679 ;
  assign n11684 = ~n11677 & ~n11683 ;
  assign n11685 = n11684 ^ n11681 ;
  assign n11686 = n11685 ^ n11679 ;
  assign n11687 = n11672 & ~n11686 ;
  assign n11688 = n11687 ^ n11672 ;
  assign n11689 = x15 & ~n11688 ;
  assign n11690 = n286 & n9655 ;
  assign n11691 = ~n11689 & ~n11690 ;
  assign n11692 = ~n11665 & n11691 ;
  assign n11693 = n1456 & ~n11692 ;
  assign n11694 = n280 & n1503 ;
  assign n11695 = n9291 & n11694 ;
  assign n11696 = ~n2469 & ~n2945 ;
  assign n11697 = ~n2156 & ~n11696 ;
  assign n11698 = n9306 & ~n11673 ;
  assign n11699 = ~n11697 & ~n11698 ;
  assign n11700 = ~n9779 & n11699 ;
  assign n11701 = ~n891 & n1657 ;
  assign n11702 = ~n11678 & ~n11701 ;
  assign n11703 = ~x9 & ~n11702 ;
  assign n11704 = n9337 & n10179 ;
  assign n11705 = ~n11703 & ~n11704 ;
  assign n11706 = ~n9874 & n11705 ;
  assign n11707 = n1254 & ~n11706 ;
  assign n11708 = n11700 & ~n11707 ;
  assign n11709 = n247 & ~n11708 ;
  assign n11710 = ~n11695 & ~n11709 ;
  assign n11711 = ~n153 & n2277 ;
  assign n11712 = n2397 & n10312 ;
  assign n11713 = ~n4506 & ~n11712 ;
  assign n11714 = ~n11596 & n11713 ;
  assign n11715 = ~n11711 & n11714 ;
  assign n11716 = n2483 & ~n11715 ;
  assign n11717 = n4690 ^ n2503 ;
  assign n11718 = ~x2 & n11717 ;
  assign n11719 = n11718 ^ n4690 ;
  assign n11720 = ~n11716 & ~n11719 ;
  assign n11721 = n222 & ~n11720 ;
  assign n11722 = n11710 & ~n11721 ;
  assign n11723 = ~n11693 & n11722 ;
  assign n11724 = ~n11659 & n11723 ;
  assign n11725 = n4746 & ~n11724 ;
  assign n11726 = n7087 & n10349 ;
  assign n11727 = ~n8984 & ~n9291 ;
  assign n11728 = n221 & ~n11727 ;
  assign n11729 = x6 & n11728 ;
  assign n11730 = ~n11726 & ~n11729 ;
  assign n11731 = n9884 & ~n11730 ;
  assign n11732 = ~n11725 & ~n11731 ;
  assign n11733 = n11642 & n11732 ;
  assign n11734 = ~n11587 & n11733 ;
  assign n11735 = n11734 ^ x0 ;
  assign n11736 = n11735 ^ n11734 ;
  assign n11737 = ~x6 & n1264 ;
  assign n11738 = ~n11009 & ~n11737 ;
  assign n11739 = n2075 & ~n11738 ;
  assign n11740 = n1511 & n11739 ;
  assign n11741 = n792 & n1671 ;
  assign n11742 = n8048 & n11741 ;
  assign n11743 = n1493 & n6670 ;
  assign n11744 = ~n1438 & n11743 ;
  assign n11745 = n585 & ~n2225 ;
  assign n11746 = n1698 & n11745 ;
  assign n11747 = n11746 ^ x1 ;
  assign n11748 = n11747 ^ n11746 ;
  assign n11749 = n11748 ^ x4 ;
  assign n11750 = n1435 ^ x8 ;
  assign n11751 = ~n1435 & ~n11750 ;
  assign n11752 = n11751 ^ n11746 ;
  assign n11753 = n11752 ^ n1435 ;
  assign n11754 = ~n11749 & n11753 ;
  assign n11755 = n11754 ^ n11751 ;
  assign n11756 = n11755 ^ n1435 ;
  assign n11757 = ~x4 & ~n11756 ;
  assign n11758 = n11757 ^ x4 ;
  assign n11759 = ~n11744 & n11758 ;
  assign n11760 = n1290 & ~n11759 ;
  assign n11761 = n38 & n11741 ;
  assign n11762 = ~n119 & ~n1581 ;
  assign n11763 = n2424 & ~n11762 ;
  assign n11764 = n284 & n1633 ;
  assign n11765 = n5403 & n11764 ;
  assign n11766 = ~n11763 & ~n11765 ;
  assign n11767 = n1275 & ~n11766 ;
  assign n11768 = ~n49 & n504 ;
  assign n11769 = n1670 & ~n11768 ;
  assign n11770 = n258 & n11769 ;
  assign n11771 = ~x10 & n11770 ;
  assign n11772 = ~n11767 & ~n11771 ;
  assign n11773 = ~n11761 & n11772 ;
  assign n11774 = ~n11760 & n11773 ;
  assign n11775 = ~n11742 & n11774 ;
  assign n11776 = n2005 & ~n11775 ;
  assign n11777 = n1642 & n9533 ;
  assign n11778 = n11376 & n11777 ;
  assign n11779 = n291 & ~n1562 ;
  assign n11780 = ~n8172 & ~n11779 ;
  assign n11781 = x1 & ~n11780 ;
  assign n11782 = n6817 ^ n1598 ;
  assign n11783 = n11782 ^ n1598 ;
  assign n11784 = n11783 ^ x12 ;
  assign n11785 = n11782 ^ x4 ;
  assign n11786 = n11785 ^ n11783 ;
  assign n11787 = n11786 ^ n11784 ;
  assign n11788 = ~n11784 & n11787 ;
  assign n11789 = n11788 ^ n11782 ;
  assign n11790 = n11789 ^ n11784 ;
  assign n11791 = n11782 ^ x15 ;
  assign n11792 = ~n11783 & n11791 ;
  assign n11793 = n11792 ^ n11782 ;
  assign n11794 = n11790 & ~n11793 ;
  assign n11795 = n11794 ^ n11782 ;
  assign n11796 = n11795 ^ n1598 ;
  assign n11797 = ~x13 & n11796 ;
  assign n11798 = n11781 & ~n11797 ;
  assign n11799 = ~n2289 & n10413 ;
  assign n11800 = ~n11798 & ~n11799 ;
  assign n11801 = n295 & ~n11800 ;
  assign n11802 = n1597 & n3728 ;
  assign n11803 = n1395 ^ x4 ;
  assign n11804 = n11803 ^ n1395 ;
  assign n11805 = n1395 ^ x8 ;
  assign n11806 = n11805 ^ n11803 ;
  assign n11807 = n11806 ^ x1 ;
  assign n11813 = n11807 ^ n11803 ;
  assign n11814 = n11813 ^ n1395 ;
  assign n11808 = n11807 ^ n9160 ;
  assign n11809 = n11808 ^ x1 ;
  assign n11810 = n11809 ^ n11808 ;
  assign n11811 = n11810 ^ n1395 ;
  assign n11812 = n11811 ^ n11804 ;
  assign n11815 = n11814 ^ n11812 ;
  assign n11816 = n11804 & n11815 ;
  assign n11817 = n11816 ^ n11810 ;
  assign n11818 = n11817 ^ n11814 ;
  assign n11823 = n11808 ^ n11807 ;
  assign n11819 = n11808 ^ n9462 ;
  assign n11820 = n11814 ^ n11810 ;
  assign n11821 = ~n11819 & n11820 ;
  assign n11822 = n11821 ^ n11816 ;
  assign n11824 = n11823 ^ n11822 ;
  assign n11825 = n11824 ^ n11819 ;
  assign n11826 = n11825 ^ n11810 ;
  assign n11827 = n11814 & ~n11826 ;
  assign n11828 = n11827 ^ n11804 ;
  assign n11829 = n11818 & n11828 ;
  assign n11830 = n11829 ^ n11804 ;
  assign n11831 = n11830 ^ x4 ;
  assign n11832 = n11831 ^ n11804 ;
  assign n11833 = n11802 & n11832 ;
  assign n11834 = ~n11801 & ~n11833 ;
  assign n11835 = ~n11778 & n11834 ;
  assign n11836 = ~x9 & ~n11835 ;
  assign n11837 = ~n11776 & ~n11836 ;
  assign n11838 = ~n11740 & n11837 ;
  assign n11839 = n11838 ^ n11734 ;
  assign n11840 = ~n11736 & n11839 ;
  assign n11841 = n11840 ^ n11734 ;
  assign n11842 = n11841 ^ n11263 ;
  assign n11843 = ~n11429 & ~n11842 ;
  assign n11844 = n11843 ^ n11840 ;
  assign n11845 = n11844 ^ n11734 ;
  assign n11846 = n11845 ^ n11428 ;
  assign n11847 = ~n11263 & n11846 ;
  assign n11848 = n11847 ^ n11263 ;
  assign n11849 = ~n11060 & n11848 ;
  assign n11850 = ~n399 & n3018 ;
  assign n11851 = ~n504 & n3821 ;
  assign n11852 = n11850 & n11851 ;
  assign n11853 = n343 & n5021 ;
  assign n11854 = n8020 & n11853 ;
  assign n11855 = n6824 & n9075 ;
  assign n11856 = n3896 & n11855 ;
  assign n11857 = ~n11854 & ~n11856 ;
  assign n11858 = ~n11852 & n11857 ;
  assign n11859 = n10719 ^ x13 ;
  assign n11860 = n11859 ^ n10719 ;
  assign n11861 = n10719 ^ n431 ;
  assign n11862 = n11861 ^ n10719 ;
  assign n11863 = ~n11860 & n11862 ;
  assign n11864 = n11863 ^ n10719 ;
  assign n11865 = x1 & ~n11864 ;
  assign n11866 = n11865 ^ n10719 ;
  assign n11867 = ~n11858 & ~n11866 ;
  assign n11868 = n3896 & n8573 ;
  assign n11869 = n3661 & n5961 ;
  assign n11870 = ~n11868 & ~n11869 ;
  assign n11871 = ~x1 & n5465 ;
  assign n11872 = ~n5264 & ~n11871 ;
  assign n11873 = ~n11870 & ~n11872 ;
  assign n11874 = ~n11867 & ~n11873 ;
  assign n11875 = ~n11849 & n11874 ;
  assign n11876 = ~n10718 & n11875 ;
  assign n11877 = n11876 ^ n10679 ;
  assign n11878 = n10681 & n11877 ;
  assign n11879 = n11878 ^ n10679 ;
  assign n11880 = n8967 & n11879 ;
  assign n11881 = n11880 ^ n8841 ;
  assign n11882 = n8843 & n11881 ;
  assign n11883 = n11882 ^ n8841 ;
  assign n11884 = n5709 & n11883 ;
  assign y0 = ~n11884 ;
endmodule
