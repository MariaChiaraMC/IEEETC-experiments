module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 ;
  assign n8 = ~x1 & ~x5 ;
  assign n9 = x3 & ~n8 ;
  assign n7 = ~x0 & x2 ;
  assign n10 = n9 ^ n7 ;
  assign n11 = n10 ^ n7 ;
  assign n12 = x0 & ~x5 ;
  assign n13 = x0 & ~x1 ;
  assign n14 = x2 & n13 ;
  assign n15 = ~n12 & ~n14 ;
  assign n16 = n15 ^ n7 ;
  assign n17 = n11 & ~n16 ;
  assign n18 = n17 ^ n7 ;
  assign n19 = x4 & n18 ;
  assign n20 = x1 ^ x0 ;
  assign n23 = x5 ^ x4 ;
  assign n21 = x5 ^ x3 ;
  assign n22 = n21 ^ x4 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ n20 ;
  assign n26 = n20 & ~n25 ;
  assign n27 = n26 ^ x5 ;
  assign n28 = n27 ^ n20 ;
  assign n29 = x1 & ~n22 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = n28 & n30 ;
  assign n32 = n31 ^ x5 ;
  assign n33 = n32 ^ x2 ;
  assign n34 = n33 ^ n32 ;
  assign n35 = n34 ^ n19 ;
  assign n36 = ~x1 & ~x3 ;
  assign n37 = n36 ^ n12 ;
  assign n38 = n12 & n37 ;
  assign n39 = n38 ^ n32 ;
  assign n40 = n39 ^ n12 ;
  assign n41 = ~n35 & n40 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = n42 ^ n12 ;
  assign n44 = ~n19 & n43 ;
  assign n45 = n44 ^ n19 ;
  assign y0 = ~n45 ;
endmodule
