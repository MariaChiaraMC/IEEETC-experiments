module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 ;
  assign n9 = x3 ^ x1 ;
  assign n10 = x5 ^ x3 ;
  assign n11 = n10 ^ x5 ;
  assign n12 = x5 & ~x6 ;
  assign n13 = n12 ^ x5 ;
  assign n14 = n11 & ~n13 ;
  assign n15 = n14 ^ x5 ;
  assign n16 = n9 & ~n15 ;
  assign n17 = n16 ^ x1 ;
  assign n18 = x4 ^ x1 ;
  assign n19 = n18 ^ x1 ;
  assign n20 = n18 ^ n9 ;
  assign n21 = n20 ^ x6 ;
  assign n22 = n21 ^ x5 ;
  assign n23 = n22 ^ x1 ;
  assign n24 = n19 & n23 ;
  assign n25 = n24 ^ n22 ;
  assign n27 = n22 ^ x6 ;
  assign n26 = n21 ^ x7 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = n27 ^ n22 ;
  assign n30 = n29 ^ n21 ;
  assign n31 = ~n28 & n30 ;
  assign n32 = n31 ^ n22 ;
  assign n33 = n21 ^ n18 ;
  assign n34 = n33 ^ x1 ;
  assign n35 = n34 ^ n25 ;
  assign n36 = n32 & ~n35 ;
  assign n37 = n36 ^ n19 ;
  assign n38 = n25 & n37 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n39 ^ x4 ;
  assign n41 = n40 ^ n19 ;
  assign n42 = ~n17 & ~n41 ;
  assign n43 = x6 ^ x5 ;
  assign n44 = ~x3 & ~n43 ;
  assign n45 = ~x1 & ~x7 ;
  assign n46 = n45 ^ x4 ;
  assign n47 = x6 ^ x4 ;
  assign n48 = n47 ^ x4 ;
  assign n49 = n48 ^ n44 ;
  assign n50 = n46 & ~n49 ;
  assign n51 = n50 ^ n45 ;
  assign n52 = n44 & n51 ;
  assign n53 = n42 & ~n52 ;
  assign n54 = ~x2 & ~n53 ;
  assign n55 = x4 & ~x6 ;
  assign n56 = x2 & ~x3 ;
  assign n57 = x6 & ~n56 ;
  assign n58 = x5 & ~n57 ;
  assign n59 = ~n55 & n58 ;
  assign n60 = x2 & ~x4 ;
  assign n61 = x6 ^ x3 ;
  assign n62 = n61 ^ x3 ;
  assign n63 = n62 ^ n60 ;
  assign n64 = x7 ^ x5 ;
  assign n65 = x7 & n64 ;
  assign n66 = n65 ^ x3 ;
  assign n67 = n66 ^ x7 ;
  assign n68 = n63 & ~n67 ;
  assign n69 = n68 ^ n65 ;
  assign n70 = n69 ^ x7 ;
  assign n71 = n60 & n70 ;
  assign n72 = n71 ^ n60 ;
  assign n73 = ~n59 & ~n72 ;
  assign n74 = ~x1 & ~n73 ;
  assign n75 = ~n54 & ~n74 ;
  assign y0 = ~n75 ;
endmodule
