module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n15 = x5 ^ x1 ;
  assign n9 = x5 ^ x4 ;
  assign n10 = n9 ^ x6 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = n9 ^ x5 ;
  assign n13 = n12 ^ x1 ;
  assign n14 = ~n11 & ~n13 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n9 ^ x3 ;
  assign n18 = n17 ^ x1 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n10 ^ x2 ;
  assign n21 = n20 ^ x5 ;
  assign n22 = n17 & ~n21 ;
  assign n23 = n22 ^ n15 ;
  assign n24 = n19 & n23 ;
  assign n25 = n24 ^ n17 ;
  assign n26 = n16 & n25 ;
  assign n27 = n26 ^ n14 ;
  assign n28 = n27 ^ n15 ;
  assign n29 = x7 & n28 ;
  assign n30 = ~x0 & ~n29 ;
  assign y0 = ~n30 ;
endmodule
