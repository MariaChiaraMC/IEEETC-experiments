module top( x0 , x1 , x2 , x3 , x4 , y0 );
  input x0 , x1 , x2 , x3 , x4 ;
  output y0 ;
  wire n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 ;
  assign n6 = x2 ^ x0 ;
  assign n13 = x3 ^ x1 ;
  assign n14 = x4 ^ x3 ;
  assign n15 = n13 & ~n14 ;
  assign n16 = n15 ^ x1 ;
  assign n8 = ~x3 & ~x4 ;
  assign n7 = x3 & x4 ;
  assign n9 = n8 ^ n7 ;
  assign n10 = x1 & n9 ;
  assign n11 = n10 ^ n8 ;
  assign n12 = n11 ^ x2 ;
  assign n17 = n16 ^ n12 ;
  assign n18 = ~n6 & ~n17 ;
  assign n19 = n18 ^ n11 ;
  assign y0 = ~n19 ;
endmodule
