module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 ;
  assign n17 = x4 & ~x5 ;
  assign n18 = ~x1 & n17 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = n19 ^ x0 ;
  assign n37 = n20 ^ n19 ;
  assign n21 = ~x14 & x15 ;
  assign n22 = ~x12 & x13 ;
  assign n23 = ~n21 & ~n22 ;
  assign n24 = ~x10 & ~x11 ;
  assign n25 = ~x8 & x9 ;
  assign n26 = n24 & n25 ;
  assign n27 = x6 & x7 ;
  assign n28 = ~n26 & n27 ;
  assign n29 = n18 & ~n28 ;
  assign n30 = ~n23 & n29 ;
  assign n31 = n30 ^ n20 ;
  assign n32 = n31 ^ n19 ;
  assign n33 = n20 ^ n18 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = ~n32 & n35 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = n38 ^ n32 ;
  assign n40 = x5 ^ x4 ;
  assign n41 = n40 ^ x7 ;
  assign n43 = n41 ^ x5 ;
  assign n42 = n41 ^ x7 ;
  assign n44 = n43 ^ n42 ;
  assign n52 = n44 ^ n41 ;
  assign n53 = n52 ^ n43 ;
  assign n54 = n53 ^ n43 ;
  assign n64 = x11 ^ x10 ;
  assign n55 = x10 ^ x6 ;
  assign n56 = n55 ^ x11 ;
  assign n57 = n56 ^ x11 ;
  assign n58 = n57 ^ x10 ;
  assign n59 = n56 ^ x9 ;
  assign n60 = n59 ^ x8 ;
  assign n61 = n60 ^ n56 ;
  assign n62 = n61 ^ n58 ;
  assign n63 = ~n58 & n62 ;
  assign n65 = n64 ^ n63 ;
  assign n66 = n65 ^ n58 ;
  assign n67 = x10 ^ x8 ;
  assign n68 = n63 ^ n58 ;
  assign n69 = n67 & ~n68 ;
  assign n70 = n69 ^ x10 ;
  assign n71 = n66 & ~n70 ;
  assign n72 = n71 ^ x10 ;
  assign n73 = n72 ^ x10 ;
  assign n74 = n73 ^ n41 ;
  assign n75 = n74 ^ n41 ;
  assign n76 = n75 ^ n43 ;
  assign n77 = ~n54 & ~n76 ;
  assign n45 = x8 & ~x9 ;
  assign n46 = x6 & n45 ;
  assign n47 = n24 & n46 ;
  assign n48 = n47 ^ n41 ;
  assign n49 = n48 ^ n44 ;
  assign n50 = n49 ^ n43 ;
  assign n51 = n44 & n50 ;
  assign n78 = n77 ^ n51 ;
  assign n79 = n78 ^ n44 ;
  assign n80 = n51 ^ n43 ;
  assign n81 = n80 ^ n53 ;
  assign n82 = ~n43 & ~n81 ;
  assign n83 = n82 ^ n51 ;
  assign n84 = n79 & n83 ;
  assign n85 = n84 ^ n77 ;
  assign n86 = n85 ^ n82 ;
  assign n87 = n86 ^ n44 ;
  assign n88 = n87 ^ n43 ;
  assign n89 = n88 ^ n53 ;
  assign n90 = n89 ^ x5 ;
  assign n91 = ~n23 & ~n90 ;
  assign n92 = x13 ^ x12 ;
  assign n93 = n21 ^ x13 ;
  assign n94 = n93 ^ n21 ;
  assign n95 = x14 & ~x15 ;
  assign n96 = n95 ^ n21 ;
  assign n97 = n94 & n96 ;
  assign n98 = n97 ^ n21 ;
  assign n99 = n92 & n98 ;
  assign n100 = ~x11 & n99 ;
  assign n101 = ~x10 & x13 ;
  assign n102 = x14 ^ x12 ;
  assign n103 = n101 & n102 ;
  assign n104 = x15 & n103 ;
  assign n105 = ~n100 & ~n104 ;
  assign n106 = x5 & ~x7 ;
  assign n107 = ~n24 & n106 ;
  assign n108 = x6 & n107 ;
  assign n109 = ~n105 & n108 ;
  assign n110 = ~x5 & x7 ;
  assign n111 = n46 & n110 ;
  assign n112 = ~x4 & n111 ;
  assign n113 = ~n109 & ~n112 ;
  assign n114 = ~n91 & n113 ;
  assign n115 = ~x1 & ~n114 ;
  assign n116 = x1 & x7 ;
  assign n117 = x9 & x10 ;
  assign n118 = x1 & ~x13 ;
  assign n119 = ~n117 & n118 ;
  assign n120 = x8 & ~n119 ;
  assign n121 = ~x8 & ~x13 ;
  assign n122 = ~x14 & ~x15 ;
  assign n123 = ~n121 & ~n122 ;
  assign n124 = ~x12 & ~n123 ;
  assign n125 = ~x9 & n24 ;
  assign n126 = n125 ^ x11 ;
  assign n127 = n124 & ~n126 ;
  assign n128 = ~n120 & n127 ;
  assign n129 = ~x1 & ~x13 ;
  assign n130 = ~x14 & n121 ;
  assign n131 = ~n129 & ~n130 ;
  assign n132 = n131 ^ x14 ;
  assign n133 = ~x15 & ~n132 ;
  assign n134 = n133 ^ x14 ;
  assign n135 = n128 & ~n134 ;
  assign n136 = ~n116 & ~n135 ;
  assign n137 = n17 & ~n136 ;
  assign n138 = ~x6 & n137 ;
  assign n139 = ~n115 & ~n138 ;
  assign n140 = n139 ^ n19 ;
  assign n141 = n36 ^ n32 ;
  assign n142 = ~n140 & ~n141 ;
  assign n143 = n142 ^ n19 ;
  assign n144 = ~n39 & ~n143 ;
  assign n145 = n144 ^ n19 ;
  assign n146 = n145 ^ x2 ;
  assign n147 = n146 ^ n19 ;
  assign n148 = ~x3 & ~n147 ;
  assign y0 = n148 ;
endmodule
