module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 ;
  assign n36 = x7 & x10 ;
  assign n37 = x3 & x4 ;
  assign n38 = n36 & n37 ;
  assign n16 = x5 & x7 ;
  assign n17 = ~x14 & n16 ;
  assign n18 = ~x0 & ~x2 ;
  assign n19 = ~x3 & ~x6 ;
  assign n20 = n18 & n19 ;
  assign n21 = n17 & n20 ;
  assign n22 = x3 & x14 ;
  assign n23 = x0 & x6 ;
  assign n24 = n22 & n23 ;
  assign n25 = x9 ^ x7 ;
  assign n26 = n24 & n25 ;
  assign n27 = ~x5 & n26 ;
  assign n28 = ~n21 & ~n27 ;
  assign n29 = ~x4 & ~x10 ;
  assign n30 = ~n28 & n29 ;
  assign n39 = n38 ^ n30 ;
  assign n40 = n39 ^ n30 ;
  assign n31 = x6 & ~x14 ;
  assign n32 = ~x9 & n31 ;
  assign n33 = n18 & n32 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ n30 ;
  assign n41 = n40 ^ n35 ;
  assign n42 = n30 ^ x5 ;
  assign n43 = n42 ^ n30 ;
  assign n44 = n43 ^ n40 ;
  assign n45 = n40 & ~n44 ;
  assign n46 = n45 ^ n40 ;
  assign n47 = n41 & n46 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = n48 ^ n30 ;
  assign n50 = n49 ^ n40 ;
  assign n51 = x1 & n50 ;
  assign n52 = n51 ^ n30 ;
  assign n53 = x8 & n52 ;
  assign n54 = ~x12 & n53 ;
  assign n55 = ~x0 & ~x8 ;
  assign n56 = ~x1 & x2 ;
  assign n57 = ~x4 & ~x5 ;
  assign n58 = ~x6 & n57 ;
  assign n59 = n22 & n36 ;
  assign n60 = n58 & n59 ;
  assign n61 = ~x7 & ~x10 ;
  assign n62 = ~x3 & n61 ;
  assign n63 = x4 & x5 ;
  assign n64 = n62 & n63 ;
  assign n65 = n32 & n64 ;
  assign n66 = ~n60 & ~n65 ;
  assign n67 = n56 & ~n66 ;
  assign n68 = n31 & n38 ;
  assign n69 = n19 & n61 ;
  assign n70 = ~x4 & n69 ;
  assign n71 = ~n68 & ~n70 ;
  assign n72 = ~x2 & ~x5 ;
  assign n73 = ~x1 & ~x9 ;
  assign n74 = n72 & n73 ;
  assign n75 = ~n71 & n74 ;
  assign n76 = ~n67 & ~n75 ;
  assign n77 = ~x12 & ~n76 ;
  assign n78 = x1 & ~x12 ;
  assign n79 = x9 & n37 ;
  assign n80 = n78 & n79 ;
  assign n81 = ~x14 & n80 ;
  assign n82 = x10 ^ x7 ;
  assign n83 = x6 & n82 ;
  assign n84 = n83 ^ x2 ;
  assign n85 = x5 ^ x2 ;
  assign n86 = n82 ^ x10 ;
  assign n87 = n86 ^ n85 ;
  assign n88 = ~n85 & ~n87 ;
  assign n89 = n88 ^ x2 ;
  assign n90 = n89 ^ n85 ;
  assign n91 = n84 & ~n90 ;
  assign n92 = n91 ^ x2 ;
  assign n93 = n92 ^ x2 ;
  assign n94 = n81 & n93 ;
  assign n95 = x9 & x10 ;
  assign n96 = ~x14 & n95 ;
  assign n97 = n19 & n63 ;
  assign n98 = n96 & n97 ;
  assign n99 = n56 & n98 ;
  assign n100 = ~n94 & ~n99 ;
  assign n101 = ~n77 & n100 ;
  assign n102 = n55 & ~n101 ;
  assign n103 = x7 & ~x9 ;
  assign n104 = x14 & n103 ;
  assign n105 = ~x3 & n56 ;
  assign n106 = n104 & ~n105 ;
  assign n107 = ~x2 & x3 ;
  assign n108 = n57 & ~n107 ;
  assign n109 = ~x8 & ~x10 ;
  assign n110 = ~n78 & n109 ;
  assign n111 = n108 & n110 ;
  assign n112 = n23 & n111 ;
  assign n113 = n106 & n112 ;
  assign n114 = ~n102 & ~n113 ;
  assign n115 = ~n54 & n114 ;
  assign n116 = ~x13 & ~n115 ;
  assign n117 = ~x12 & n55 ;
  assign n118 = x14 & n56 ;
  assign n119 = n97 & n118 ;
  assign n120 = n117 & n119 ;
  assign n121 = n95 & n120 ;
  assign n122 = ~n116 & ~n121 ;
  assign n123 = ~x11 & ~n122 ;
  assign y0 = n123 ;
endmodule
