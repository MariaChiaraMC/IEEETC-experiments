module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 ;
  assign n10 = x4 & x7 ;
  assign n11 = ~x0 & n10 ;
  assign n12 = x6 ^ x3 ;
  assign n13 = n12 ^ x6 ;
  assign n14 = x6 ^ x2 ;
  assign n15 = ~n13 & n14 ;
  assign n16 = n15 ^ x6 ;
  assign n17 = x1 & ~x6 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = ~n16 & n18 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = x5 & n20 ;
  assign n22 = n21 ^ x5 ;
  assign n23 = n11 & n22 ;
  assign y0 = n23 ;
endmodule
