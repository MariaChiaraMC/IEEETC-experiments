module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 ;
  assign n25 = ~x6 & ~x7 ;
  assign n26 = ~x9 & n25 ;
  assign n27 = ~x8 & ~x22 ;
  assign n28 = n26 & n27 ;
  assign n29 = ~x1 & ~x2 ;
  assign n30 = ~x12 & n29 ;
  assign n31 = n30 ^ x0 ;
  assign n32 = x15 & x17 ;
  assign n33 = x16 & n32 ;
  assign n34 = ~x13 & n33 ;
  assign n35 = x13 & ~x15 ;
  assign n36 = ~x16 & ~x17 ;
  assign n37 = n35 & n36 ;
  assign n38 = ~n34 & ~n37 ;
  assign n39 = ~x10 & x11 ;
  assign n40 = x14 & n39 ;
  assign n41 = x5 ^ x3 ;
  assign n42 = ~x4 & n41 ;
  assign n43 = ~x3 & ~x5 ;
  assign n44 = x0 & n43 ;
  assign n45 = ~n42 & ~n44 ;
  assign n46 = n40 & ~n45 ;
  assign n47 = ~n38 & n46 ;
  assign n48 = ~x16 & n35 ;
  assign n49 = ~x14 & x17 ;
  assign n50 = n39 & n49 ;
  assign n51 = n48 & n50 ;
  assign n52 = ~x14 & ~x17 ;
  assign n53 = ~x11 & ~x13 ;
  assign n54 = ~x16 & n53 ;
  assign n55 = n52 & n54 ;
  assign n56 = x10 & x15 ;
  assign n57 = n55 & n56 ;
  assign n58 = ~n51 & ~n57 ;
  assign n59 = ~x4 & n44 ;
  assign n60 = ~n58 & n59 ;
  assign n61 = ~n47 & ~n60 ;
  assign n62 = n61 ^ n31 ;
  assign n63 = n62 ^ n30 ;
  assign n64 = n63 ^ n62 ;
  assign n125 = x23 & n43 ;
  assign n126 = ~x4 & n125 ;
  assign n127 = n29 & n126 ;
  assign n128 = x10 & n127 ;
  assign n65 = x14 & x17 ;
  assign n66 = x1 & ~n52 ;
  assign n67 = ~n65 & n66 ;
  assign n68 = ~x2 & ~x3 ;
  assign n69 = n68 ^ x4 ;
  assign n70 = x17 ^ x5 ;
  assign n71 = n70 ^ x17 ;
  assign n72 = x17 ^ x1 ;
  assign n73 = ~n71 & n72 ;
  assign n74 = n73 ^ x17 ;
  assign n75 = n74 ^ n68 ;
  assign n76 = ~n69 & n75 ;
  assign n77 = n76 ^ n73 ;
  assign n78 = n77 ^ x17 ;
  assign n79 = n78 ^ x4 ;
  assign n80 = n68 & ~n79 ;
  assign n81 = n80 ^ n68 ;
  assign n82 = ~n67 & ~n81 ;
  assign n83 = n48 & ~n82 ;
  assign n84 = ~x4 & ~x5 ;
  assign n85 = ~x23 & n84 ;
  assign n86 = n29 & n85 ;
  assign n87 = n86 ^ x1 ;
  assign n88 = x14 & n34 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = n89 ^ n86 ;
  assign n91 = n90 ^ n89 ;
  assign n92 = ~x15 & ~x16 ;
  assign n95 = n84 ^ x13 ;
  assign n96 = n95 ^ x13 ;
  assign n93 = x13 ^ x2 ;
  assign n94 = n93 ^ x13 ;
  assign n97 = n96 ^ n94 ;
  assign n98 = x14 & x23 ;
  assign n99 = n98 ^ x13 ;
  assign n100 = n99 ^ x13 ;
  assign n101 = n100 ^ n96 ;
  assign n102 = n96 & n101 ;
  assign n103 = n102 ^ n96 ;
  assign n104 = ~n97 & n103 ;
  assign n105 = n104 ^ n102 ;
  assign n106 = n105 ^ x13 ;
  assign n107 = n106 ^ n96 ;
  assign n108 = ~x3 & n107 ;
  assign n109 = n108 ^ x13 ;
  assign n110 = n92 & n109 ;
  assign n111 = n110 ^ n89 ;
  assign n112 = n111 ^ n87 ;
  assign n113 = ~n91 & ~n112 ;
  assign n114 = n113 ^ n110 ;
  assign n115 = ~n48 & ~n110 ;
  assign n116 = n115 ^ n87 ;
  assign n117 = ~n114 & ~n116 ;
  assign n118 = n117 ^ n115 ;
  assign n119 = ~n87 & n118 ;
  assign n120 = n119 ^ n113 ;
  assign n121 = n120 ^ x1 ;
  assign n122 = n121 ^ n110 ;
  assign n123 = ~n83 & ~n122 ;
  assign n124 = n39 & ~n123 ;
  assign n129 = n128 ^ n124 ;
  assign n130 = n129 ^ x12 ;
  assign n151 = n130 ^ n129 ;
  assign n131 = x17 ^ x16 ;
  assign n132 = n131 ^ x14 ;
  assign n133 = n132 ^ x15 ;
  assign n134 = n133 ^ n53 ;
  assign n135 = x17 ^ x15 ;
  assign n136 = x15 ^ x14 ;
  assign n137 = n136 ^ n135 ;
  assign n138 = ~n135 & n137 ;
  assign n139 = n138 ^ x15 ;
  assign n140 = n139 ^ n135 ;
  assign n141 = ~n134 & ~n140 ;
  assign n142 = n141 ^ n138 ;
  assign n143 = n142 ^ n135 ;
  assign n144 = n53 & ~n143 ;
  assign n145 = n144 ^ n130 ;
  assign n146 = n145 ^ n129 ;
  assign n147 = n130 ^ n124 ;
  assign n148 = n147 ^ n144 ;
  assign n149 = n148 ^ n146 ;
  assign n150 = n146 & ~n149 ;
  assign n152 = n151 ^ n150 ;
  assign n153 = n152 ^ n146 ;
  assign n154 = ~x14 & n33 ;
  assign n155 = ~x15 & n36 ;
  assign n156 = ~n154 & ~n155 ;
  assign n157 = n156 ^ x13 ;
  assign n158 = n157 ^ n156 ;
  assign n159 = n158 ^ x11 ;
  assign n160 = n52 ^ x15 ;
  assign n161 = ~n52 & n160 ;
  assign n162 = n161 ^ n156 ;
  assign n163 = n162 ^ n52 ;
  assign n164 = n159 & n163 ;
  assign n165 = n164 ^ n161 ;
  assign n166 = n165 ^ n52 ;
  assign n167 = x11 & ~n166 ;
  assign n168 = n167 ^ x11 ;
  assign n169 = n168 ^ n129 ;
  assign n170 = n150 ^ n146 ;
  assign n171 = n169 & n170 ;
  assign n172 = n171 ^ n129 ;
  assign n173 = ~n153 & n172 ;
  assign n174 = n173 ^ n129 ;
  assign n175 = n174 ^ n128 ;
  assign n176 = n175 ^ n129 ;
  assign n177 = n176 ^ n62 ;
  assign n178 = n177 ^ n31 ;
  assign n179 = n64 & n178 ;
  assign n180 = n179 ^ n176 ;
  assign n181 = x21 ^ x20 ;
  assign n182 = n181 ^ x21 ;
  assign n183 = x18 & x19 ;
  assign n184 = n183 ^ x21 ;
  assign n185 = n182 & ~n184 ;
  assign n186 = n185 ^ x21 ;
  assign n187 = x10 & ~n186 ;
  assign n188 = ~x13 & ~n187 ;
  assign n189 = x11 & n126 ;
  assign n190 = ~n188 & n189 ;
  assign n191 = n190 ^ x10 ;
  assign n192 = n190 ^ n154 ;
  assign n193 = n192 ^ n154 ;
  assign n194 = ~x4 & ~x14 ;
  assign n196 = x15 & ~x17 ;
  assign n195 = x13 & n125 ;
  assign n197 = n196 ^ n195 ;
  assign n198 = n41 & n54 ;
  assign n199 = n198 ^ n195 ;
  assign n200 = n199 ^ n198 ;
  assign n201 = ~x16 & x17 ;
  assign n202 = n201 ^ n198 ;
  assign n203 = n200 & ~n202 ;
  assign n204 = n203 ^ n198 ;
  assign n205 = n197 & ~n204 ;
  assign n206 = n205 ^ n196 ;
  assign n207 = n194 & n206 ;
  assign n208 = n207 ^ n154 ;
  assign n209 = ~n193 & ~n208 ;
  assign n210 = n209 ^ n154 ;
  assign n211 = n191 & n210 ;
  assign n212 = n211 ^ x10 ;
  assign n213 = ~n176 & ~n212 ;
  assign n214 = n213 ^ n31 ;
  assign n215 = ~n180 & n214 ;
  assign n216 = n215 ^ n213 ;
  assign n217 = n31 & n216 ;
  assign n218 = n217 ^ n179 ;
  assign n219 = n218 ^ x0 ;
  assign n220 = n219 ^ n176 ;
  assign n221 = n28 & n220 ;
  assign y0 = n221 ;
endmodule
