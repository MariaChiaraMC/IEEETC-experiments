module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 ;
  output y0 ;
  wire n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 ;
  assign n23 = x0 & ~x1 ;
  assign n24 = x3 & n23 ;
  assign n25 = ~x0 & ~x2 ;
  assign n26 = x1 & n25 ;
  assign n27 = ~n24 & ~n26 ;
  assign n28 = ~x3 & x5 ;
  assign n29 = x3 & ~x5 ;
  assign n30 = ~n28 & ~n29 ;
  assign n31 = ~n27 & n30 ;
  assign n32 = ~x4 & n31 ;
  assign n234 = ~x19 & ~x20 ;
  assign n44 = x11 ^ x10 ;
  assign n45 = x13 ^ x11 ;
  assign n46 = n45 ^ x11 ;
  assign n47 = n46 ^ n44 ;
  assign n48 = ~x6 & ~x7 ;
  assign n49 = n48 ^ x12 ;
  assign n50 = ~x12 & ~n49 ;
  assign n51 = n50 ^ x11 ;
  assign n52 = n51 ^ x12 ;
  assign n53 = ~n47 & ~n52 ;
  assign n54 = n53 ^ n50 ;
  assign n55 = n54 ^ x12 ;
  assign n56 = n44 & ~n55 ;
  assign n57 = ~x9 & n56 ;
  assign n58 = ~x12 & ~x13 ;
  assign n59 = x9 & n58 ;
  assign n60 = n48 & n59 ;
  assign n61 = ~x0 & n60 ;
  assign n62 = ~x10 & ~x11 ;
  assign n63 = n61 & n62 ;
  assign n64 = ~n57 & ~n63 ;
  assign n65 = ~x8 & ~n64 ;
  assign n34 = ~x1 & x2 ;
  assign n35 = x0 & ~n34 ;
  assign n66 = n65 ^ n35 ;
  assign n36 = n35 ^ x3 ;
  assign n41 = n36 ^ n35 ;
  assign n67 = n41 ^ x5 ;
  assign n68 = n66 & n67 ;
  assign n33 = x1 & x2 ;
  assign n37 = n36 ^ x4 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = n38 ^ n33 ;
  assign n40 = ~n33 & ~n39 ;
  assign n74 = n68 ^ n40 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = n42 ^ n33 ;
  assign n69 = n35 ^ n33 ;
  assign n70 = n69 ^ n68 ;
  assign n71 = n70 ^ n66 ;
  assign n72 = n71 ^ x5 ;
  assign n73 = ~n43 & n72 ;
  assign n75 = n74 ^ n73 ;
  assign n76 = n75 ^ n69 ;
  assign n77 = n76 ^ n66 ;
  assign n78 = n77 ^ n41 ;
  assign n79 = x5 & n78 ;
  assign n151 = x3 ^ x1 ;
  assign n80 = x11 & x13 ;
  assign n81 = x7 & n80 ;
  assign n82 = ~x12 & n81 ;
  assign n83 = ~x8 & x9 ;
  assign n84 = x11 & ~x12 ;
  assign n85 = x13 & n62 ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = n83 & ~n86 ;
  assign n88 = x11 & ~x16 ;
  assign n89 = ~x9 & x10 ;
  assign n90 = x9 & x11 ;
  assign n91 = ~n89 & ~n90 ;
  assign n92 = ~n88 & n91 ;
  assign n93 = ~x6 & n92 ;
  assign n94 = x13 & ~n93 ;
  assign n95 = ~x12 & ~n90 ;
  assign n96 = x6 & ~n95 ;
  assign n97 = x10 & x11 ;
  assign n98 = x8 & n97 ;
  assign n99 = ~n96 & ~n98 ;
  assign n100 = x7 & ~n99 ;
  assign n101 = ~x8 & ~x15 ;
  assign n102 = x9 & x10 ;
  assign n103 = ~x12 & n102 ;
  assign n104 = ~x13 & ~n103 ;
  assign n105 = ~n101 & ~n104 ;
  assign n106 = ~x9 & ~x10 ;
  assign n107 = ~x13 & ~n106 ;
  assign n108 = ~x8 & ~n88 ;
  assign n109 = ~n107 & n108 ;
  assign n110 = n48 & ~n109 ;
  assign n111 = x12 & ~n80 ;
  assign n112 = ~x6 & n111 ;
  assign n113 = ~x17 & ~n112 ;
  assign n114 = ~n110 & n113 ;
  assign n115 = ~n105 & n114 ;
  assign n116 = ~n100 & n115 ;
  assign n117 = ~n94 & n116 ;
  assign n118 = x2 & ~n117 ;
  assign n119 = ~n87 & ~n118 ;
  assign n120 = ~n82 & n119 ;
  assign n121 = n120 ^ x2 ;
  assign n122 = n121 ^ x1 ;
  assign n130 = n122 ^ n121 ;
  assign n123 = n84 & n102 ;
  assign n124 = n123 ^ n122 ;
  assign n125 = n124 ^ n121 ;
  assign n126 = n122 ^ n120 ;
  assign n127 = n126 ^ n123 ;
  assign n128 = n127 ^ n125 ;
  assign n129 = n125 & n128 ;
  assign n131 = n130 ^ n129 ;
  assign n132 = n131 ^ n125 ;
  assign n133 = n121 ^ x13 ;
  assign n134 = n129 ^ n125 ;
  assign n135 = ~n133 & n134 ;
  assign n136 = n135 ^ n121 ;
  assign n137 = ~n132 & n136 ;
  assign n138 = n137 ^ n121 ;
  assign n139 = n138 ^ x2 ;
  assign n140 = n139 ^ n121 ;
  assign n141 = x4 & ~n140 ;
  assign n142 = x4 ^ x2 ;
  assign n143 = n142 ^ x4 ;
  assign n144 = x1 & x4 ;
  assign n145 = n144 ^ x4 ;
  assign n146 = ~n143 & ~n145 ;
  assign n147 = n146 ^ x4 ;
  assign n148 = ~x0 & ~n147 ;
  assign n149 = ~n141 & ~n148 ;
  assign n150 = n149 ^ x3 ;
  assign n152 = n151 ^ n150 ;
  assign n153 = n152 ^ x2 ;
  assign n154 = n153 ^ n152 ;
  assign n155 = n152 ^ n150 ;
  assign n156 = n155 ^ x3 ;
  assign n157 = ~n154 & ~n156 ;
  assign n158 = n157 ^ n150 ;
  assign n159 = ~x12 & x13 ;
  assign n160 = n150 & n159 ;
  assign n161 = n160 ^ x3 ;
  assign n162 = n158 & ~n161 ;
  assign n163 = n162 ^ n160 ;
  assign n164 = ~x3 & n163 ;
  assign n165 = n164 ^ n157 ;
  assign n166 = n165 ^ n149 ;
  assign n167 = n166 ^ n150 ;
  assign n168 = n79 & n167 ;
  assign n169 = ~x10 & x11 ;
  assign n170 = n59 & n169 ;
  assign n171 = x8 & n48 ;
  assign n172 = n170 & n171 ;
  assign n173 = n24 & n172 ;
  assign n174 = ~x5 & ~n173 ;
  assign n175 = ~x11 & n58 ;
  assign n176 = ~x4 & n175 ;
  assign n177 = n48 & n176 ;
  assign n178 = n25 & n177 ;
  assign n179 = n83 & n178 ;
  assign n180 = ~x3 & ~x8 ;
  assign n181 = ~x11 & n180 ;
  assign n182 = ~x2 & x8 ;
  assign n183 = n169 & n182 ;
  assign n184 = ~n181 & ~n183 ;
  assign n185 = x1 & n61 ;
  assign n186 = ~n184 & n185 ;
  assign n187 = ~n144 & ~n186 ;
  assign n188 = n187 ^ x4 ;
  assign n189 = n188 ^ n187 ;
  assign n190 = n187 ^ n23 ;
  assign n191 = n189 & ~n190 ;
  assign n192 = n191 ^ n187 ;
  assign n193 = x2 & x21 ;
  assign n194 = x3 & ~n193 ;
  assign n195 = ~n187 & n194 ;
  assign n196 = n195 ^ n179 ;
  assign n197 = ~n192 & ~n196 ;
  assign n198 = n197 ^ n195 ;
  assign n199 = ~n179 & n198 ;
  assign n200 = n199 ^ n179 ;
  assign n201 = n174 & ~n200 ;
  assign n202 = ~n168 & ~n201 ;
  assign n203 = x10 & n175 ;
  assign n204 = n48 & n203 ;
  assign n205 = ~x8 & n204 ;
  assign n206 = x3 & ~n205 ;
  assign n207 = n25 ^ x4 ;
  assign n208 = n207 ^ n25 ;
  assign n209 = x0 & ~x3 ;
  assign n210 = n209 ^ n25 ;
  assign n211 = n208 & n210 ;
  assign n212 = n211 ^ n25 ;
  assign n213 = ~x1 & n212 ;
  assign n214 = ~n206 & n213 ;
  assign n215 = ~x0 & n144 ;
  assign n216 = ~x5 & n215 ;
  assign n217 = ~x5 & n23 ;
  assign n218 = n151 & ~n217 ;
  assign n219 = ~x4 & n218 ;
  assign n220 = n219 ^ n217 ;
  assign n221 = n172 & n220 ;
  assign n222 = ~x9 & n169 ;
  assign n223 = ~n204 & ~n222 ;
  assign n224 = n217 & ~n223 ;
  assign n225 = n89 & n177 ;
  assign n226 = x1 & n225 ;
  assign n227 = ~n224 & ~n226 ;
  assign n228 = n180 & ~n227 ;
  assign n229 = ~n221 & ~n228 ;
  assign n230 = ~n216 & n229 ;
  assign n231 = x2 & ~n230 ;
  assign n232 = ~n214 & ~n231 ;
  assign n233 = ~n202 & n232 ;
  assign n235 = n234 ^ n233 ;
  assign n236 = n235 ^ n233 ;
  assign n237 = n233 ^ x18 ;
  assign n238 = ~n236 & n237 ;
  assign n239 = n238 ^ n233 ;
  assign n240 = ~n32 & n239 ;
  assign n241 = x14 & ~n240 ;
  assign y0 = n241 ;
endmodule
