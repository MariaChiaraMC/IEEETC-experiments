module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 ;
  assign n11 = x5 & ~x8 ;
  assign n12 = x0 & x2 ;
  assign n13 = x7 & n12 ;
  assign n14 = x6 & x9 ;
  assign n15 = ~x3 & ~x4 ;
  assign n16 = n14 & n15 ;
  assign n17 = n13 & n16 ;
  assign n18 = n11 & n17 ;
  assign n19 = ~x3 & ~x7 ;
  assign n20 = x4 & x5 ;
  assign n21 = n12 & n20 ;
  assign n22 = x5 & x8 ;
  assign n23 = x0 & ~x2 ;
  assign n24 = n22 & n23 ;
  assign n25 = ~n21 & ~n24 ;
  assign n26 = n19 & ~n25 ;
  assign n27 = ~x2 & ~x7 ;
  assign n46 = ~n20 & ~n27 ;
  assign n28 = n22 & n27 ;
  assign n29 = ~x4 & ~x5 ;
  assign n32 = ~x2 & ~x8 ;
  assign n30 = x4 & ~x8 ;
  assign n31 = x2 & ~n30 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = n33 ^ n32 ;
  assign n35 = n32 ^ n22 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n34 & ~n36 ;
  assign n38 = n37 ^ n32 ;
  assign n39 = ~n29 & n38 ;
  assign n40 = n39 ^ n32 ;
  assign n41 = x7 & n40 ;
  assign n42 = ~n28 & ~n41 ;
  assign n47 = n46 ^ n42 ;
  assign n48 = n47 ^ n42 ;
  assign n43 = x5 & ~x7 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = n44 ^ n42 ;
  assign n49 = n48 ^ n45 ;
  assign n50 = n42 ^ x8 ;
  assign n51 = n50 ^ n42 ;
  assign n52 = n51 ^ n48 ;
  assign n53 = ~n48 & n52 ;
  assign n54 = n53 ^ n48 ;
  assign n55 = n49 & ~n54 ;
  assign n56 = n55 ^ n53 ;
  assign n57 = n56 ^ n42 ;
  assign n58 = n57 ^ n48 ;
  assign n59 = ~x3 & n58 ;
  assign n60 = n59 ^ n42 ;
  assign n61 = ~x0 & ~n60 ;
  assign n62 = ~x5 & n12 ;
  assign n63 = x7 & ~x8 ;
  assign n64 = n62 & n63 ;
  assign n65 = ~n28 & ~n64 ;
  assign n66 = n65 ^ x4 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = n67 ^ x3 ;
  assign n69 = ~x5 & x7 ;
  assign n70 = n69 ^ n23 ;
  assign n71 = n23 & n70 ;
  assign n72 = n71 ^ n65 ;
  assign n73 = n72 ^ n23 ;
  assign n74 = n68 & ~n73 ;
  assign n75 = n74 ^ n71 ;
  assign n76 = n75 ^ n23 ;
  assign n77 = x3 & n76 ;
  assign n78 = ~n61 & ~n77 ;
  assign n79 = ~n26 & n78 ;
  assign n80 = n14 & ~n79 ;
  assign n81 = ~x0 & x2 ;
  assign n82 = x8 & n81 ;
  assign n83 = x5 ^ x4 ;
  assign n84 = x7 & ~n83 ;
  assign n85 = n84 ^ x4 ;
  assign n86 = n85 ^ n84 ;
  assign n87 = n84 ^ n43 ;
  assign n88 = n87 ^ n84 ;
  assign n89 = ~n86 & n88 ;
  assign n90 = n89 ^ n84 ;
  assign n91 = x9 & n90 ;
  assign n92 = n91 ^ n84 ;
  assign n93 = n82 & n92 ;
  assign n94 = ~x4 & ~x9 ;
  assign n95 = x0 & ~x8 ;
  assign n96 = ~x5 & n27 ;
  assign n97 = n95 & n96 ;
  assign n98 = n94 & n97 ;
  assign n99 = ~n93 & ~n98 ;
  assign n100 = x3 & ~n99 ;
  assign n101 = ~x6 & x9 ;
  assign n102 = x7 & n95 ;
  assign n103 = ~x3 & x4 ;
  assign n104 = n102 & n103 ;
  assign n105 = x7 & x8 ;
  assign n106 = ~n19 & ~n105 ;
  assign n107 = ~x4 & ~n106 ;
  assign n108 = ~x0 & n107 ;
  assign n109 = ~n104 & ~n108 ;
  assign n110 = x2 & ~n109 ;
  assign n111 = ~x5 & n110 ;
  assign n112 = ~x3 & ~x8 ;
  assign n113 = x0 & x8 ;
  assign n114 = ~n112 & ~n113 ;
  assign n115 = ~n15 & n96 ;
  assign n116 = ~n114 & n115 ;
  assign n117 = ~x2 & n19 ;
  assign n118 = n95 & n117 ;
  assign n119 = x3 & x4 ;
  assign n120 = x2 ^ x0 ;
  assign n121 = n120 ^ x7 ;
  assign n122 = n121 ^ x8 ;
  assign n123 = n122 ^ x7 ;
  assign n124 = n123 ^ x8 ;
  assign n125 = x8 & n124 ;
  assign n126 = n125 ^ n122 ;
  assign n127 = n126 ^ x8 ;
  assign n128 = n122 ^ x2 ;
  assign n129 = x5 & ~n128 ;
  assign n130 = n129 ^ n122 ;
  assign n131 = ~n127 & ~n130 ;
  assign n132 = n131 ^ n122 ;
  assign n133 = n119 & ~n132 ;
  assign n134 = ~n118 & ~n133 ;
  assign n135 = ~n116 & n134 ;
  assign n136 = ~n111 & n135 ;
  assign n137 = n101 & ~n136 ;
  assign n138 = ~n100 & ~n137 ;
  assign n139 = ~n80 & n138 ;
  assign n140 = x5 & n105 ;
  assign n141 = ~x2 & x3 ;
  assign n142 = n140 & n141 ;
  assign n143 = n142 ^ x8 ;
  assign n144 = n143 ^ x0 ;
  assign n155 = n144 ^ n143 ;
  assign n145 = x3 & x5 ;
  assign n146 = ~x3 & ~x5 ;
  assign n147 = ~n145 & ~n146 ;
  assign n148 = n27 & ~n147 ;
  assign n149 = n148 ^ n144 ;
  assign n150 = n149 ^ n143 ;
  assign n151 = n144 ^ n142 ;
  assign n152 = n151 ^ n148 ;
  assign n153 = n152 ^ n150 ;
  assign n154 = ~n150 & n153 ;
  assign n156 = n155 ^ n154 ;
  assign n157 = n156 ^ n150 ;
  assign n158 = x3 ^ x2 ;
  assign n159 = n69 ^ x3 ;
  assign n160 = n159 ^ n69 ;
  assign n161 = n69 ^ n43 ;
  assign n162 = ~n160 & n161 ;
  assign n163 = n162 ^ n69 ;
  assign n164 = n158 & n163 ;
  assign n165 = n164 ^ n143 ;
  assign n166 = n154 ^ n150 ;
  assign n167 = n165 & ~n166 ;
  assign n168 = n167 ^ n143 ;
  assign n169 = ~n157 & ~n168 ;
  assign n170 = n169 ^ n143 ;
  assign n171 = n170 ^ x8 ;
  assign n172 = n171 ^ n143 ;
  assign n173 = n94 & ~n172 ;
  assign n174 = n173 ^ x9 ;
  assign n175 = n174 ^ n173 ;
  assign n176 = ~x3 & x5 ;
  assign n177 = n102 & n176 ;
  assign n178 = ~x3 & n105 ;
  assign n179 = ~x7 & ~x8 ;
  assign n180 = ~n178 & ~n179 ;
  assign n181 = n62 & ~n180 ;
  assign n182 = x2 & x3 ;
  assign n183 = n140 & n182 ;
  assign n184 = ~n181 & ~n183 ;
  assign n185 = ~n177 & n184 ;
  assign n186 = x4 & ~n185 ;
  assign n187 = x8 & n29 ;
  assign n188 = ~n22 & ~n29 ;
  assign n189 = ~x0 & n182 ;
  assign n190 = ~n188 & n189 ;
  assign n191 = ~n187 & ~n190 ;
  assign n192 = ~x0 & ~x2 ;
  assign n193 = ~x3 & ~n192 ;
  assign n194 = x7 & ~n141 ;
  assign n195 = ~n193 & n194 ;
  assign n196 = ~n191 & n195 ;
  assign n197 = ~n186 & ~n196 ;
  assign n198 = n197 ^ n173 ;
  assign n199 = n198 ^ n173 ;
  assign n200 = ~n175 & ~n199 ;
  assign n201 = n200 ^ n173 ;
  assign n202 = x6 & n201 ;
  assign n203 = n202 ^ n173 ;
  assign n204 = n139 & ~n203 ;
  assign n205 = n204 ^ x1 ;
  assign n206 = n205 ^ n204 ;
  assign n207 = ~x6 & ~x8 ;
  assign n208 = n15 & ~n207 ;
  assign n209 = ~x4 & x9 ;
  assign n210 = x6 & x8 ;
  assign n211 = ~n207 & ~n210 ;
  assign n212 = x9 & n176 ;
  assign n213 = n211 & n212 ;
  assign n214 = ~n209 & ~n213 ;
  assign n215 = x3 & ~x4 ;
  assign n216 = ~x6 & x8 ;
  assign n217 = n215 & ~n216 ;
  assign n218 = ~n11 & n217 ;
  assign n219 = ~n214 & ~n218 ;
  assign n220 = ~n208 & n219 ;
  assign n221 = x6 & ~x9 ;
  assign n222 = ~n145 & ~n221 ;
  assign n223 = ~x4 & ~x8 ;
  assign n224 = x5 & x6 ;
  assign n225 = n223 & ~n224 ;
  assign n226 = ~n222 & n225 ;
  assign n227 = ~n220 & ~n226 ;
  assign n228 = n23 & ~n227 ;
  assign n229 = ~x0 & x9 ;
  assign n230 = ~n32 & n176 ;
  assign n231 = ~n211 & n230 ;
  assign n232 = ~x4 & n231 ;
  assign n233 = ~x5 & x6 ;
  assign n234 = x3 & x6 ;
  assign n235 = ~n233 & ~n234 ;
  assign n236 = ~n103 & ~n215 ;
  assign n237 = n32 & n236 ;
  assign n238 = ~n235 & n237 ;
  assign n239 = ~n232 & ~n238 ;
  assign n240 = n229 & ~n239 ;
  assign n241 = ~x5 & n30 ;
  assign n242 = n14 & n141 ;
  assign n243 = n241 & n242 ;
  assign n244 = x7 & ~n243 ;
  assign n245 = ~n240 & n244 ;
  assign n246 = ~n228 & n245 ;
  assign n247 = ~x0 & ~x9 ;
  assign n248 = ~x2 & ~x6 ;
  assign n249 = n187 ^ x3 ;
  assign n250 = n249 ^ n187 ;
  assign n251 = ~n22 & ~n241 ;
  assign n252 = n251 ^ n187 ;
  assign n253 = ~n250 & ~n252 ;
  assign n254 = n253 ^ n187 ;
  assign n255 = n248 & n254 ;
  assign n265 = ~n20 & n188 ;
  assign n266 = n234 & n265 ;
  assign n256 = x6 ^ x4 ;
  assign n257 = n146 ^ x6 ;
  assign n258 = n257 ^ n146 ;
  assign n259 = n146 ^ n145 ;
  assign n260 = n259 ^ n146 ;
  assign n261 = ~n258 & n260 ;
  assign n262 = n261 ^ n146 ;
  assign n263 = n256 & n262 ;
  assign n264 = n263 ^ n146 ;
  assign n267 = n266 ^ n264 ;
  assign n268 = n267 ^ n266 ;
  assign n269 = n266 ^ x8 ;
  assign n270 = n269 ^ n266 ;
  assign n271 = n268 & ~n270 ;
  assign n272 = n271 ^ n266 ;
  assign n273 = x2 & n272 ;
  assign n274 = n273 ^ n266 ;
  assign n275 = ~n255 & ~n274 ;
  assign n276 = n247 & ~n275 ;
  assign n277 = n94 & n147 ;
  assign n278 = ~n22 & ~n216 ;
  assign n279 = n277 & ~n278 ;
  assign n280 = x4 & x9 ;
  assign n281 = ~x9 & ~n119 ;
  assign n282 = ~n280 & ~n281 ;
  assign n283 = n210 & ~n282 ;
  assign n284 = n283 ^ x5 ;
  assign n285 = n284 ^ n283 ;
  assign n286 = n285 ^ n279 ;
  assign n287 = ~x8 & ~n280 ;
  assign n288 = n236 & n287 ;
  assign n289 = x8 & n209 ;
  assign n290 = x3 & n289 ;
  assign n291 = ~n288 & ~n290 ;
  assign n292 = n291 ^ x6 ;
  assign n293 = ~n291 & ~n292 ;
  assign n294 = n293 ^ n283 ;
  assign n295 = n294 ^ n291 ;
  assign n296 = n286 & ~n295 ;
  assign n297 = n296 ^ n293 ;
  assign n298 = n297 ^ n291 ;
  assign n299 = ~n279 & ~n298 ;
  assign n300 = n299 ^ n279 ;
  assign n301 = n12 & n300 ;
  assign n302 = ~n276 & ~n301 ;
  assign n303 = n246 & n302 ;
  assign n304 = ~x5 & x8 ;
  assign n305 = n12 & n221 ;
  assign n306 = x9 ^ x2 ;
  assign n307 = n306 ^ x9 ;
  assign n308 = n247 ^ x9 ;
  assign n309 = ~n307 & n308 ;
  assign n310 = n309 ^ x9 ;
  assign n311 = ~x6 & n310 ;
  assign n312 = ~n305 & ~n311 ;
  assign n313 = n304 & ~n312 ;
  assign n314 = x2 & x9 ;
  assign n315 = n95 & ~n314 ;
  assign n316 = ~n101 & ~n221 ;
  assign n317 = ~x5 & n316 ;
  assign n318 = n315 & n317 ;
  assign n319 = n229 ^ n11 ;
  assign n320 = x5 & n216 ;
  assign n321 = n320 ^ n319 ;
  assign n322 = n321 ^ n229 ;
  assign n323 = n322 ^ n321 ;
  assign n324 = n321 ^ n305 ;
  assign n325 = n324 ^ n319 ;
  assign n326 = n323 & ~n325 ;
  assign n327 = n326 ^ n305 ;
  assign n328 = n248 & ~n305 ;
  assign n329 = n328 ^ n319 ;
  assign n330 = ~n327 & ~n329 ;
  assign n331 = n330 ^ n328 ;
  assign n332 = ~n319 & n331 ;
  assign n333 = n332 ^ n326 ;
  assign n334 = n333 ^ n11 ;
  assign n335 = n334 ^ n305 ;
  assign n336 = ~n318 & n335 ;
  assign n337 = ~n313 & n336 ;
  assign n338 = n103 & ~n337 ;
  assign n339 = ~n11 & n314 ;
  assign n340 = ~x0 & n211 ;
  assign n341 = n340 ^ n210 ;
  assign n342 = n339 & ~n341 ;
  assign n343 = x5 & ~x9 ;
  assign n344 = n192 & ~n211 ;
  assign n345 = n343 & n344 ;
  assign n346 = ~n342 & ~n345 ;
  assign n347 = n15 & ~n346 ;
  assign n348 = n62 & n101 ;
  assign n349 = x8 & n348 ;
  assign n350 = ~n347 & ~n349 ;
  assign n351 = ~x7 & n350 ;
  assign n352 = ~x2 & ~x4 ;
  assign n353 = n320 ^ x6 ;
  assign n354 = n353 ^ n320 ;
  assign n355 = n320 ^ n304 ;
  assign n356 = n355 ^ n320 ;
  assign n357 = n354 & n356 ;
  assign n358 = n357 ^ n320 ;
  assign n359 = x9 & n358 ;
  assign n360 = n359 ^ n320 ;
  assign n361 = n352 & n360 ;
  assign n362 = ~x4 & x6 ;
  assign n363 = n11 & n362 ;
  assign n364 = n207 & ~n209 ;
  assign n365 = n364 ^ n343 ;
  assign n366 = n364 ^ x2 ;
  assign n367 = n364 & n366 ;
  assign n368 = n367 ^ n364 ;
  assign n369 = ~n365 & n368 ;
  assign n370 = n369 ^ n367 ;
  assign n371 = n370 ^ n364 ;
  assign n372 = n371 ^ x2 ;
  assign n373 = ~n363 & n372 ;
  assign n374 = n373 ^ x2 ;
  assign n375 = ~n361 & ~n374 ;
  assign n376 = n375 ^ x0 ;
  assign n377 = n376 ^ n375 ;
  assign n378 = x4 ^ x2 ;
  assign n379 = n221 ^ x4 ;
  assign n380 = n379 ^ n221 ;
  assign n381 = n221 ^ x9 ;
  assign n382 = n381 ^ n221 ;
  assign n383 = n380 & n382 ;
  assign n384 = n383 ^ n221 ;
  assign n385 = n378 & n384 ;
  assign n386 = n385 ^ n221 ;
  assign n387 = n304 & n386 ;
  assign n388 = n387 ^ n375 ;
  assign n389 = ~n377 & ~n388 ;
  assign n390 = n389 ^ n375 ;
  assign n391 = x3 & ~n390 ;
  assign n392 = n351 & ~n391 ;
  assign n393 = ~n338 & n392 ;
  assign n394 = ~n303 & ~n393 ;
  assign n395 = ~x5 & n280 ;
  assign n396 = n12 & n216 ;
  assign n399 = n396 ^ n32 ;
  assign n400 = n399 ^ n396 ;
  assign n397 = n396 ^ x6 ;
  assign n398 = n397 ^ n396 ;
  assign n401 = n400 ^ n398 ;
  assign n402 = n396 ^ x0 ;
  assign n403 = n402 ^ n396 ;
  assign n404 = n403 ^ n400 ;
  assign n405 = n400 & ~n404 ;
  assign n406 = n405 ^ n400 ;
  assign n407 = n401 & n406 ;
  assign n408 = n407 ^ n405 ;
  assign n409 = n408 ^ n396 ;
  assign n410 = n409 ^ n400 ;
  assign n411 = x3 & n410 ;
  assign n412 = n411 ^ n396 ;
  assign n413 = n395 & n412 ;
  assign n414 = ~n394 & ~n413 ;
  assign n415 = n414 ^ n204 ;
  assign n416 = n206 & n415 ;
  assign n417 = n416 ^ n204 ;
  assign n418 = ~n18 & n417 ;
  assign y0 = ~n418 ;
endmodule
