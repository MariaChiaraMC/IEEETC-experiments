module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n10 = x2 & x3 ;
  assign n11 = x0 & n10 ;
  assign n12 = ~x4 & n11 ;
  assign n13 = ~x5 & ~n12 ;
  assign n14 = x8 ^ x7 ;
  assign n15 = x6 & n14 ;
  assign n16 = n15 ^ x7 ;
  assign n17 = ~n13 & n16 ;
  assign n18 = ~x0 & x3 ;
  assign n19 = n18 ^ x7 ;
  assign n20 = x4 ^ x1 ;
  assign n21 = n20 ^ x4 ;
  assign n22 = x4 ^ x2 ;
  assign n23 = ~n21 & n22 ;
  assign n24 = n23 ^ x4 ;
  assign n25 = n24 ^ n18 ;
  assign n26 = n19 & ~n25 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = n27 ^ x4 ;
  assign n29 = n28 ^ x7 ;
  assign n30 = n18 & ~n29 ;
  assign n31 = n30 ^ n18 ;
  assign n32 = ~n17 & ~n31 ;
  assign y0 = ~n32 ;
endmodule
