module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 ;
  assign n39 = ~x1 & x4 ;
  assign n40 = x0 & ~x1 ;
  assign n29 = x6 & ~x9 ;
  assign n41 = x7 & n29 ;
  assign n42 = ~x2 & ~x5 ;
  assign n43 = n41 & n42 ;
  assign n44 = n40 & n43 ;
  assign n45 = ~n39 & ~n44 ;
  assign n46 = ~x7 & x9 ;
  assign n47 = ~x6 & n46 ;
  assign n48 = x2 & x5 ;
  assign n49 = n47 & n48 ;
  assign n50 = x4 & ~n49 ;
  assign n51 = n50 ^ x2 ;
  assign n52 = n51 ^ n50 ;
  assign n11 = x7 & x9 ;
  assign n12 = ~x5 & n11 ;
  assign n13 = x6 & n12 ;
  assign n53 = n50 ^ n13 ;
  assign n54 = n53 ^ n50 ;
  assign n55 = ~n52 & n54 ;
  assign n56 = n55 ^ n50 ;
  assign n57 = ~x0 & ~n56 ;
  assign n58 = n57 ^ n50 ;
  assign n59 = ~n45 & ~n58 ;
  assign n14 = ~x1 & ~x2 ;
  assign n15 = n13 & n14 ;
  assign n16 = ~x6 & ~x7 ;
  assign n17 = ~x9 & n16 ;
  assign n18 = x1 & x2 ;
  assign n19 = n17 & n18 ;
  assign n20 = ~x0 & ~n19 ;
  assign n21 = x5 & ~n20 ;
  assign n22 = ~n15 & ~n21 ;
  assign n23 = x5 & x7 ;
  assign n24 = x0 & n23 ;
  assign n25 = ~x2 & ~x6 ;
  assign n26 = x1 & x9 ;
  assign n27 = n25 & n26 ;
  assign n28 = n27 ^ n23 ;
  assign n30 = ~x1 & x2 ;
  assign n31 = n29 & n30 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = ~n28 & n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n24 & n34 ;
  assign n36 = n35 ^ x0 ;
  assign n37 = ~x4 & ~n36 ;
  assign n38 = ~n22 & n37 ;
  assign n60 = n59 ^ n38 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = ~x0 & n42 ;
  assign n63 = n17 & n62 ;
  assign n64 = x6 & x7 ;
  assign n65 = x0 & x9 ;
  assign n66 = n48 & n65 ;
  assign n67 = n64 & n66 ;
  assign n68 = ~n63 & ~n67 ;
  assign n69 = n39 & ~n68 ;
  assign n70 = n69 ^ n59 ;
  assign n71 = n70 ^ n59 ;
  assign n72 = ~n61 & ~n71 ;
  assign n73 = n72 ^ n59 ;
  assign n74 = x8 & ~n73 ;
  assign n75 = n74 ^ n59 ;
  assign n226 = x8 & n17 ;
  assign n115 = x8 & ~x9 ;
  assign n100 = ~x8 & x9 ;
  assign n356 = ~x7 & n100 ;
  assign n357 = ~n115 & ~n356 ;
  assign n358 = n357 ^ n41 ;
  assign n359 = n358 ^ n41 ;
  assign n360 = n41 ^ x6 ;
  assign n361 = n360 ^ n41 ;
  assign n362 = ~n359 & ~n361 ;
  assign n363 = n362 ^ n41 ;
  assign n364 = x5 & n363 ;
  assign n365 = n364 ^ n41 ;
  assign n366 = ~n226 & ~n365 ;
  assign n367 = ~x0 & x1 ;
  assign n368 = ~n366 & n367 ;
  assign n86 = ~x8 & ~x9 ;
  assign n96 = x6 & ~x7 ;
  assign n222 = n86 & n96 ;
  assign n369 = x1 & ~x5 ;
  assign n370 = n222 & n369 ;
  assign n76 = x0 & x1 ;
  assign n87 = ~x6 & x7 ;
  assign n197 = n87 & n115 ;
  assign n371 = n76 & n197 ;
  assign n372 = n371 ^ x5 ;
  assign n373 = n372 ^ n371 ;
  assign n374 = n373 ^ n370 ;
  assign n219 = x9 ^ x7 ;
  assign n375 = ~x0 & ~x1 ;
  assign n376 = n375 ^ x9 ;
  assign n377 = n376 ^ x8 ;
  assign n378 = n377 ^ n375 ;
  assign n379 = n378 ^ n219 ;
  assign n380 = n76 ^ x8 ;
  assign n381 = n76 & ~n380 ;
  assign n382 = n381 ^ n375 ;
  assign n383 = n382 ^ n76 ;
  assign n384 = n379 & n383 ;
  assign n385 = n384 ^ n381 ;
  assign n386 = n385 ^ n76 ;
  assign n387 = n219 & n386 ;
  assign n388 = n387 ^ x6 ;
  assign n389 = n387 & n388 ;
  assign n390 = n389 ^ n371 ;
  assign n391 = n390 ^ n387 ;
  assign n392 = ~n374 & n391 ;
  assign n393 = n392 ^ n389 ;
  assign n394 = n393 ^ n387 ;
  assign n395 = ~n370 & n394 ;
  assign n396 = n395 ^ n370 ;
  assign n397 = ~n368 & ~n396 ;
  assign n398 = ~x2 & ~n397 ;
  assign n399 = ~x4 & n398 ;
  assign n116 = ~x4 & n115 ;
  assign n164 = ~x1 & x6 ;
  assign n400 = x5 ^ x0 ;
  assign n401 = x7 ^ x5 ;
  assign n402 = ~n400 & ~n401 ;
  assign n403 = n164 & n402 ;
  assign n404 = n116 & n403 ;
  assign n405 = ~n399 & ~n404 ;
  assign n247 = ~x0 & x4 ;
  assign n77 = x8 & x9 ;
  assign n143 = n86 ^ n77 ;
  assign n406 = x5 & n143 ;
  assign n407 = n406 ^ n77 ;
  assign n408 = n247 & n407 ;
  assign n409 = n64 & n408 ;
  assign n104 = ~x6 & n77 ;
  assign n105 = ~x7 & n104 ;
  assign n410 = n105 ^ x0 ;
  assign n411 = n410 ^ n105 ;
  assign n88 = n86 & n87 ;
  assign n412 = x7 & n77 ;
  assign n413 = ~n88 & ~n412 ;
  assign n414 = n413 ^ x6 ;
  assign n415 = n414 ^ n413 ;
  assign n416 = n413 ^ n356 ;
  assign n417 = n416 ^ n413 ;
  assign n418 = ~n415 & n417 ;
  assign n419 = n418 ^ n413 ;
  assign n420 = x4 & ~n419 ;
  assign n421 = n420 ^ n413 ;
  assign n422 = n421 ^ n105 ;
  assign n423 = n411 & ~n422 ;
  assign n424 = n423 ^ n105 ;
  assign n425 = n369 & n424 ;
  assign n426 = ~n409 & ~n425 ;
  assign n427 = ~x4 & ~x5 ;
  assign n428 = x8 ^ x6 ;
  assign n429 = x0 & n428 ;
  assign n430 = n429 ^ x6 ;
  assign n431 = n427 & ~n430 ;
  assign n432 = ~x9 & n431 ;
  assign n131 = ~x0 & ~x7 ;
  assign n79 = ~x4 & x6 ;
  assign n327 = x8 & ~n79 ;
  assign n433 = x5 & x9 ;
  assign n434 = ~n327 & n433 ;
  assign n250 = x4 & x6 ;
  assign n435 = n115 & n250 ;
  assign n436 = ~x7 & ~n435 ;
  assign n437 = ~n434 & n436 ;
  assign n438 = ~n131 & ~n437 ;
  assign n439 = x4 & ~x5 ;
  assign n440 = ~x0 & x6 ;
  assign n441 = ~x8 & n440 ;
  assign n442 = ~n104 & ~n441 ;
  assign n443 = n439 & ~n442 ;
  assign n444 = ~n438 & ~n443 ;
  assign n445 = ~n432 & n444 ;
  assign n168 = ~x6 & ~x8 ;
  assign n446 = n65 & n439 ;
  assign n447 = n168 & n446 ;
  assign n83 = ~x0 & x8 ;
  assign n278 = x4 & ~x9 ;
  assign n268 = x4 & ~x6 ;
  assign n280 = ~n79 & ~n268 ;
  assign n448 = ~n280 & n433 ;
  assign n449 = ~n278 & ~n448 ;
  assign n450 = n83 & ~n449 ;
  assign n451 = x7 & ~n450 ;
  assign n452 = ~n447 & n451 ;
  assign n453 = ~n445 & ~n452 ;
  assign n454 = n453 ^ x1 ;
  assign n455 = n454 ^ n453 ;
  assign n456 = n455 ^ n426 ;
  assign n457 = n23 & n116 ;
  assign n267 = x7 & x8 ;
  assign n460 = n267 ^ n86 ;
  assign n461 = n460 ^ n267 ;
  assign n458 = n267 ^ x7 ;
  assign n459 = n458 ^ n267 ;
  assign n462 = n461 ^ n459 ;
  assign n463 = n267 ^ x5 ;
  assign n464 = n463 ^ n267 ;
  assign n465 = n464 ^ n461 ;
  assign n466 = n461 & ~n465 ;
  assign n467 = n466 ^ n461 ;
  assign n468 = ~n462 & n467 ;
  assign n469 = n468 ^ n466 ;
  assign n470 = n469 ^ n267 ;
  assign n471 = n470 ^ n461 ;
  assign n472 = x4 & n471 ;
  assign n473 = n472 ^ n267 ;
  assign n474 = n473 ^ x0 ;
  assign n475 = n474 ^ n473 ;
  assign n476 = n475 ^ n457 ;
  assign n477 = x5 & n86 ;
  assign n478 = ~n12 & ~n477 ;
  assign n479 = n478 ^ x4 ;
  assign n480 = x4 & ~n479 ;
  assign n481 = n480 ^ n473 ;
  assign n482 = n481 ^ x4 ;
  assign n483 = n476 & n482 ;
  assign n484 = n483 ^ n480 ;
  assign n485 = n484 ^ x4 ;
  assign n486 = ~n457 & n485 ;
  assign n487 = n486 ^ n457 ;
  assign n488 = n487 ^ x6 ;
  assign n489 = x6 & n488 ;
  assign n490 = n489 ^ n453 ;
  assign n491 = n490 ^ x6 ;
  assign n492 = n456 & n491 ;
  assign n493 = n492 ^ n489 ;
  assign n494 = n493 ^ x6 ;
  assign n495 = n426 & n494 ;
  assign n496 = n495 ^ n426 ;
  assign n497 = x2 & ~n496 ;
  assign n270 = x7 ^ x6 ;
  assign n322 = x8 & n270 ;
  assign n498 = x9 & n40 ;
  assign n499 = n322 & n498 ;
  assign n89 = n40 & n88 ;
  assign n500 = ~x5 & ~n89 ;
  assign n501 = ~n499 & n500 ;
  assign n502 = x9 ^ x8 ;
  assign n503 = n64 ^ x9 ;
  assign n504 = n503 ^ n64 ;
  assign n505 = n504 ^ n502 ;
  assign n506 = n96 ^ n76 ;
  assign n507 = n76 & n506 ;
  assign n508 = n507 ^ n64 ;
  assign n509 = n508 ^ n76 ;
  assign n510 = ~n505 & n509 ;
  assign n511 = n510 ^ n507 ;
  assign n512 = n511 ^ n76 ;
  assign n513 = n502 & n512 ;
  assign n514 = n501 & ~n513 ;
  assign n515 = ~x2 & x4 ;
  assign n516 = n88 & n375 ;
  assign n329 = x7 & n168 ;
  assign n517 = n26 & n329 ;
  assign n518 = x5 & ~n517 ;
  assign n519 = ~n516 & n518 ;
  assign n520 = n515 & ~n519 ;
  assign n521 = ~n514 & n520 ;
  assign n522 = x6 & n86 ;
  assign n523 = ~n104 & ~n522 ;
  assign n524 = ~x5 & n131 ;
  assign n525 = n39 & n524 ;
  assign n526 = ~n523 & n525 ;
  assign n527 = ~n521 & ~n526 ;
  assign n528 = ~n497 & n527 ;
  assign n529 = n405 & n528 ;
  assign n78 = ~x7 & n77 ;
  assign n80 = n78 & n79 ;
  assign n81 = n76 & n80 ;
  assign n82 = x1 & x4 ;
  assign n84 = n82 & n83 ;
  assign n85 = n41 & n84 ;
  assign n90 = x4 & n89 ;
  assign n91 = ~n85 & ~n90 ;
  assign n92 = ~n81 & n91 ;
  assign n93 = x2 & ~n92 ;
  assign n94 = ~x4 & n87 ;
  assign n95 = ~x1 & n94 ;
  assign n97 = n82 & n96 ;
  assign n98 = ~n95 & ~n97 ;
  assign n99 = ~x0 & ~x2 ;
  assign n101 = n99 & n100 ;
  assign n102 = ~n98 & n101 ;
  assign n103 = n102 ^ n93 ;
  assign n106 = ~n25 & ~n105 ;
  assign n107 = x7 & n86 ;
  assign n108 = ~x2 & ~n107 ;
  assign n109 = n82 & ~n108 ;
  assign n110 = ~n106 & n109 ;
  assign n111 = x7 & n99 ;
  assign n112 = n100 ^ x1 ;
  assign n113 = n100 ^ x4 ;
  assign n114 = n113 ^ x4 ;
  assign n117 = n116 ^ x4 ;
  assign n118 = ~n114 & n117 ;
  assign n119 = n118 ^ x4 ;
  assign n120 = ~n112 & ~n119 ;
  assign n121 = n120 ^ x1 ;
  assign n122 = n121 ^ n39 ;
  assign n123 = n122 ^ n121 ;
  assign n124 = n121 ^ n86 ;
  assign n125 = n124 ^ n121 ;
  assign n126 = n123 & n125 ;
  assign n127 = n126 ^ n121 ;
  assign n128 = x6 & ~n127 ;
  assign n129 = n128 ^ n121 ;
  assign n130 = n111 & ~n129 ;
  assign n132 = n77 ^ x2 ;
  assign n133 = n132 ^ x6 ;
  assign n140 = n133 ^ n77 ;
  assign n134 = n133 ^ x1 ;
  assign n135 = n134 ^ n77 ;
  assign n136 = x6 ^ x1 ;
  assign n137 = n136 ^ x1 ;
  assign n138 = n137 ^ n135 ;
  assign n139 = ~n135 & ~n138 ;
  assign n141 = n140 ^ n139 ;
  assign n142 = n141 ^ n135 ;
  assign n144 = n139 ^ n135 ;
  assign n145 = n143 & ~n144 ;
  assign n146 = n145 ^ n77 ;
  assign n147 = ~n142 & n146 ;
  assign n148 = n147 ^ n77 ;
  assign n149 = n148 ^ n77 ;
  assign n150 = n149 ^ x4 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = n151 ^ n131 ;
  assign n153 = x2 & ~x6 ;
  assign n154 = n30 ^ x6 ;
  assign n155 = n154 ^ n30 ;
  assign n156 = n30 ^ x1 ;
  assign n157 = n156 ^ n30 ;
  assign n158 = ~n155 & ~n157 ;
  assign n159 = n158 ^ n30 ;
  assign n160 = ~x8 & n159 ;
  assign n161 = n160 ^ n30 ;
  assign n162 = ~n153 & n161 ;
  assign n163 = ~x9 & n162 ;
  assign n165 = n164 ^ x9 ;
  assign n166 = n18 ^ x8 ;
  assign n167 = n166 ^ x8 ;
  assign n169 = n168 ^ x8 ;
  assign n170 = n167 & n169 ;
  assign n171 = n170 ^ x8 ;
  assign n172 = n171 ^ n164 ;
  assign n173 = ~n165 & ~n172 ;
  assign n174 = n173 ^ n170 ;
  assign n175 = n174 ^ x8 ;
  assign n176 = n175 ^ x9 ;
  assign n177 = ~n164 & n176 ;
  assign n178 = n177 ^ n164 ;
  assign n179 = n178 ^ n163 ;
  assign n180 = ~n163 & ~n179 ;
  assign n181 = n180 ^ n149 ;
  assign n182 = n181 ^ n163 ;
  assign n183 = ~n152 & n182 ;
  assign n184 = n183 ^ n180 ;
  assign n185 = n184 ^ n163 ;
  assign n186 = n131 & ~n185 ;
  assign n187 = n186 ^ n131 ;
  assign n188 = ~n130 & ~n187 ;
  assign n194 = x7 & ~x9 ;
  assign n195 = x2 & ~n194 ;
  assign n189 = ~x2 & ~n46 ;
  assign n190 = ~x4 & ~x6 ;
  assign n191 = ~x8 & n190 ;
  assign n192 = ~n189 & n191 ;
  assign n193 = n192 ^ x4 ;
  assign n196 = n195 ^ n193 ;
  assign n204 = n196 ^ n193 ;
  assign n198 = n197 ^ n196 ;
  assign n199 = n198 ^ n193 ;
  assign n200 = n196 ^ n192 ;
  assign n201 = n200 ^ n197 ;
  assign n202 = n201 ^ n199 ;
  assign n203 = n199 & ~n202 ;
  assign n205 = n204 ^ n203 ;
  assign n206 = n205 ^ n199 ;
  assign n207 = ~x8 & n64 ;
  assign n208 = ~n29 & ~n207 ;
  assign n209 = n208 ^ n193 ;
  assign n210 = n203 ^ n199 ;
  assign n211 = n209 & n210 ;
  assign n212 = n211 ^ n193 ;
  assign n213 = ~n206 & n212 ;
  assign n214 = n213 ^ n193 ;
  assign n215 = n214 ^ x4 ;
  assign n216 = n215 ^ n193 ;
  assign n217 = n216 ^ x1 ;
  assign n218 = n217 ^ n216 ;
  assign n220 = n190 & ~n219 ;
  assign n221 = x8 & n220 ;
  assign n227 = ~x4 & ~x8 ;
  assign n228 = n11 & n227 ;
  assign n229 = ~n226 & ~n228 ;
  assign n223 = ~n41 & ~n47 ;
  assign n224 = x8 & ~n223 ;
  assign n225 = ~n222 & ~n224 ;
  assign n230 = n229 ^ n225 ;
  assign n231 = n230 ^ n229 ;
  assign n232 = n229 ^ x4 ;
  assign n233 = n232 ^ n229 ;
  assign n234 = ~n231 & n233 ;
  assign n235 = n234 ^ n229 ;
  assign n236 = ~x2 & ~n235 ;
  assign n237 = n236 ^ n229 ;
  assign n238 = ~n221 & n237 ;
  assign n239 = n238 ^ n216 ;
  assign n240 = ~n218 & ~n239 ;
  assign n241 = n240 ^ n216 ;
  assign n242 = x0 & n241 ;
  assign n243 = n188 & ~n242 ;
  assign n244 = ~n110 & n243 ;
  assign n245 = n244 ^ x5 ;
  assign n246 = n245 ^ n244 ;
  assign n251 = n46 & n250 ;
  assign n252 = n251 ^ x0 ;
  assign n248 = n47 & n247 ;
  assign n249 = n248 ^ x8 ;
  assign n253 = n252 ^ n249 ;
  assign n254 = n252 ^ n248 ;
  assign n255 = n254 ^ x0 ;
  assign n256 = n253 & ~n255 ;
  assign n257 = n256 ^ n248 ;
  assign n258 = ~n94 & ~n248 ;
  assign n259 = n258 ^ x0 ;
  assign n260 = ~n257 & n259 ;
  assign n261 = n260 ^ n258 ;
  assign n262 = x0 & n261 ;
  assign n263 = n262 ^ n256 ;
  assign n264 = n263 ^ x8 ;
  assign n265 = n264 ^ n248 ;
  assign n266 = n30 & n265 ;
  assign n269 = n267 & n268 ;
  assign n271 = x6 ^ x2 ;
  assign n272 = n270 & ~n271 ;
  assign n273 = n272 ^ x2 ;
  assign n274 = n227 & n273 ;
  assign n275 = ~n269 & ~n274 ;
  assign n276 = x0 & n26 ;
  assign n277 = ~n275 & n276 ;
  assign n279 = n14 & n267 ;
  assign n281 = n280 ^ x4 ;
  assign n282 = n281 ^ n280 ;
  assign n283 = n280 ^ x9 ;
  assign n284 = n283 ^ n280 ;
  assign n285 = ~n282 & n284 ;
  assign n286 = n285 ^ n280 ;
  assign n287 = x0 & ~n286 ;
  assign n288 = n287 ^ n280 ;
  assign n289 = n279 & ~n288 ;
  assign n290 = ~n278 & n289 ;
  assign n291 = ~n277 & ~n290 ;
  assign n292 = ~n266 & n291 ;
  assign n293 = n153 & n227 ;
  assign n296 = n293 ^ n250 ;
  assign n297 = n296 ^ n293 ;
  assign n294 = n293 ^ x8 ;
  assign n295 = n294 ^ n293 ;
  assign n298 = n297 ^ n295 ;
  assign n299 = n293 ^ x2 ;
  assign n300 = n299 ^ n293 ;
  assign n301 = n300 ^ n297 ;
  assign n302 = n297 & ~n301 ;
  assign n303 = n302 ^ n297 ;
  assign n304 = n298 & n303 ;
  assign n305 = n304 ^ n302 ;
  assign n306 = n305 ^ n293 ;
  assign n307 = n306 ^ n297 ;
  assign n308 = ~x7 & n307 ;
  assign n309 = n308 ^ n293 ;
  assign n310 = x1 & n309 ;
  assign n311 = n96 & n227 ;
  assign n312 = n250 & n267 ;
  assign n313 = ~n311 & ~n312 ;
  assign n314 = x2 & ~n313 ;
  assign n315 = ~n310 & ~n314 ;
  assign n316 = n315 ^ x0 ;
  assign n317 = n316 ^ n315 ;
  assign n318 = n317 ^ x9 ;
  assign n319 = n30 & n79 ;
  assign n320 = x7 & n319 ;
  assign n321 = ~x4 & ~n16 ;
  assign n323 = ~n227 & ~n322 ;
  assign n324 = ~n321 & ~n323 ;
  assign n325 = n324 ^ x1 ;
  assign n326 = n325 ^ n324 ;
  assign n328 = ~x7 & x8 ;
  assign n330 = ~n328 & ~n329 ;
  assign n331 = ~n327 & ~n330 ;
  assign n332 = n331 ^ n324 ;
  assign n333 = n326 & n332 ;
  assign n334 = n333 ^ n324 ;
  assign n335 = ~x2 & n334 ;
  assign n336 = n335 ^ n320 ;
  assign n337 = ~n320 & n336 ;
  assign n338 = n337 ^ n315 ;
  assign n339 = n338 ^ n320 ;
  assign n340 = ~n318 & ~n339 ;
  assign n341 = n340 ^ n337 ;
  assign n342 = n341 ^ n320 ;
  assign n343 = ~x9 & ~n342 ;
  assign n344 = n343 ^ x9 ;
  assign n345 = n292 & n344 ;
  assign n346 = n345 ^ n244 ;
  assign n347 = ~n246 & n346 ;
  assign n348 = n347 ^ n244 ;
  assign n349 = n348 ^ n93 ;
  assign n350 = n103 & ~n349 ;
  assign n351 = n350 ^ n347 ;
  assign n352 = n351 ^ n244 ;
  assign n353 = n352 ^ n102 ;
  assign n354 = ~n93 & ~n353 ;
  assign n355 = n354 ^ n93 ;
  assign n530 = n529 ^ n355 ;
  assign n531 = ~x3 & ~n530 ;
  assign n532 = n531 ^ n355 ;
  assign n533 = ~n75 & ~n532 ;
  assign y0 = ~n533 ;
endmodule
