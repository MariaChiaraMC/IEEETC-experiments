module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 ;
  assign n17 = x6 & x7 ;
  assign n18 = ~x10 & ~x11 ;
  assign n19 = ~x8 & ~x9 ;
  assign n20 = x8 & x9 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = n18 & n21 ;
  assign n23 = n17 & ~n22 ;
  assign n24 = x4 & ~n23 ;
  assign n25 = ~x14 & ~x15 ;
  assign n27 = ~x12 & ~x13 ;
  assign n28 = x5 & ~n17 ;
  assign n29 = n27 & ~n28 ;
  assign n26 = ~x6 & x7 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n29 ^ x5 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = ~n31 & n33 ;
  assign n35 = n34 ^ n29 ;
  assign n36 = n25 & ~n35 ;
  assign n37 = n36 ^ n29 ;
  assign n38 = n24 & n37 ;
  assign n39 = ~x4 & ~x5 ;
  assign n40 = ~x8 & x9 ;
  assign n41 = n17 & n40 ;
  assign n42 = n39 & n41 ;
  assign n43 = ~n38 & ~n42 ;
  assign n44 = x6 ^ x4 ;
  assign n45 = n22 ^ x6 ;
  assign n46 = n45 ^ n22 ;
  assign n47 = n46 ^ n44 ;
  assign n48 = x10 & x11 ;
  assign n49 = ~n18 & ~n48 ;
  assign n50 = n49 ^ n19 ;
  assign n51 = n19 & n50 ;
  assign n52 = n51 ^ n22 ;
  assign n53 = n52 ^ n19 ;
  assign n54 = n47 & n53 ;
  assign n55 = n54 ^ n51 ;
  assign n56 = n55 ^ n19 ;
  assign n57 = ~n44 & n56 ;
  assign n58 = n57 ^ x4 ;
  assign n59 = x7 & n58 ;
  assign n60 = x7 ^ x4 ;
  assign n61 = x6 & ~x10 ;
  assign n62 = x11 & n61 ;
  assign n63 = x14 & n62 ;
  assign n64 = n63 ^ x7 ;
  assign n65 = n64 ^ n63 ;
  assign n66 = ~x6 & ~n21 ;
  assign n67 = n18 & ~n66 ;
  assign n68 = n67 ^ n63 ;
  assign n69 = n65 & ~n68 ;
  assign n70 = n69 ^ n63 ;
  assign n71 = n60 & n70 ;
  assign n72 = n71 ^ x4 ;
  assign n73 = ~n59 & n72 ;
  assign n74 = n27 & ~n73 ;
  assign n75 = x15 & ~n74 ;
  assign n76 = ~x12 & x14 ;
  assign n77 = x7 & n76 ;
  assign n78 = x9 ^ x8 ;
  assign n79 = n78 ^ x10 ;
  assign n80 = n79 ^ x11 ;
  assign n81 = n80 ^ x11 ;
  assign n82 = n80 ^ x6 ;
  assign n84 = n82 ^ x10 ;
  assign n85 = n84 ^ x11 ;
  assign n83 = n82 ^ x11 ;
  assign n86 = n85 ^ n83 ;
  assign n87 = n86 ^ n81 ;
  assign n88 = ~n81 & ~n87 ;
  assign n89 = n88 ^ n82 ;
  assign n90 = n89 ^ n81 ;
  assign n91 = x9 & ~n85 ;
  assign n92 = n91 ^ n82 ;
  assign n93 = ~n90 & n92 ;
  assign n94 = n93 ^ n82 ;
  assign n95 = n94 ^ n80 ;
  assign n96 = n77 & ~n95 ;
  assign n97 = x6 & x10 ;
  assign n98 = x12 & ~x14 ;
  assign n99 = ~n76 & ~n98 ;
  assign n100 = n97 & ~n99 ;
  assign n101 = ~x11 & n100 ;
  assign n102 = ~x13 & ~n101 ;
  assign n105 = ~x14 & n17 ;
  assign n103 = n17 & ~n99 ;
  assign n104 = x11 & n103 ;
  assign n106 = n105 ^ n104 ;
  assign n107 = x12 ^ x10 ;
  assign n108 = n107 ^ x10 ;
  assign n109 = n108 ^ n106 ;
  assign n110 = x8 & ~x9 ;
  assign n111 = n110 ^ x10 ;
  assign n112 = n111 ^ n104 ;
  assign n113 = n104 & ~n112 ;
  assign n114 = n113 ^ x10 ;
  assign n115 = n114 ^ n104 ;
  assign n116 = ~n109 & n115 ;
  assign n117 = n116 ^ n113 ;
  assign n118 = n117 ^ n104 ;
  assign n119 = n106 & n118 ;
  assign n120 = n119 ^ n105 ;
  assign n121 = n102 & ~n120 ;
  assign n122 = ~n96 & n121 ;
  assign n123 = x4 & ~n122 ;
  assign n124 = ~x15 & ~n123 ;
  assign n125 = n62 & n98 ;
  assign n126 = x13 & ~n125 ;
  assign n127 = ~n105 & n126 ;
  assign n128 = ~n124 & ~n127 ;
  assign n129 = ~x6 & n19 ;
  assign n130 = ~n18 & ~n129 ;
  assign n131 = ~n18 & ~n20 ;
  assign n132 = n66 & ~n131 ;
  assign n133 = ~n48 & ~n132 ;
  assign n134 = ~n130 & n133 ;
  assign n135 = x7 & ~n134 ;
  assign n136 = x14 ^ x4 ;
  assign n137 = n136 ^ x4 ;
  assign n138 = n27 ^ x4 ;
  assign n139 = n137 & ~n138 ;
  assign n140 = n139 ^ x4 ;
  assign n141 = x4 & ~n26 ;
  assign n142 = n141 ^ n135 ;
  assign n143 = n140 & ~n142 ;
  assign n144 = n143 ^ n141 ;
  assign n145 = ~n135 & n144 ;
  assign n146 = n145 ^ n135 ;
  assign n147 = ~n128 & n146 ;
  assign n148 = x5 & ~n147 ;
  assign n149 = ~n75 & n148 ;
  assign n150 = n43 & ~n149 ;
  assign n151 = ~x0 & ~x3 ;
  assign n152 = ~x1 & n151 ;
  assign n153 = ~x2 & n152 ;
  assign n154 = ~n150 & n153 ;
  assign y0 = n154 ;
endmodule
