module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 ;
  assign n9 = x1 & ~x5 ;
  assign n10 = x4 & n9 ;
  assign n11 = n10 ^ x6 ;
  assign n18 = n11 ^ n10 ;
  assign n12 = n11 ^ x1 ;
  assign n13 = n12 ^ n10 ;
  assign n14 = x2 ^ x1 ;
  assign n15 = n14 ^ x1 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = n13 & n16 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = n19 ^ n13 ;
  assign n21 = ~x4 & x5 ;
  assign n22 = n21 ^ n10 ;
  assign n23 = n17 ^ n13 ;
  assign n24 = n22 & n23 ;
  assign n25 = n24 ^ n10 ;
  assign n26 = ~n20 & n25 ;
  assign n27 = n26 ^ n10 ;
  assign n28 = n27 ^ n10 ;
  assign n29 = ~x0 & ~n28 ;
  assign n30 = ~x2 & n21 ;
  assign n31 = ~x1 & n30 ;
  assign n32 = ~x6 & n31 ;
  assign n33 = n32 ^ x3 ;
  assign n34 = n33 ^ n32 ;
  assign n35 = n34 ^ x7 ;
  assign n36 = x2 & n10 ;
  assign n37 = x6 & n36 ;
  assign n38 = n37 ^ x0 ;
  assign n39 = ~n37 & ~n38 ;
  assign n40 = n39 ^ n32 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = ~n35 & n41 ;
  assign n43 = n42 ^ n39 ;
  assign n44 = n43 ^ n37 ;
  assign n45 = x7 & ~n44 ;
  assign n46 = n45 ^ x7 ;
  assign n47 = ~n29 & n46 ;
  assign n48 = ~x0 & ~x7 ;
  assign n49 = n36 ^ n31 ;
  assign n50 = x6 & n49 ;
  assign n51 = n50 ^ n36 ;
  assign n52 = n48 & n51 ;
  assign n53 = ~x3 & n52 ;
  assign n54 = ~n47 & ~n53 ;
  assign y0 = ~n54 ;
endmodule
