module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 ;
  assign n17 = x4 & x5 ;
  assign n18 = x3 & ~x6 ;
  assign n19 = x1 & ~n18 ;
  assign n20 = n17 & ~n19 ;
  assign n21 = x5 & ~x6 ;
  assign n22 = x1 & ~n21 ;
  assign n23 = ~n17 & ~n22 ;
  assign n24 = x10 & ~x11 ;
  assign n25 = ~x8 & ~x12 ;
  assign n26 = x9 & n25 ;
  assign n27 = ~x3 & n26 ;
  assign n28 = n24 & n27 ;
  assign n29 = ~n23 & n28 ;
  assign n30 = x14 & x15 ;
  assign n31 = x14 ^ x13 ;
  assign n32 = n31 ^ x15 ;
  assign n33 = n30 & n32 ;
  assign n34 = n33 ^ n32 ;
  assign n35 = n29 & n34 ;
  assign n36 = ~n20 & ~n35 ;
  assign y0 = ~n36 ;
endmodule
