module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n7 = x5 ^ x3 ;
  assign n8 = x1 ^ x0 ;
  assign n9 = n8 ^ x5 ;
  assign n10 = ~x5 & n9 ;
  assign n11 = n10 ^ x5 ;
  assign n12 = n7 & ~n11 ;
  assign n13 = n12 ^ n10 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = n14 ^ n8 ;
  assign n16 = ~x1 & n15 ;
  assign n17 = n16 ^ n8 ;
  assign n18 = n17 ^ x3 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = n19 ^ n18 ;
  assign n24 = n18 ^ x4 ;
  assign n25 = ~n18 & ~n24 ;
  assign n21 = ~x0 & ~x1 ;
  assign n22 = x3 & ~n21 ;
  assign n28 = n25 ^ n22 ;
  assign n23 = n22 ^ n20 ;
  assign n26 = n25 ^ n18 ;
  assign n27 = n23 & ~n26 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n20 & n29 ;
  assign n31 = n30 ^ n25 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = n32 ^ x3 ;
  assign y0 = n33 ;
endmodule
