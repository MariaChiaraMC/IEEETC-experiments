module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 ;
  assign n8 = x3 ^ x0 ;
  assign n7 = x2 ^ x0 ;
  assign n9 = n8 ^ n7 ;
  assign n10 = n9 ^ x1 ;
  assign n11 = n10 ^ x4 ;
  assign n12 = n11 ^ n10 ;
  assign n18 = n10 ^ n8 ;
  assign n19 = n18 ^ x0 ;
  assign n14 = n11 ^ x1 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = n15 ^ x0 ;
  assign n13 = n12 ^ x0 ;
  assign n17 = n16 ^ n13 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = ~n12 & n20 ;
  assign n22 = n21 ^ n12 ;
  assign n23 = n22 ^ x0 ;
  assign n24 = n19 ^ x0 ;
  assign n30 = n16 ^ n8 ;
  assign n31 = ~x0 & n30 ;
  assign n25 = n8 ^ x5 ;
  assign n26 = n25 ^ n11 ;
  assign n27 = n16 ^ x0 ;
  assign n28 = n27 ^ n19 ;
  assign n29 = ~n26 & ~n28 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = n32 ^ n26 ;
  assign n34 = n33 ^ n8 ;
  assign n35 = n34 ^ n12 ;
  assign n36 = n35 ^ n16 ;
  assign n37 = n36 ^ n19 ;
  assign n38 = n24 & ~n37 ;
  assign n39 = n38 ^ n29 ;
  assign n40 = n39 ^ n26 ;
  assign n41 = n40 ^ n12 ;
  assign n42 = n41 ^ n16 ;
  assign n43 = n23 & ~n42 ;
  assign n44 = n43 ^ n31 ;
  assign n45 = n44 ^ n8 ;
  assign n46 = n45 ^ x0 ;
  assign n47 = n46 ^ x3 ;
  assign n48 = n47 ^ n8 ;
  assign y0 = n48 ;
endmodule
