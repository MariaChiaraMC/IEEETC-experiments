module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 ;
  assign n11 = x4 & ~x7 ;
  assign n12 = ~x0 & ~x2 ;
  assign n13 = n11 & n12 ;
  assign n14 = x1 & x3 ;
  assign n15 = x8 & ~x9 ;
  assign n16 = n14 & n15 ;
  assign n17 = n13 & n16 ;
  assign n18 = ~x2 & n14 ;
  assign n19 = ~x4 & ~x7 ;
  assign n20 = x8 & n19 ;
  assign n21 = n18 & n20 ;
  assign n22 = ~x3 & ~x8 ;
  assign n23 = ~x1 & x2 ;
  assign n24 = x4 & x7 ;
  assign n25 = n23 & n24 ;
  assign n26 = n22 & n25 ;
  assign n27 = ~n21 & ~n26 ;
  assign n28 = x0 & x9 ;
  assign n29 = ~n27 & n28 ;
  assign n30 = ~n17 & ~n29 ;
  assign n31 = ~x6 & ~n30 ;
  assign n32 = x2 & x7 ;
  assign n33 = ~x4 & x6 ;
  assign n34 = n32 & n33 ;
  assign n35 = x0 & n34 ;
  assign n36 = ~x1 & x9 ;
  assign n37 = n36 ^ x3 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = x1 & ~x9 ;
  assign n40 = n39 ^ n36 ;
  assign n41 = ~n38 & n40 ;
  assign n42 = n41 ^ n36 ;
  assign n43 = n35 & n42 ;
  assign n44 = ~x2 & ~x3 ;
  assign n45 = ~x7 & ~x9 ;
  assign n46 = x4 & ~x6 ;
  assign n47 = n45 & n46 ;
  assign n48 = ~x1 & n47 ;
  assign n49 = x7 & ~n36 ;
  assign n50 = x6 ^ x4 ;
  assign n51 = n39 ^ x4 ;
  assign n52 = ~n50 & ~n51 ;
  assign n53 = n49 & n52 ;
  assign n54 = ~n48 & ~n53 ;
  assign n55 = n44 & ~n54 ;
  assign n56 = x7 ^ x4 ;
  assign n57 = x4 ^ x3 ;
  assign n58 = n57 ^ n56 ;
  assign n59 = x7 ^ x6 ;
  assign n60 = n59 ^ x6 ;
  assign n61 = ~x6 & x9 ;
  assign n62 = n61 ^ x6 ;
  assign n63 = ~n60 & n62 ;
  assign n64 = n63 ^ x6 ;
  assign n65 = n64 ^ n56 ;
  assign n66 = ~n58 & ~n65 ;
  assign n67 = n66 ^ n63 ;
  assign n68 = n67 ^ x6 ;
  assign n69 = n68 ^ n57 ;
  assign n70 = ~n56 & n69 ;
  assign n71 = n70 ^ n56 ;
  assign n72 = n23 & ~n71 ;
  assign n73 = ~x3 & ~x9 ;
  assign n74 = x4 & x9 ;
  assign n75 = ~n73 & ~n74 ;
  assign n76 = ~x4 & ~x9 ;
  assign n77 = x6 & ~x7 ;
  assign n78 = ~x2 & n77 ;
  assign n79 = ~x1 & n78 ;
  assign n80 = ~n76 & n79 ;
  assign n81 = n75 & n80 ;
  assign n82 = ~n72 & ~n81 ;
  assign n83 = ~n55 & n82 ;
  assign n84 = x0 & ~n83 ;
  assign n85 = n18 & n47 ;
  assign n86 = ~x0 & ~x3 ;
  assign n87 = x9 & n86 ;
  assign n88 = ~x1 & ~x6 ;
  assign n89 = n32 & n88 ;
  assign n90 = n89 ^ x4 ;
  assign n91 = n90 ^ n89 ;
  assign n92 = n91 ^ n87 ;
  assign n93 = ~x2 & x7 ;
  assign n94 = x1 & ~n93 ;
  assign n95 = ~x6 & n94 ;
  assign n96 = n95 ^ n79 ;
  assign n97 = ~n79 & n96 ;
  assign n98 = n97 ^ n89 ;
  assign n99 = n98 ^ n79 ;
  assign n100 = n92 & n99 ;
  assign n101 = n100 ^ n97 ;
  assign n102 = n101 ^ n79 ;
  assign n103 = n87 & ~n102 ;
  assign n104 = n103 ^ n87 ;
  assign n105 = ~n85 & ~n104 ;
  assign n106 = ~n84 & n105 ;
  assign n107 = n106 ^ x8 ;
  assign n108 = n107 ^ n106 ;
  assign n157 = n75 & n88 ;
  assign n118 = ~x3 & x6 ;
  assign n158 = x4 & n118 ;
  assign n159 = ~n39 & n158 ;
  assign n160 = ~n157 & ~n159 ;
  assign n161 = n93 & ~n160 ;
  assign n109 = n33 & n45 ;
  assign n162 = x2 & x9 ;
  assign n163 = n11 & n162 ;
  assign n164 = ~x3 & ~n163 ;
  assign n165 = ~n109 & n164 ;
  assign n112 = x6 & ~x9 ;
  assign n166 = n93 & n112 ;
  assign n167 = ~n34 & ~n166 ;
  assign n168 = x9 ^ x4 ;
  assign n169 = x9 ^ x2 ;
  assign n170 = n169 ^ x2 ;
  assign n171 = n32 ^ x2 ;
  assign n172 = n170 & ~n171 ;
  assign n173 = n172 ^ x2 ;
  assign n174 = ~n168 & ~n173 ;
  assign n175 = ~x6 & n174 ;
  assign n176 = x3 & ~n175 ;
  assign n177 = n167 & n176 ;
  assign n178 = x1 & ~n177 ;
  assign n179 = ~n165 & n178 ;
  assign n180 = ~n161 & ~n179 ;
  assign n110 = x2 & x3 ;
  assign n111 = n109 & n110 ;
  assign n116 = x6 & x7 ;
  assign n117 = ~x6 & ~x7 ;
  assign n119 = ~x2 & x9 ;
  assign n120 = ~n118 & n119 ;
  assign n121 = ~n117 & n120 ;
  assign n122 = ~n116 & n121 ;
  assign n113 = x3 & n112 ;
  assign n114 = n113 ^ x9 ;
  assign n115 = n32 & ~n114 ;
  assign n123 = n122 ^ n115 ;
  assign n124 = n123 ^ n122 ;
  assign n125 = n44 & n117 ;
  assign n126 = n125 ^ n122 ;
  assign n127 = n126 ^ n122 ;
  assign n128 = ~n124 & ~n127 ;
  assign n129 = n128 ^ n122 ;
  assign n130 = x4 & ~n129 ;
  assign n131 = n130 ^ n122 ;
  assign n132 = ~n111 & ~n131 ;
  assign n133 = x1 & ~n132 ;
  assign n134 = x2 & ~x3 ;
  assign n135 = n33 & n134 ;
  assign n137 = n135 ^ n36 ;
  assign n136 = n135 ^ n46 ;
  assign n138 = n137 ^ n136 ;
  assign n139 = n138 ^ n137 ;
  assign n140 = n139 ^ n135 ;
  assign n141 = n138 ^ n73 ;
  assign n142 = x2 & ~n141 ;
  assign n143 = n137 ^ n135 ;
  assign n144 = ~n139 & n143 ;
  assign n145 = n144 ^ n140 ;
  assign n146 = n142 & n145 ;
  assign n147 = n146 ^ n144 ;
  assign n148 = n140 & n147 ;
  assign n149 = n148 ^ n144 ;
  assign n150 = n149 ^ n36 ;
  assign n151 = ~x7 & n150 ;
  assign n152 = ~x1 & x7 ;
  assign n153 = ~x9 & n152 ;
  assign n154 = n135 & n153 ;
  assign n155 = ~n151 & ~n154 ;
  assign n156 = ~n133 & n155 ;
  assign n181 = n180 ^ n156 ;
  assign n182 = ~x0 & n181 ;
  assign n183 = n182 ^ n180 ;
  assign n184 = n183 ^ n106 ;
  assign n185 = ~n108 & n184 ;
  assign n186 = n185 ^ n106 ;
  assign n187 = ~n43 & n186 ;
  assign n188 = n187 ^ x5 ;
  assign n189 = n188 ^ n187 ;
  assign n190 = ~x3 & x8 ;
  assign n191 = x9 ^ x6 ;
  assign n192 = x0 & x2 ;
  assign n193 = n192 ^ x9 ;
  assign n194 = n193 ^ n192 ;
  assign n195 = n192 ^ n12 ;
  assign n196 = ~n194 & n195 ;
  assign n197 = n196 ^ n192 ;
  assign n198 = n191 & n197 ;
  assign n199 = n152 & n198 ;
  assign n200 = n190 & n199 ;
  assign n206 = ~x7 & ~x8 ;
  assign n207 = x3 & n206 ;
  assign n208 = n162 & n207 ;
  assign n209 = x1 & n15 ;
  assign n210 = n86 & n209 ;
  assign n211 = n93 & n210 ;
  assign n212 = ~n208 & ~n211 ;
  assign n201 = x7 & ~x8 ;
  assign n202 = n73 & n201 ;
  assign n203 = x8 & x9 ;
  assign n204 = n14 & n203 ;
  assign n205 = ~n202 & ~n204 ;
  assign n213 = n212 ^ n205 ;
  assign n214 = n213 ^ n212 ;
  assign n215 = n212 ^ x2 ;
  assign n216 = n215 ^ n212 ;
  assign n217 = ~n214 & n216 ;
  assign n218 = n217 ^ n212 ;
  assign n219 = x0 & ~n218 ;
  assign n220 = n219 ^ n212 ;
  assign n221 = n46 & ~n220 ;
  assign n222 = ~n36 & ~n209 ;
  assign n223 = ~x8 & ~n39 ;
  assign n224 = n77 & ~n223 ;
  assign n225 = x2 & n224 ;
  assign n226 = n222 & n225 ;
  assign n227 = ~x8 & n153 ;
  assign n228 = ~x6 & n227 ;
  assign n229 = ~n226 & ~n228 ;
  assign n230 = x0 & ~n229 ;
  assign n231 = ~n134 & n230 ;
  assign n232 = x3 & n89 ;
  assign n233 = n15 & n232 ;
  assign n234 = n192 & n201 ;
  assign n235 = n112 & n234 ;
  assign n236 = ~x1 & ~n235 ;
  assign n237 = ~x3 & ~n236 ;
  assign n238 = x9 & n117 ;
  assign n239 = n12 & n238 ;
  assign n240 = n190 & n239 ;
  assign n241 = ~n237 & ~n240 ;
  assign n242 = x7 ^ x0 ;
  assign n243 = n242 ^ x9 ;
  assign n244 = x6 ^ x2 ;
  assign n252 = n244 ^ x2 ;
  assign n253 = n252 ^ x2 ;
  assign n254 = ~n252 & n253 ;
  assign n246 = x7 ^ x2 ;
  assign n245 = n244 ^ x9 ;
  assign n247 = n246 ^ n245 ;
  assign n248 = n246 ^ n244 ;
  assign n249 = n248 ^ x2 ;
  assign n250 = n247 & ~n249 ;
  assign n257 = n254 ^ n250 ;
  assign n251 = n250 ^ n243 ;
  assign n255 = n254 ^ n252 ;
  assign n256 = n251 & ~n255 ;
  assign n258 = n257 ^ n256 ;
  assign n259 = n243 & n258 ;
  assign n260 = n259 ^ n250 ;
  assign n261 = n260 ^ n254 ;
  assign n262 = n261 ^ n256 ;
  assign n263 = ~x8 & n262 ;
  assign n264 = x0 & ~x2 ;
  assign n265 = n112 & n264 ;
  assign n266 = ~n206 & n265 ;
  assign n267 = x1 & ~n266 ;
  assign n268 = ~n263 & n267 ;
  assign n269 = ~n241 & ~n268 ;
  assign n270 = ~n233 & ~n269 ;
  assign n271 = ~n231 & n270 ;
  assign n272 = n271 ^ x4 ;
  assign n273 = n272 ^ n271 ;
  assign n278 = ~x0 & n110 ;
  assign n310 = ~x9 & n206 ;
  assign n311 = n278 & n310 ;
  assign n274 = x0 & n238 ;
  assign n275 = n44 & n274 ;
  assign n279 = n278 ^ n275 ;
  assign n280 = n279 ^ n275 ;
  assign n276 = n275 ^ n116 ;
  assign n277 = n276 ^ n275 ;
  assign n281 = n280 ^ n277 ;
  assign n282 = n275 ^ x9 ;
  assign n283 = n282 ^ n275 ;
  assign n284 = n283 ^ n280 ;
  assign n285 = n280 & ~n284 ;
  assign n286 = n285 ^ n280 ;
  assign n287 = n281 & n286 ;
  assign n288 = n287 ^ n285 ;
  assign n289 = n288 ^ n275 ;
  assign n290 = n289 ^ n280 ;
  assign n291 = x8 & n290 ;
  assign n292 = n291 ^ n275 ;
  assign n312 = n311 ^ n292 ;
  assign n313 = n312 ^ n292 ;
  assign n293 = n264 ^ x9 ;
  assign n294 = n201 ^ x3 ;
  assign n295 = n294 ^ n201 ;
  assign n296 = n201 ^ x8 ;
  assign n297 = ~n295 & n296 ;
  assign n298 = n297 ^ n201 ;
  assign n299 = n298 ^ n264 ;
  assign n300 = n293 & n299 ;
  assign n301 = n300 ^ n297 ;
  assign n302 = n301 ^ n201 ;
  assign n303 = n302 ^ x9 ;
  assign n304 = n264 & n303 ;
  assign n305 = n304 ^ n264 ;
  assign n306 = n212 & ~n305 ;
  assign n307 = ~x6 & ~n306 ;
  assign n308 = n307 ^ n292 ;
  assign n309 = n308 ^ n292 ;
  assign n314 = n313 ^ n309 ;
  assign n317 = x7 & x9 ;
  assign n318 = x8 & n317 ;
  assign n315 = n119 & n207 ;
  assign n316 = ~n264 & ~n315 ;
  assign n319 = n318 ^ n316 ;
  assign n320 = n316 ^ n278 ;
  assign n321 = n320 ^ n278 ;
  assign n322 = x3 & n310 ;
  assign n323 = x0 & ~n322 ;
  assign n324 = n323 ^ n278 ;
  assign n325 = ~n321 & n324 ;
  assign n326 = n325 ^ n278 ;
  assign n327 = ~n319 & ~n326 ;
  assign n328 = n327 ^ n318 ;
  assign n329 = x6 & n328 ;
  assign n330 = n329 ^ n292 ;
  assign n331 = n330 ^ n292 ;
  assign n332 = n331 ^ n313 ;
  assign n333 = ~n313 & n332 ;
  assign n334 = n333 ^ n313 ;
  assign n335 = n314 & ~n334 ;
  assign n336 = n335 ^ n333 ;
  assign n337 = n336 ^ n292 ;
  assign n338 = n337 ^ n313 ;
  assign n339 = x1 & n338 ;
  assign n340 = n339 ^ n292 ;
  assign n341 = n340 ^ n271 ;
  assign n342 = n273 & ~n341 ;
  assign n343 = n342 ^ n271 ;
  assign n344 = ~n221 & n343 ;
  assign n345 = ~n200 & n344 ;
  assign n346 = n345 ^ n187 ;
  assign n347 = n189 & n346 ;
  assign n348 = n347 ^ n187 ;
  assign n349 = ~n31 & n348 ;
  assign y0 = ~n349 ;
endmodule
