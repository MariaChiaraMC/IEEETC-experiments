module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 ;
  assign n13 = ~x5 & ~x9 ;
  assign n14 = ~x3 & ~x11 ;
  assign n15 = n13 & n14 ;
  assign n16 = ~x2 & ~x10 ;
  assign n17 = x1 & x4 ;
  assign n18 = n16 & n17 ;
  assign n19 = n15 & n18 ;
  assign n20 = ~x7 & ~n19 ;
  assign n21 = ~x0 & ~n20 ;
  assign n22 = x10 & x11 ;
  assign n23 = x9 & n22 ;
  assign n24 = x7 & ~n23 ;
  assign n25 = x8 & ~n24 ;
  assign n26 = ~x6 & ~n25 ;
  assign n27 = n21 & n26 ;
  assign y0 = n27 ;
endmodule
