module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 ;
  assign n9 = ~x2 & ~x6 ;
  assign n10 = n9 ^ x4 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = n11 ^ x5 ;
  assign n13 = x1 & ~x7 ;
  assign n14 = n13 ^ x6 ;
  assign n15 = x6 & n14 ;
  assign n16 = n15 ^ n9 ;
  assign n17 = n16 ^ x6 ;
  assign n18 = n12 & n17 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n19 ^ x6 ;
  assign n21 = x5 & n20 ;
  assign n37 = x5 & x7 ;
  assign n38 = x1 & ~n37 ;
  assign n39 = x4 & ~n38 ;
  assign n40 = ~x2 & ~n39 ;
  assign n43 = x2 & x4 ;
  assign n44 = n43 ^ x4 ;
  assign n45 = n44 ^ x6 ;
  assign n41 = ~x5 & x7 ;
  assign n46 = n45 ^ n41 ;
  assign n50 = n46 ^ n44 ;
  assign n51 = n44 & n50 ;
  assign n42 = n41 ^ n13 ;
  assign n47 = n46 ^ n13 ;
  assign n48 = n47 ^ n44 ;
  assign n49 = ~n42 & ~n48 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = n46 ^ n43 ;
  assign n54 = n53 ^ n13 ;
  assign n55 = n54 ^ n48 ;
  assign n56 = n49 & n55 ;
  assign n57 = n56 ^ n49 ;
  assign n58 = n52 & n57 ;
  assign n59 = n58 ^ n51 ;
  assign n60 = n59 ^ x4 ;
  assign n61 = n60 ^ n50 ;
  assign n62 = ~n40 & n61 ;
  assign n22 = x5 & n9 ;
  assign n23 = x7 & n22 ;
  assign n24 = ~x4 & x6 ;
  assign n25 = x7 ^ x5 ;
  assign n26 = n24 & ~n25 ;
  assign n27 = ~x5 & ~x6 ;
  assign n28 = x4 & n27 ;
  assign n29 = n28 ^ x2 ;
  assign n30 = n29 ^ x2 ;
  assign n31 = x7 ^ x2 ;
  assign n32 = n30 & ~n31 ;
  assign n33 = n32 ^ x2 ;
  assign n34 = x1 & n33 ;
  assign n35 = ~n26 & ~n34 ;
  assign n36 = ~n23 & n35 ;
  assign n63 = n62 ^ n36 ;
  assign n64 = x3 & n63 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = ~n21 & n65 ;
  assign n67 = ~x0 & ~n66 ;
  assign n68 = x6 ^ x2 ;
  assign n69 = x7 ^ x6 ;
  assign n70 = ~n68 & ~n69 ;
  assign n71 = x5 & n70 ;
  assign n72 = x3 & n71 ;
  assign n73 = x0 & ~n72 ;
  assign n74 = ~x0 & ~n27 ;
  assign n75 = ~x4 & ~n74 ;
  assign n76 = ~n23 & ~n75 ;
  assign n77 = ~x5 & x6 ;
  assign n78 = ~n43 & ~n77 ;
  assign n79 = n78 ^ x2 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = n78 ^ x0 ;
  assign n82 = n81 ^ n78 ;
  assign n83 = ~n80 & ~n82 ;
  assign n84 = n83 ^ n78 ;
  assign n85 = x3 & ~n84 ;
  assign n86 = n85 ^ n78 ;
  assign n87 = n76 & n86 ;
  assign n88 = ~n73 & n87 ;
  assign n89 = ~x1 & ~n88 ;
  assign n90 = ~x3 & n22 ;
  assign n91 = ~x4 & n90 ;
  assign n92 = ~n89 & ~n91 ;
  assign n93 = ~n67 & n92 ;
  assign y0 = ~n93 ;
endmodule
