module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n15 = ~x5 & ~x10 ;
  assign n16 = x2 & x6 ;
  assign n17 = x0 & n16 ;
  assign n18 = n15 & n17 ;
  assign n19 = x11 ^ x9 ;
  assign n24 = n19 ^ x9 ;
  assign n21 = x13 ^ x9 ;
  assign n20 = n19 ^ x12 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n22 ^ x9 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n20 ^ n19 ;
  assign n27 = n26 ^ x9 ;
  assign n28 = n27 ^ x9 ;
  assign n29 = n22 & ~n28 ;
  assign n30 = n29 ^ n22 ;
  assign n31 = ~n27 & n30 ;
  assign n32 = n31 ^ x9 ;
  assign n33 = n25 & n32 ;
  assign n34 = n33 ^ n29 ;
  assign n35 = n34 ^ x9 ;
  assign n36 = n35 ^ n24 ;
  assign n37 = n18 & n36 ;
  assign y0 = n37 ;
endmodule
