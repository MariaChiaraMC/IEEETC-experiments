// Benchmark "./m1.pla" written by ABC on Thu Apr 23 10:59:54 2020

module \./m1.pla  ( 
    x0, x1, x2, x3, x4, x5,
    z4  );
  input  x0, x1, x2, x3, x4, x5;
  output z4;
  wire new_n8_, new_n9_, new_n10_, new_n11_, new_n12_, new_n13_, new_n14_;
  assign new_n8_ = ~x2 & x4;
  assign new_n9_ = x3 & x5;
  assign new_n10_ = new_n8_ & ~new_n9_;
  assign new_n11_ = ~x1 & ~new_n10_;
  assign new_n12_ = x2 & ~x4;
  assign new_n13_ = x3 & ~new_n8_;
  assign new_n14_ = ~new_n12_ & new_n13_;
  assign z4 = ~new_n11_ | new_n14_;
endmodule


