module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 ;
  assign n8 = ~x3 & ~x5 ;
  assign n9 = n8 ^ x3 ;
  assign n10 = n9 ^ x0 ;
  assign n18 = n10 ^ n9 ;
  assign n11 = x4 & x6 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = n10 ^ n8 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = ~n13 & ~n16 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = n19 ^ n13 ;
  assign n21 = ~x4 & ~x5 ;
  assign n22 = ~x6 & n21 ;
  assign n23 = n22 ^ n9 ;
  assign n24 = n17 ^ n13 ;
  assign n25 = ~n23 & ~n24 ;
  assign n26 = n25 ^ n9 ;
  assign n27 = ~n20 & n26 ;
  assign n28 = n27 ^ n9 ;
  assign n29 = n28 ^ x3 ;
  assign n30 = n29 ^ n9 ;
  assign n31 = x2 & n30 ;
  assign n36 = x5 ^ x2 ;
  assign n32 = x6 ^ x4 ;
  assign n33 = n32 ^ x2 ;
  assign n34 = n33 ^ x0 ;
  assign n35 = n34 ^ x6 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = n37 ^ x6 ;
  assign n39 = n38 ^ x3 ;
  assign n46 = n39 ^ x6 ;
  assign n53 = n46 ^ x3 ;
  assign n42 = n36 ^ x2 ;
  assign n43 = n42 ^ n36 ;
  assign n44 = n43 ^ x3 ;
  assign n54 = n44 ^ n35 ;
  assign n55 = n54 ^ n46 ;
  assign n56 = n53 & ~n55 ;
  assign n48 = n44 ^ x0 ;
  assign n49 = n48 ^ n36 ;
  assign n50 = n49 ^ x3 ;
  assign n40 = n39 ^ n35 ;
  assign n41 = n40 ^ x3 ;
  assign n45 = n44 ^ n41 ;
  assign n47 = n46 ^ n45 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = x3 & ~n51 ;
  assign n57 = n56 ^ n52 ;
  assign n58 = n57 ^ n35 ;
  assign n59 = n58 ^ n39 ;
  assign n60 = n59 ^ n44 ;
  assign n61 = n52 ^ n39 ;
  assign n62 = n61 ^ n50 ;
  assign n63 = n44 ^ x3 ;
  assign n64 = n63 ^ n50 ;
  assign n65 = n55 ^ n50 ;
  assign n66 = ~n64 & ~n65 ;
  assign n67 = n66 ^ x3 ;
  assign n68 = n67 ^ n46 ;
  assign n69 = n62 & n68 ;
  assign n70 = n69 ^ x3 ;
  assign n71 = n70 ^ n44 ;
  assign n72 = ~n60 & ~n71 ;
  assign n73 = n72 ^ n52 ;
  assign n74 = n73 ^ n66 ;
  assign n75 = n74 ^ n56 ;
  assign n76 = n75 ^ n35 ;
  assign n77 = n76 ^ n39 ;
  assign n78 = n77 ^ x3 ;
  assign n79 = n78 ^ n50 ;
  assign n80 = n79 ^ x3 ;
  assign n81 = ~n31 & n80 ;
  assign n82 = ~x1 & ~n81 ;
  assign n83 = ~x2 & x3 ;
  assign n84 = x0 & x4 ;
  assign n85 = ~n21 & ~n84 ;
  assign n86 = n83 & ~n85 ;
  assign n95 = x0 & ~x3 ;
  assign n96 = ~n84 & ~n95 ;
  assign n87 = ~x4 & x6 ;
  assign n88 = n87 ^ x6 ;
  assign n89 = x6 ^ x3 ;
  assign n90 = n89 ^ x6 ;
  assign n91 = ~n88 & ~n90 ;
  assign n92 = n91 ^ x6 ;
  assign n93 = ~n8 & ~n92 ;
  assign n97 = n96 ^ n93 ;
  assign n94 = n93 ^ x0 ;
  assign n98 = n97 ^ n94 ;
  assign n99 = n98 ^ x2 ;
  assign n100 = x3 & x5 ;
  assign n101 = ~n8 & ~n100 ;
  assign n102 = n101 ^ n94 ;
  assign n103 = n102 ^ n96 ;
  assign n104 = n96 & ~n103 ;
  assign n105 = n104 ^ n94 ;
  assign n106 = n105 ^ n96 ;
  assign n107 = n99 & n106 ;
  assign n108 = n107 ^ n104 ;
  assign n109 = n108 ^ n96 ;
  assign n110 = x2 & n109 ;
  assign n111 = n110 ^ n93 ;
  assign n112 = ~n86 & ~n111 ;
  assign n113 = x1 & ~n112 ;
  assign n114 = n93 & ~n96 ;
  assign n115 = ~x0 & x6 ;
  assign n116 = n100 & n115 ;
  assign n117 = ~x4 & n116 ;
  assign n118 = ~n114 & ~n117 ;
  assign n119 = n118 ^ x2 ;
  assign n120 = n119 ^ n118 ;
  assign n121 = n120 ^ n113 ;
  assign n122 = ~x0 & ~x1 ;
  assign n123 = ~x3 & ~n122 ;
  assign n124 = n123 ^ n11 ;
  assign n125 = n11 & n124 ;
  assign n126 = n125 ^ n118 ;
  assign n127 = n126 ^ n11 ;
  assign n128 = ~n121 & ~n127 ;
  assign n129 = n128 ^ n125 ;
  assign n130 = n129 ^ n11 ;
  assign n131 = ~n113 & n130 ;
  assign n132 = n131 ^ n113 ;
  assign n133 = ~n82 & ~n132 ;
  assign y0 = ~n133 ;
endmodule
