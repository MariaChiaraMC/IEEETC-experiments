module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 ;
  assign n9 = x0 & x1 ;
  assign n10 = ~x2 & ~x3 ;
  assign n11 = n9 & n10 ;
  assign n12 = x2 & x3 ;
  assign n13 = ~n10 & ~n12 ;
  assign n14 = ~x0 & ~x1 ;
  assign n15 = ~n9 & ~n14 ;
  assign n16 = n13 & n15 ;
  assign n17 = ~n11 & ~n16 ;
  assign n18 = x4 & x5 ;
  assign n19 = ~x4 & ~x5 ;
  assign n20 = x6 & x7 ;
  assign n21 = n19 & n20 ;
  assign n22 = ~n18 & ~n21 ;
  assign n23 = ~n17 & ~n22 ;
  assign n24 = x7 ^ x6 ;
  assign n25 = n14 ^ x7 ;
  assign n26 = n24 & ~n25 ;
  assign n27 = n26 ^ x7 ;
  assign n28 = ~n9 & n27 ;
  assign n29 = n28 ^ n12 ;
  assign n30 = n10 & n18 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = ~n9 & ~n18 ;
  assign n35 = ~n14 & ~n19 ;
  assign n36 = n34 & ~n35 ;
  assign n37 = n36 ^ n31 ;
  assign n38 = n37 ^ n29 ;
  assign n39 = n33 & n38 ;
  assign n40 = n39 ^ n36 ;
  assign n41 = ~n19 & n36 ;
  assign n42 = n41 ^ n29 ;
  assign n43 = n40 & ~n42 ;
  assign n44 = n43 ^ n41 ;
  assign n45 = ~n29 & n44 ;
  assign n46 = n45 ^ n39 ;
  assign n47 = n46 ^ n12 ;
  assign n48 = n47 ^ n36 ;
  assign n49 = ~n23 & ~n48 ;
  assign n50 = ~x6 & ~x7 ;
  assign n51 = ~n35 & ~n50 ;
  assign n52 = n51 ^ n9 ;
  assign n53 = n52 ^ n13 ;
  assign n54 = n19 ^ n18 ;
  assign n55 = n9 & n54 ;
  assign n56 = n55 ^ n18 ;
  assign n57 = n53 & n56 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = n58 ^ n18 ;
  assign n60 = n59 ^ n9 ;
  assign n61 = n13 & n60 ;
  assign n62 = n49 & ~n61 ;
  assign n63 = x5 ^ x4 ;
  assign n64 = n12 & n14 ;
  assign n65 = ~n11 & ~n64 ;
  assign n66 = ~n50 & ~n65 ;
  assign n67 = n28 ^ x3 ;
  assign n68 = n67 ^ x2 ;
  assign n69 = n68 ^ n28 ;
  assign n70 = n69 ^ n66 ;
  assign n71 = n15 & n20 ;
  assign n72 = n71 ^ x2 ;
  assign n73 = n71 & ~n72 ;
  assign n74 = n73 ^ n28 ;
  assign n75 = n74 ^ n71 ;
  assign n76 = n70 & n75 ;
  assign n77 = n76 ^ n73 ;
  assign n78 = n77 ^ n71 ;
  assign n79 = ~n66 & n78 ;
  assign n80 = n79 ^ n66 ;
  assign n81 = n63 & n80 ;
  assign n82 = n62 & ~n81 ;
  assign y0 = ~n82 ;
endmodule
