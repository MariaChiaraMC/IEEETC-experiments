module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 ;
  assign n20 = x18 ^ x15 ;
  assign n21 = n20 ^ x18 ;
  assign n22 = ~x10 & x15 ;
  assign n23 = ~x6 & ~x7 ;
  assign n24 = x8 & x9 ;
  assign n25 = n23 & ~n24 ;
  assign n26 = n22 & n25 ;
  assign n27 = ~x2 & n26 ;
  assign n28 = x18 & ~n27 ;
  assign n29 = x4 & n25 ;
  assign n30 = ~x15 & ~n29 ;
  assign n31 = ~x3 & n30 ;
  assign n32 = n28 & ~n31 ;
  assign n33 = n32 ^ x14 ;
  assign n34 = n33 ^ x18 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = n35 ^ n21 ;
  assign n37 = n21 & n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = n33 ^ n32 ;
  assign n50 = ~x8 & n23 ;
  assign n48 = ~n32 & n39 ;
  assign n40 = x1 & ~x11 ;
  assign n41 = ~x12 & n40 ;
  assign n42 = x3 & ~x10 ;
  assign n43 = ~x5 & n42 ;
  assign n44 = n41 & ~n43 ;
  assign n45 = n35 ^ n32 ;
  assign n46 = n45 ^ n21 ;
  assign n47 = n44 & ~n46 ;
  assign n49 = n48 ^ n47 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = n51 ^ n32 ;
  assign n53 = n39 & n52 ;
  assign n54 = n53 ^ n47 ;
  assign n55 = n38 & n54 ;
  assign n56 = n55 ^ n47 ;
  assign n57 = n56 ^ n48 ;
  assign n58 = n57 ^ n53 ;
  assign n59 = n58 ^ n32 ;
  assign n60 = n59 ^ x14 ;
  assign y0 = n60 ;
endmodule
