module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 ;
  output y0 ;
  wire n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 ;
  assign n24 = ~x0 & x1 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = n25 ^ x2 ;
  assign n27 = n26 ^ n25 ;
  assign n31 = n25 ^ x3 ;
  assign n32 = n25 & n31 ;
  assign n28 = x0 & ~x1 ;
  assign n29 = x5 & ~n28 ;
  assign n35 = n32 ^ n29 ;
  assign n30 = n29 ^ n27 ;
  assign n33 = n32 ^ n25 ;
  assign n34 = n30 & n33 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = n27 & n36 ;
  assign n38 = n37 ^ n32 ;
  assign n39 = n38 ^ n34 ;
  assign n40 = n39 ^ x5 ;
  assign n41 = ~x4 & n40 ;
  assign n42 = ~x19 & ~x20 ;
  assign n43 = n42 ^ x18 ;
  assign n44 = n43 ^ x18 ;
  assign n45 = ~x1 & x5 ;
  assign n46 = ~x8 & ~x11 ;
  assign n47 = x10 & n46 ;
  assign n48 = ~x9 & n47 ;
  assign n49 = ~x6 & ~x7 ;
  assign n50 = ~x12 & ~x13 ;
  assign n51 = ~x4 & n50 ;
  assign n52 = n49 & n51 ;
  assign n53 = n28 & n52 ;
  assign n54 = n48 & n53 ;
  assign n55 = ~n45 & ~n54 ;
  assign n56 = x11 & ~x12 ;
  assign n57 = ~x8 & x9 ;
  assign n58 = n56 & n57 ;
  assign n59 = ~x0 & ~n58 ;
  assign n60 = x15 & ~n59 ;
  assign n61 = ~x0 & ~x2 ;
  assign n63 = x9 & x10 ;
  assign n64 = ~n57 & ~n63 ;
  assign n62 = x13 ^ x12 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = n65 ^ x13 ;
  assign n72 = n66 ^ n62 ;
  assign n73 = n72 ^ x13 ;
  assign n74 = n73 ^ x13 ;
  assign n75 = n62 ^ x11 ;
  assign n76 = n75 ^ n62 ;
  assign n77 = n76 ^ x13 ;
  assign n78 = ~n74 & n77 ;
  assign n67 = ~x10 & ~x11 ;
  assign n68 = n67 ^ n62 ;
  assign n69 = n68 ^ n66 ;
  assign n70 = n69 ^ x13 ;
  assign n71 = n66 & ~n70 ;
  assign n79 = n78 ^ n71 ;
  assign n80 = n79 ^ n66 ;
  assign n81 = n71 ^ x13 ;
  assign n82 = n81 ^ n73 ;
  assign n83 = x13 & ~n82 ;
  assign n84 = n83 ^ n71 ;
  assign n85 = n80 & n84 ;
  assign n86 = n85 ^ n78 ;
  assign n87 = n86 ^ n83 ;
  assign n88 = n87 ^ n66 ;
  assign n89 = n88 ^ x13 ;
  assign n90 = n89 ^ n73 ;
  assign n91 = n90 ^ x12 ;
  assign n92 = n61 & n91 ;
  assign n93 = ~n60 & ~n92 ;
  assign n94 = ~n55 & ~n93 ;
  assign n95 = n56 & n63 ;
  assign n96 = x1 & x13 ;
  assign n97 = ~n95 & ~n96 ;
  assign n98 = ~x2 & x15 ;
  assign n99 = ~n97 & n98 ;
  assign n100 = x4 & ~n99 ;
  assign n101 = ~n94 & n100 ;
  assign n102 = x5 & ~n101 ;
  assign n103 = n24 & n52 ;
  assign n104 = ~x10 & x11 ;
  assign n105 = x15 & n104 ;
  assign n106 = x8 & x9 ;
  assign n107 = n105 & n106 ;
  assign n108 = ~n48 & ~n107 ;
  assign n109 = n103 & ~n108 ;
  assign n110 = x5 & x15 ;
  assign n111 = x1 & n110 ;
  assign n112 = x4 & ~n111 ;
  assign n113 = n61 & ~n112 ;
  assign n114 = x15 & n47 ;
  assign n115 = n103 & n114 ;
  assign n116 = ~x1 & x2 ;
  assign n117 = x5 & n116 ;
  assign n118 = ~n115 & ~n117 ;
  assign n119 = x17 & ~n118 ;
  assign n120 = ~n113 & ~n119 ;
  assign n121 = ~n109 & n120 ;
  assign n122 = ~x0 & ~x15 ;
  assign n123 = x12 ^ x6 ;
  assign n124 = ~x13 & n123 ;
  assign n125 = n124 ^ x6 ;
  assign n126 = n122 & ~n125 ;
  assign n127 = x8 & ~x10 ;
  assign n128 = ~x12 & ~n127 ;
  assign n129 = x16 & n49 ;
  assign n130 = ~n128 & n129 ;
  assign n131 = ~x13 & ~n130 ;
  assign n132 = ~x0 & n131 ;
  assign n133 = ~n126 & ~n132 ;
  assign n134 = x15 & n63 ;
  assign n138 = x9 & ~n67 ;
  assign n135 = ~x9 & n104 ;
  assign n136 = ~x8 & n135 ;
  assign n137 = x16 & n136 ;
  assign n139 = n138 ^ n137 ;
  assign n140 = n139 ^ x13 ;
  assign n148 = n140 ^ n139 ;
  assign n141 = x6 & ~n46 ;
  assign n142 = n141 ^ n140 ;
  assign n143 = n142 ^ n139 ;
  assign n144 = n140 ^ n137 ;
  assign n145 = n144 ^ n141 ;
  assign n146 = n145 ^ n143 ;
  assign n147 = ~n143 & ~n146 ;
  assign n149 = n148 ^ n147 ;
  assign n150 = n149 ^ n143 ;
  assign n151 = n139 ^ n127 ;
  assign n152 = n147 ^ n143 ;
  assign n153 = ~n151 & ~n152 ;
  assign n154 = n153 ^ n139 ;
  assign n155 = ~n150 & n154 ;
  assign n156 = n155 ^ n139 ;
  assign n157 = n156 ^ n138 ;
  assign n158 = n157 ^ n139 ;
  assign n159 = n158 ^ x7 ;
  assign n160 = n159 ^ n158 ;
  assign n161 = n160 ^ n134 ;
  assign n162 = x15 ^ x8 ;
  assign n163 = n162 ^ x16 ;
  assign n164 = ~x11 & ~x13 ;
  assign n165 = ~x9 & x10 ;
  assign n166 = n164 & n165 ;
  assign n167 = n166 ^ n104 ;
  assign n168 = x15 & ~n167 ;
  assign n169 = n168 ^ n166 ;
  assign n170 = ~n163 & n169 ;
  assign n171 = n170 ^ n168 ;
  assign n172 = n171 ^ n166 ;
  assign n173 = n172 ^ x15 ;
  assign n174 = ~x16 & n173 ;
  assign n175 = ~n114 & ~n174 ;
  assign n176 = n175 ^ x6 ;
  assign n177 = ~n175 & n176 ;
  assign n178 = n177 ^ n158 ;
  assign n179 = n178 ^ n175 ;
  assign n180 = n161 & ~n179 ;
  assign n181 = n180 ^ n177 ;
  assign n182 = n181 ^ n175 ;
  assign n183 = ~n134 & ~n182 ;
  assign n184 = n183 ^ n134 ;
  assign n185 = ~x12 & n184 ;
  assign n186 = ~n133 & ~n185 ;
  assign n187 = x2 & ~n55 ;
  assign n188 = ~n186 & n187 ;
  assign n189 = n121 & ~n188 ;
  assign n190 = ~n102 & n189 ;
  assign n191 = ~x3 & ~n190 ;
  assign n192 = ~x1 & ~x2 ;
  assign n193 = x15 ^ x0 ;
  assign n194 = n193 ^ x15 ;
  assign n195 = x21 ^ x15 ;
  assign n196 = n194 & ~n195 ;
  assign n197 = n196 ^ x15 ;
  assign n198 = x3 & n197 ;
  assign n199 = x4 & ~n198 ;
  assign n200 = n192 & ~n199 ;
  assign n201 = x1 & x3 ;
  assign n202 = x2 & n201 ;
  assign n203 = ~n52 & ~n202 ;
  assign n204 = n46 & n63 ;
  assign n205 = ~n201 & ~n204 ;
  assign n206 = n205 ^ x15 ;
  assign n207 = n206 ^ n205 ;
  assign n208 = n205 ^ n136 ;
  assign n209 = n208 ^ n205 ;
  assign n210 = n207 & n209 ;
  assign n211 = n210 ^ n205 ;
  assign n212 = ~x2 & ~n211 ;
  assign n213 = n212 ^ n205 ;
  assign n214 = ~n203 & ~n213 ;
  assign n215 = ~n200 & ~n214 ;
  assign n216 = x5 & ~n215 ;
  assign n217 = x22 & n202 ;
  assign n218 = ~x3 & ~n192 ;
  assign n219 = x1 ^ x0 ;
  assign n220 = ~n218 & n219 ;
  assign n221 = ~x5 & n220 ;
  assign n222 = ~n217 & ~n221 ;
  assign n223 = x4 & ~n222 ;
  assign n224 = x3 & ~x5 ;
  assign n225 = n106 & n224 ;
  assign n226 = ~x0 & n225 ;
  assign n227 = n116 & n226 ;
  assign n228 = n52 & n227 ;
  assign n229 = n104 & n228 ;
  assign n230 = ~n223 & ~n229 ;
  assign n231 = ~n216 & n230 ;
  assign n232 = ~n191 & n231 ;
  assign n233 = n232 ^ x18 ;
  assign n234 = n44 & n233 ;
  assign n235 = n234 ^ x18 ;
  assign n236 = x14 & n235 ;
  assign n237 = ~n41 & n236 ;
  assign y0 = ~n237 ;
endmodule
