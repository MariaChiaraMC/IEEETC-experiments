module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 ;
  assign n20 = ~x7 & x16 ;
  assign n21 = n20 ^ x9 ;
  assign n22 = n21 ^ x9 ;
  assign n23 = x17 ^ x9 ;
  assign n24 = n23 ^ x9 ;
  assign n25 = n22 & ~n24 ;
  assign n26 = n25 ^ x9 ;
  assign n27 = ~x18 & n26 ;
  assign n28 = n27 ^ x9 ;
  assign n29 = x8 & n28 ;
  assign n30 = ~x17 & ~x18 ;
  assign n31 = x6 & x16 ;
  assign n32 = n30 & ~n31 ;
  assign n33 = x8 & ~x18 ;
  assign n34 = x17 & ~n33 ;
  assign n35 = x7 & ~n34 ;
  assign n36 = ~n32 & n35 ;
  assign n37 = ~n29 & ~n36 ;
  assign n38 = x16 ^ x6 ;
  assign n39 = ~n30 & n38 ;
  assign n40 = x9 & ~x18 ;
  assign n41 = x7 & ~n40 ;
  assign n42 = n34 & ~n41 ;
  assign n43 = x15 & ~n42 ;
  assign n44 = ~n39 & n43 ;
  assign n45 = n37 & n44 ;
  assign n46 = ~x2 & ~x10 ;
  assign n47 = n46 ^ x16 ;
  assign n48 = n46 ^ n30 ;
  assign n49 = n48 ^ n30 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = x6 & ~n40 ;
  assign n52 = n51 ^ x8 ;
  assign n53 = ~x8 & n52 ;
  assign n54 = n53 ^ n30 ;
  assign n55 = n54 ^ x8 ;
  assign n56 = ~n50 & ~n55 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n57 ^ x8 ;
  assign n59 = ~n47 & ~n58 ;
  assign n60 = n59 ^ n46 ;
  assign n61 = n45 & n60 ;
  assign n62 = x7 & ~x17 ;
  assign n63 = ~x6 & x16 ;
  assign n64 = n33 & n63 ;
  assign n65 = n62 & n64 ;
  assign n66 = ~x7 & x17 ;
  assign n67 = n66 ^ x18 ;
  assign n68 = n67 ^ n38 ;
  assign n69 = ~n62 & ~n68 ;
  assign n70 = n69 ^ n62 ;
  assign n71 = n66 ^ x8 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = n67 & ~n72 ;
  assign n74 = n73 ^ n67 ;
  assign n75 = n74 ^ n38 ;
  assign n76 = ~n70 & ~n75 ;
  assign n77 = ~n65 & ~n76 ;
  assign n78 = x4 & ~x9 ;
  assign n79 = ~n77 & n78 ;
  assign n80 = ~x16 & n30 ;
  assign n81 = n80 ^ x3 ;
  assign n82 = n81 ^ x3 ;
  assign n83 = n82 ^ x15 ;
  assign n84 = x3 & ~x5 ;
  assign n85 = ~x10 & n84 ;
  assign n86 = x12 & x13 ;
  assign n87 = x11 & n86 ;
  assign n88 = ~n85 & ~n87 ;
  assign n89 = n88 ^ x1 ;
  assign n90 = x1 & n89 ;
  assign n91 = n90 ^ x3 ;
  assign n92 = n91 ^ x1 ;
  assign n93 = ~n83 & n92 ;
  assign n94 = n93 ^ n90 ;
  assign n95 = n94 ^ x1 ;
  assign n96 = ~x15 & n95 ;
  assign n97 = n96 ^ x15 ;
  assign n98 = ~n79 & ~n97 ;
  assign n99 = ~x0 & ~x14 ;
  assign n100 = ~n98 & n99 ;
  assign n101 = ~n61 & n100 ;
  assign y0 = n101 ;
endmodule
