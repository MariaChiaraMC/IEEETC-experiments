module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 ;
  assign n8 = ~x0 & ~x4 ;
  assign n9 = x3 & n8 ;
  assign n10 = x6 ^ x5 ;
  assign n11 = n10 ^ x1 ;
  assign n12 = n11 ^ x2 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = x6 ^ x1 ;
  assign n15 = n14 ^ x1 ;
  assign n16 = ~x2 & n15 ;
  assign n17 = n16 ^ x1 ;
  assign n18 = ~n13 & ~n17 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n19 ^ x1 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = n9 & n21 ;
  assign y0 = n22 ;
endmodule
