module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n13 = x10 & x11 ;
  assign n14 = ~x9 & n13 ;
  assign n15 = x6 & ~n14 ;
  assign n16 = x7 & ~x8 ;
  assign n17 = x6 & ~n16 ;
  assign n18 = x4 & n17 ;
  assign n19 = ~n15 & ~n18 ;
  assign n20 = x7 & ~x11 ;
  assign n21 = n20 ^ x5 ;
  assign n22 = ~x0 & ~n21 ;
  assign n23 = n19 & n22 ;
  assign n24 = x6 ^ x4 ;
  assign n25 = n16 ^ x6 ;
  assign n26 = n25 ^ n16 ;
  assign n27 = x9 & ~n13 ;
  assign n28 = n27 ^ n16 ;
  assign n29 = ~n26 & n28 ;
  assign n30 = n29 ^ n16 ;
  assign n31 = n24 & ~n30 ;
  assign n32 = n31 ^ x4 ;
  assign n33 = n23 & n32 ;
  assign y0 = n33 ;
endmodule
