module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 ;
  assign n13 = x2 & x4 ;
  assign n14 = x5 & n13 ;
  assign n15 = ~x4 & x11 ;
  assign n16 = n15 ^ x3 ;
  assign n17 = n16 ^ x3 ;
  assign n18 = x10 ^ x3 ;
  assign n19 = n18 ^ x3 ;
  assign n20 = ~n17 & n19 ;
  assign n21 = n20 ^ x3 ;
  assign n22 = ~x2 & ~n21 ;
  assign n23 = n22 ^ x3 ;
  assign n24 = ~n14 & n23 ;
  assign n25 = x8 & ~n24 ;
  assign n26 = x11 ^ x10 ;
  assign n27 = x11 ^ x5 ;
  assign n28 = n27 ^ x5 ;
  assign n29 = x5 ^ x2 ;
  assign n30 = n28 & n29 ;
  assign n31 = n30 ^ x5 ;
  assign n32 = ~n26 & n31 ;
  assign n33 = n32 ^ x10 ;
  assign n34 = ~n25 & n33 ;
  assign n35 = x7 ^ x4 ;
  assign n45 = n35 ^ x3 ;
  assign n37 = n35 ^ x8 ;
  assign n46 = n45 ^ n37 ;
  assign n38 = n37 ^ x7 ;
  assign n47 = n46 ^ n38 ;
  assign n48 = n47 ^ n38 ;
  assign n49 = n48 ^ n37 ;
  assign n50 = n49 ^ n35 ;
  assign n52 = n50 ^ n35 ;
  assign n55 = n52 ^ n50 ;
  assign n56 = n47 ^ x2 ;
  assign n57 = n56 ^ x5 ;
  assign n36 = n35 ^ x5 ;
  assign n58 = n57 ^ n36 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n39 ^ n35 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n41 ^ n35 ;
  assign n43 = n42 ^ n36 ;
  assign n59 = n58 ^ n43 ;
  assign n60 = n59 ^ n50 ;
  assign n61 = ~n55 & ~n60 ;
  assign n44 = n43 ^ n40 ;
  assign n51 = n50 ^ n40 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = ~n44 & ~n53 ;
  assign n62 = n61 ^ n54 ;
  assign n63 = n62 ^ n57 ;
  assign n64 = n63 ^ n40 ;
  assign n65 = n64 ^ n50 ;
  assign n66 = n40 ^ n36 ;
  assign n67 = n66 ^ n43 ;
  assign n68 = n67 ^ n52 ;
  assign n69 = n67 ^ n50 ;
  assign n70 = n69 ^ n52 ;
  assign n71 = n68 & n70 ;
  assign n72 = n71 ^ n54 ;
  assign n73 = n72 ^ n36 ;
  assign n74 = n73 ^ n40 ;
  assign n75 = ~n52 & n74 ;
  assign n76 = n75 ^ n50 ;
  assign n77 = n65 & n76 ;
  assign n78 = n77 ^ n54 ;
  assign n79 = n78 ^ n40 ;
  assign n80 = n79 ^ n50 ;
  assign n81 = n80 ^ n52 ;
  assign n82 = n81 ^ x4 ;
  assign n83 = n82 ^ n42 ;
  assign n84 = x9 ^ x8 ;
  assign n85 = n84 ^ x9 ;
  assign n86 = x7 & ~n13 ;
  assign n87 = x5 & ~x11 ;
  assign n88 = ~x3 & x4 ;
  assign n89 = n87 & ~n88 ;
  assign n90 = ~n86 & n89 ;
  assign n91 = n90 ^ x9 ;
  assign n92 = ~n85 & n91 ;
  assign n93 = n92 ^ x9 ;
  assign n94 = ~x7 & ~x9 ;
  assign n95 = n94 ^ n83 ;
  assign n96 = ~n93 & ~n95 ;
  assign n97 = n96 ^ n94 ;
  assign n98 = ~n83 & n97 ;
  assign n99 = n98 ^ n83 ;
  assign n100 = n34 & ~n99 ;
  assign y0 = n100 ;
endmodule
