module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 ;
  output y0 ;
  wire n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 ;
  assign n24 = x0 & ~x1 ;
  assign n25 = x2 & ~x3 ;
  assign n26 = ~x2 & x3 ;
  assign n27 = ~n25 & ~n26 ;
  assign n28 = n24 & ~n27 ;
  assign n29 = n28 ^ x5 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = n30 ^ x4 ;
  assign n32 = ~x2 & ~x3 ;
  assign n33 = ~x0 & x1 ;
  assign n34 = n33 ^ n32 ;
  assign n35 = n32 & n34 ;
  assign n36 = n35 ^ n28 ;
  assign n37 = n36 ^ n32 ;
  assign n38 = n31 & n37 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n39 ^ n32 ;
  assign n41 = ~x4 & n40 ;
  assign n300 = ~x19 & ~x20 ;
  assign n42 = x8 & ~x10 ;
  assign n43 = x9 & n42 ;
  assign n44 = x11 & n43 ;
  assign n45 = n25 & n33 ;
  assign n46 = ~x6 & ~x7 ;
  assign n47 = ~x12 & ~x13 ;
  assign n48 = n46 & n47 ;
  assign n49 = ~x15 & n48 ;
  assign n50 = n45 & n49 ;
  assign n51 = n44 & n50 ;
  assign n52 = ~x7 & ~x10 ;
  assign n53 = x8 & x10 ;
  assign n54 = ~x13 & ~n53 ;
  assign n55 = ~n52 & n54 ;
  assign n56 = x11 & ~x15 ;
  assign n57 = ~x16 & n56 ;
  assign n58 = ~x6 & n47 ;
  assign n59 = n58 ^ x13 ;
  assign n60 = n57 & n59 ;
  assign n61 = ~n55 & n60 ;
  assign n62 = x6 & x13 ;
  assign n63 = ~x17 & ~n62 ;
  assign n64 = ~x8 & ~x10 ;
  assign n65 = x11 & n64 ;
  assign n66 = x13 & ~x15 ;
  assign n67 = x9 & x10 ;
  assign n68 = ~x8 & n67 ;
  assign n69 = n66 & ~n68 ;
  assign n70 = ~n65 & n69 ;
  assign n71 = n63 & ~n70 ;
  assign n72 = x9 & n66 ;
  assign n73 = ~x6 & ~x13 ;
  assign n74 = x16 & n73 ;
  assign n75 = x7 & n74 ;
  assign n76 = ~n72 & ~n75 ;
  assign n77 = n76 ^ x12 ;
  assign n78 = n77 ^ n76 ;
  assign n81 = ~x11 & ~x13 ;
  assign n96 = n64 & n81 ;
  assign n97 = ~n56 & ~n96 ;
  assign n98 = n46 & ~n97 ;
  assign n79 = x15 ^ x10 ;
  assign n80 = n79 ^ x15 ;
  assign n82 = n81 ^ x15 ;
  assign n83 = n80 & ~n82 ;
  assign n84 = n83 ^ x15 ;
  assign n85 = x8 & ~n84 ;
  assign n86 = n46 & n85 ;
  assign n87 = x7 & x11 ;
  assign n88 = n53 ^ x13 ;
  assign n89 = n88 ^ n53 ;
  assign n90 = x16 & n64 ;
  assign n91 = n90 ^ n53 ;
  assign n92 = n89 & n91 ;
  assign n93 = n92 ^ n53 ;
  assign n94 = n87 & n93 ;
  assign n95 = ~n86 & ~n94 ;
  assign n99 = n98 ^ n95 ;
  assign n100 = n99 ^ n95 ;
  assign n101 = ~x11 & ~n53 ;
  assign n102 = ~x15 & ~n42 ;
  assign n103 = x6 & x7 ;
  assign n104 = ~n102 & ~n103 ;
  assign n105 = ~n101 & ~n104 ;
  assign n106 = n105 ^ n95 ;
  assign n107 = n106 ^ n95 ;
  assign n108 = ~n100 & ~n107 ;
  assign n109 = n108 ^ n95 ;
  assign n110 = x9 & n109 ;
  assign n111 = n110 ^ n95 ;
  assign n112 = n111 ^ n76 ;
  assign n113 = ~n78 & n112 ;
  assign n114 = n113 ^ n76 ;
  assign n115 = n71 & n114 ;
  assign n116 = ~x1 & ~n115 ;
  assign n117 = ~n61 & ~n116 ;
  assign n118 = x4 & ~n117 ;
  assign n119 = ~x1 & ~x4 ;
  assign n120 = ~x21 & n119 ;
  assign n121 = x0 & x4 ;
  assign n122 = ~x16 & n121 ;
  assign n123 = ~n120 & ~n122 ;
  assign n124 = ~n24 & n123 ;
  assign n125 = ~n118 & n124 ;
  assign n126 = n25 & ~n125 ;
  assign n127 = x4 & ~x15 ;
  assign n128 = n33 & n127 ;
  assign n129 = ~x3 & n128 ;
  assign n134 = x9 & ~x11 ;
  assign n135 = n64 & n134 ;
  assign n136 = x12 & ~n135 ;
  assign n137 = x13 & ~n136 ;
  assign n138 = x4 & ~n137 ;
  assign n130 = x11 & n67 ;
  assign n131 = ~x12 & n130 ;
  assign n132 = ~x13 & ~n131 ;
  assign n133 = n127 & ~n132 ;
  assign n139 = n138 ^ n133 ;
  assign n140 = n139 ^ x1 ;
  assign n148 = n140 ^ n139 ;
  assign n141 = ~x16 & n119 ;
  assign n142 = n141 ^ n140 ;
  assign n143 = n142 ^ n139 ;
  assign n144 = n140 ^ n133 ;
  assign n145 = n144 ^ n141 ;
  assign n146 = n145 ^ n143 ;
  assign n147 = ~n143 & n146 ;
  assign n149 = n148 ^ n147 ;
  assign n150 = n149 ^ n143 ;
  assign n151 = n139 ^ x0 ;
  assign n152 = n147 ^ n143 ;
  assign n153 = ~n151 & ~n152 ;
  assign n154 = n153 ^ n139 ;
  assign n155 = ~n150 & ~n154 ;
  assign n156 = n155 ^ n139 ;
  assign n157 = n156 ^ n138 ;
  assign n158 = n157 ^ n139 ;
  assign n159 = n32 & ~n158 ;
  assign n160 = x5 & ~n159 ;
  assign n161 = ~x4 & n33 ;
  assign n164 = n48 ^ x1 ;
  assign n165 = n164 ^ x1 ;
  assign n162 = x4 ^ x1 ;
  assign n163 = n162 ^ x1 ;
  assign n166 = n165 ^ n163 ;
  assign n167 = ~x9 & ~x10 ;
  assign n168 = x11 & n167 ;
  assign n169 = ~n134 & ~n168 ;
  assign n170 = ~x8 & ~n169 ;
  assign n171 = ~n44 & ~n170 ;
  assign n172 = n171 ^ x1 ;
  assign n173 = n172 ^ x1 ;
  assign n174 = n173 ^ n165 ;
  assign n175 = n165 & ~n174 ;
  assign n176 = n175 ^ n165 ;
  assign n177 = ~n166 & n176 ;
  assign n178 = n177 ^ n175 ;
  assign n179 = n178 ^ x1 ;
  assign n180 = n179 ^ n165 ;
  assign n181 = ~x0 & n180 ;
  assign n182 = n181 ^ x1 ;
  assign n183 = x3 & n182 ;
  assign n184 = ~n161 & ~n183 ;
  assign n185 = n184 ^ x2 ;
  assign n186 = n185 ^ n184 ;
  assign n187 = n186 ^ n160 ;
  assign n188 = x1 ^ x0 ;
  assign n189 = x13 ^ x9 ;
  assign n190 = n189 ^ n49 ;
  assign n191 = n65 ^ x4 ;
  assign n192 = ~n190 & ~n191 ;
  assign n193 = n192 ^ n190 ;
  assign n194 = n193 ^ x4 ;
  assign n196 = n65 ^ x9 ;
  assign n197 = n196 ^ n65 ;
  assign n195 = n190 ^ n49 ;
  assign n198 = n197 ^ n195 ;
  assign n199 = n65 ^ x12 ;
  assign n200 = n199 ^ n197 ;
  assign n201 = n198 & ~n200 ;
  assign n202 = n201 ^ n199 ;
  assign n203 = n202 ^ n195 ;
  assign n204 = n195 ^ x4 ;
  assign n205 = ~x4 & ~n204 ;
  assign n206 = n205 ^ n197 ;
  assign n207 = n206 ^ n199 ;
  assign n208 = n207 ^ x4 ;
  assign n209 = ~n203 & n208 ;
  assign n210 = n209 ^ n197 ;
  assign n211 = n210 ^ n65 ;
  assign n212 = n211 ^ n199 ;
  assign n213 = n194 & ~n212 ;
  assign n214 = n213 ^ n205 ;
  assign n215 = n214 ^ x4 ;
  assign n216 = n215 ^ x1 ;
  assign n217 = n216 ^ n215 ;
  assign n218 = n215 ^ n127 ;
  assign n219 = ~n217 & n218 ;
  assign n220 = n219 ^ n215 ;
  assign n221 = ~n188 & n220 ;
  assign n222 = n221 ^ x0 ;
  assign n223 = n222 ^ x3 ;
  assign n224 = n222 & n223 ;
  assign n225 = n224 ^ n184 ;
  assign n226 = n225 ^ n222 ;
  assign n227 = ~n187 & ~n226 ;
  assign n228 = n227 ^ n224 ;
  assign n229 = n228 ^ n222 ;
  assign n230 = n160 & n229 ;
  assign n231 = n230 ^ n160 ;
  assign n232 = ~n129 & n231 ;
  assign n233 = ~n126 & n232 ;
  assign n234 = x2 & x22 ;
  assign n235 = x3 & n121 ;
  assign n236 = ~n234 & n235 ;
  assign n237 = ~x4 & n47 ;
  assign n238 = x0 & x1 ;
  assign n239 = n238 ^ x1 ;
  assign n240 = n239 ^ x1 ;
  assign n241 = x2 ^ x1 ;
  assign n242 = n241 ^ x1 ;
  assign n243 = n240 & n242 ;
  assign n244 = n243 ^ x1 ;
  assign n245 = ~x3 & ~n244 ;
  assign n246 = n245 ^ x1 ;
  assign n247 = n44 & ~n246 ;
  assign n248 = ~x1 & n26 ;
  assign n249 = ~x9 & ~n248 ;
  assign n250 = ~x0 & n249 ;
  assign n251 = ~x11 & ~n250 ;
  assign n252 = ~x0 & ~x1 ;
  assign n253 = n25 & ~n252 ;
  assign n254 = ~x0 & n26 ;
  assign n255 = ~n253 & ~n254 ;
  assign n256 = ~n167 & ~n255 ;
  assign n257 = n251 & n256 ;
  assign n258 = ~x8 & n257 ;
  assign n259 = ~n247 & ~n258 ;
  assign n260 = n46 & ~n259 ;
  assign n261 = ~n248 & ~n253 ;
  assign n262 = n53 & ~n261 ;
  assign n263 = n134 & n262 ;
  assign n264 = ~n260 & ~n263 ;
  assign n265 = n237 & ~n264 ;
  assign n266 = x4 & ~n25 ;
  assign n267 = n24 & n266 ;
  assign n268 = ~x5 & ~n267 ;
  assign n269 = ~n265 & n268 ;
  assign n270 = ~n236 & n269 ;
  assign n271 = ~n233 & ~n270 ;
  assign n273 = ~x2 & ~x15 ;
  assign n274 = n24 & n273 ;
  assign n275 = ~n45 & ~n274 ;
  assign n272 = ~x8 & n24 ;
  assign n276 = n275 ^ n272 ;
  assign n277 = n276 ^ x4 ;
  assign n286 = n277 ^ n276 ;
  assign n278 = n26 & n134 ;
  assign n279 = n48 & n278 ;
  assign n280 = n279 ^ n277 ;
  assign n281 = n280 ^ n276 ;
  assign n282 = n279 ^ n272 ;
  assign n283 = n282 ^ n279 ;
  assign n284 = n283 ^ n281 ;
  assign n285 = ~n281 & ~n284 ;
  assign n287 = n286 ^ n285 ;
  assign n288 = n287 ^ n281 ;
  assign n289 = n25 & n168 ;
  assign n290 = n289 ^ n276 ;
  assign n291 = n285 ^ n281 ;
  assign n292 = n290 & ~n291 ;
  assign n293 = n292 ^ n276 ;
  assign n294 = ~n288 & ~n293 ;
  assign n295 = n294 ^ n276 ;
  assign n296 = n295 ^ n272 ;
  assign n297 = n296 ^ n276 ;
  assign n298 = ~n271 & ~n297 ;
  assign n299 = ~n51 & n298 ;
  assign n301 = n300 ^ n299 ;
  assign n302 = n301 ^ n299 ;
  assign n303 = n299 ^ x18 ;
  assign n304 = ~n302 & n303 ;
  assign n305 = n304 ^ n299 ;
  assign n306 = ~n41 & n305 ;
  assign n307 = x14 & ~n306 ;
  assign y0 = n307 ;
endmodule
