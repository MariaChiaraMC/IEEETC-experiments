module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 ;
  assign n9 = x0 & ~x3 ;
  assign n14 = x6 & x7 ;
  assign n15 = ~x5 & ~n14 ;
  assign n10 = ~x2 & x5 ;
  assign n11 = ~x6 & ~x7 ;
  assign n12 = x1 & ~n11 ;
  assign n13 = n10 & n12 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = ~x1 & x2 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = n19 ^ n13 ;
  assign n21 = ~n17 & n20 ;
  assign n22 = n21 ^ n13 ;
  assign n23 = x4 & n22 ;
  assign n24 = n23 ^ n13 ;
  assign n25 = n9 & n24 ;
  assign y0 = n25 ;
endmodule
