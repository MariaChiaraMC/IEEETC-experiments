module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 ;
  assign n16 = x4 & x6 ;
  assign n17 = x2 & ~x8 ;
  assign n18 = ~x1 & x5 ;
  assign n19 = n17 & n18 ;
  assign n20 = ~x0 & n19 ;
  assign n21 = ~n16 & ~n20 ;
  assign n22 = ~x12 & x13 ;
  assign n23 = n22 ^ x11 ;
  assign n24 = x14 ^ x4 ;
  assign n25 = n24 ^ x14 ;
  assign n26 = ~x9 & ~x10 ;
  assign n27 = ~x14 & n26 ;
  assign n28 = n27 ^ x14 ;
  assign n29 = ~n25 & n28 ;
  assign n30 = n29 ^ x14 ;
  assign n31 = n30 ^ n22 ;
  assign n32 = ~n23 & n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ x14 ;
  assign n35 = n34 ^ x11 ;
  assign n36 = n22 & ~n35 ;
  assign n37 = n36 ^ n22 ;
  assign n38 = ~n21 & n37 ;
  assign n39 = x9 & x10 ;
  assign n40 = ~x3 & n39 ;
  assign n41 = n40 ^ x6 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = x1 & ~x2 ;
  assign n44 = x0 & n43 ;
  assign n45 = ~x5 & n44 ;
  assign n46 = x4 & ~n45 ;
  assign n47 = x3 & x7 ;
  assign n48 = ~n46 & n47 ;
  assign n49 = n48 ^ n40 ;
  assign n50 = n42 & n49 ;
  assign n51 = n50 ^ n40 ;
  assign n52 = n38 & n51 ;
  assign y0 = n52 ;
endmodule
