module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 ;
  assign n85 = x3 & ~x5 ;
  assign n61 = ~x4 & x6 ;
  assign n86 = x1 & x7 ;
  assign n87 = n61 & ~n86 ;
  assign n88 = ~x2 & n87 ;
  assign n89 = x2 & x4 ;
  assign n90 = ~x1 & n89 ;
  assign n91 = ~x6 & n90 ;
  assign n92 = ~n88 & ~n91 ;
  assign n93 = n85 & ~n92 ;
  assign n9 = x4 & ~x7 ;
  assign n15 = ~x3 & ~x6 ;
  assign n73 = x2 & n15 ;
  assign n94 = n9 & n73 ;
  assign n95 = x3 & ~x4 ;
  assign n96 = ~n89 & ~n95 ;
  assign n97 = n96 ^ x6 ;
  assign n98 = n97 ^ n96 ;
  assign n99 = x7 ^ x4 ;
  assign n100 = n99 ^ x4 ;
  assign n101 = n100 ^ n96 ;
  assign n102 = n101 ^ n96 ;
  assign n103 = n102 ^ n98 ;
  assign n30 = x2 & x3 ;
  assign n104 = n99 ^ n30 ;
  assign n105 = n104 ^ n98 ;
  assign n106 = ~n99 & ~n105 ;
  assign n107 = n106 ^ n96 ;
  assign n108 = ~n103 & n107 ;
  assign n109 = n108 ^ n106 ;
  assign n110 = n109 ^ n96 ;
  assign n111 = n110 ^ n99 ;
  assign n112 = n98 & ~n111 ;
  assign n113 = n112 ^ n106 ;
  assign n114 = n113 ^ n99 ;
  assign n115 = ~x1 & ~n114 ;
  assign n116 = ~n94 & ~n115 ;
  assign n117 = x5 & ~n116 ;
  assign n118 = ~x5 & ~x6 ;
  assign n119 = n89 & n118 ;
  assign n120 = ~x7 & ~n119 ;
  assign n16 = n15 ^ x2 ;
  assign n121 = n15 ^ x4 ;
  assign n122 = n121 ^ x4 ;
  assign n123 = n122 ^ n16 ;
  assign n124 = n61 ^ x3 ;
  assign n125 = n61 & n124 ;
  assign n126 = n125 ^ x4 ;
  assign n127 = n126 ^ n61 ;
  assign n128 = ~n123 & n127 ;
  assign n129 = n128 ^ n125 ;
  assign n130 = n129 ^ n61 ;
  assign n131 = n16 & n130 ;
  assign n132 = n131 ^ n15 ;
  assign n133 = x5 & n132 ;
  assign n134 = n95 & n118 ;
  assign n135 = x2 & n134 ;
  assign n136 = x7 & ~n135 ;
  assign n137 = ~n133 & n136 ;
  assign n138 = x3 ^ x2 ;
  assign n139 = n138 ^ x5 ;
  assign n140 = n139 ^ x4 ;
  assign n141 = x6 ^ x2 ;
  assign n142 = n141 ^ x2 ;
  assign n143 = x5 ^ x2 ;
  assign n144 = n143 ^ x2 ;
  assign n145 = n142 & ~n144 ;
  assign n146 = n145 ^ x2 ;
  assign n147 = n146 ^ n139 ;
  assign n148 = ~n140 & n147 ;
  assign n149 = n148 ^ n145 ;
  assign n150 = n149 ^ x2 ;
  assign n151 = n150 ^ x4 ;
  assign n152 = ~n139 & ~n151 ;
  assign n153 = n152 ^ n139 ;
  assign n154 = n137 & n153 ;
  assign n155 = x1 & ~n154 ;
  assign n156 = ~n120 & n155 ;
  assign n157 = ~n117 & ~n156 ;
  assign n158 = ~n93 & n157 ;
  assign n58 = ~x1 & ~x2 ;
  assign n59 = x3 & x7 ;
  assign n60 = ~x6 & n59 ;
  assign n62 = ~n60 & ~n61 ;
  assign n63 = n58 & ~n62 ;
  assign n64 = x4 & n60 ;
  assign n26 = ~x3 & x7 ;
  assign n27 = x6 & n26 ;
  assign n65 = n27 ^ x4 ;
  assign n66 = n65 ^ n27 ;
  assign n67 = n27 ^ n15 ;
  assign n68 = ~n66 & n67 ;
  assign n69 = n68 ^ n27 ;
  assign n70 = x2 & n69 ;
  assign n71 = ~n64 & ~n70 ;
  assign n72 = x1 & ~n71 ;
  assign n74 = ~x4 & x7 ;
  assign n75 = n73 & n74 ;
  assign n28 = x1 & ~x2 ;
  assign n76 = n9 & n28 ;
  assign n77 = x6 ^ x3 ;
  assign n78 = n76 & ~n77 ;
  assign n79 = ~n75 & ~n78 ;
  assign n80 = ~n72 & n79 ;
  assign n81 = ~n63 & n80 ;
  assign n10 = x2 & x6 ;
  assign n11 = n10 ^ x1 ;
  assign n12 = n10 ^ x3 ;
  assign n13 = n12 ^ x3 ;
  assign n14 = n13 ^ n11 ;
  assign n17 = n15 & ~n16 ;
  assign n18 = n17 ^ x3 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n14 & n19 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n21 ^ n15 ;
  assign n23 = ~n11 & n22 ;
  assign n24 = n23 ^ n10 ;
  assign n25 = n9 & n24 ;
  assign n29 = n27 & n28 ;
  assign n31 = x7 ^ x1 ;
  assign n32 = n30 & n31 ;
  assign n33 = x6 & ~n32 ;
  assign n34 = ~x4 & ~n33 ;
  assign n35 = x3 ^ x1 ;
  assign n43 = n35 ^ x3 ;
  assign n44 = n43 ^ x3 ;
  assign n45 = ~n43 & ~n44 ;
  assign n36 = n35 ^ x7 ;
  assign n37 = n36 ^ x2 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = n36 ^ n35 ;
  assign n40 = n39 ^ x3 ;
  assign n41 = ~n38 & ~n40 ;
  assign n48 = n45 ^ n41 ;
  assign n42 = n41 ^ x6 ;
  assign n46 = n45 ^ n43 ;
  assign n47 = n42 & ~n46 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = x6 & n49 ;
  assign n51 = n50 ^ n41 ;
  assign n52 = n51 ^ n45 ;
  assign n53 = n52 ^ n47 ;
  assign n54 = n53 ^ x6 ;
  assign n55 = n34 & n54 ;
  assign n56 = ~n29 & ~n55 ;
  assign n57 = ~n25 & n56 ;
  assign n82 = n81 ^ n57 ;
  assign n83 = ~x5 & n82 ;
  assign n84 = n83 ^ n81 ;
  assign n159 = n158 ^ n84 ;
  assign n160 = n159 ^ n158 ;
  assign n161 = n58 & n64 ;
  assign n162 = n161 ^ n158 ;
  assign n163 = n162 ^ n158 ;
  assign n164 = n160 & ~n163 ;
  assign n165 = n164 ^ n158 ;
  assign n166 = ~x0 & n165 ;
  assign n167 = n166 ^ n158 ;
  assign y0 = ~n167 ;
endmodule
