module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 ;
  assign n13 = x9 & ~x11 ;
  assign n14 = x2 & n13 ;
  assign n15 = x7 & x8 ;
  assign n16 = x4 & ~x10 ;
  assign n17 = n15 & n16 ;
  assign n18 = ~x5 & x6 ;
  assign n19 = ~x3 & n18 ;
  assign n20 = n17 & n19 ;
  assign n21 = n14 & n20 ;
  assign n22 = x5 & ~x6 ;
  assign n23 = ~x8 & ~x11 ;
  assign n24 = x4 & n23 ;
  assign n25 = x7 & n24 ;
  assign n26 = x3 & n25 ;
  assign n27 = n26 ^ x9 ;
  assign n28 = n27 ^ x2 ;
  assign n65 = n28 ^ n27 ;
  assign n35 = x8 ^ x7 ;
  assign n29 = x4 ^ x2 ;
  assign n30 = x8 ^ x4 ;
  assign n31 = n30 ^ x3 ;
  assign n32 = n31 ^ x4 ;
  assign n33 = n29 & ~n32 ;
  assign n34 = n33 ^ n31 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = x10 ^ x4 ;
  assign n38 = x3 ^ x2 ;
  assign n39 = n38 ^ x4 ;
  assign n40 = n39 ^ n31 ;
  assign n41 = ~n37 & ~n40 ;
  assign n42 = n41 ^ x10 ;
  assign n43 = n42 ^ x4 ;
  assign n44 = n43 ^ n39 ;
  assign n45 = n44 ^ n31 ;
  assign n46 = n45 ^ n29 ;
  assign n47 = n40 ^ n35 ;
  assign n48 = n39 ^ n29 ;
  assign n49 = n48 ^ n35 ;
  assign n50 = n47 & n49 ;
  assign n51 = n50 ^ n39 ;
  assign n52 = n51 ^ n31 ;
  assign n53 = n46 & ~n52 ;
  assign n54 = n53 ^ n35 ;
  assign n55 = ~n36 & ~n54 ;
  assign n56 = n55 ^ n53 ;
  assign n57 = n56 ^ n35 ;
  assign n58 = ~x11 & ~n57 ;
  assign n59 = n58 ^ n28 ;
  assign n60 = n59 ^ n27 ;
  assign n61 = n28 ^ n26 ;
  assign n62 = n61 ^ n58 ;
  assign n63 = n62 ^ n60 ;
  assign n64 = ~n60 & ~n63 ;
  assign n66 = n65 ^ n64 ;
  assign n67 = n66 ^ n60 ;
  assign n68 = ~x7 & n23 ;
  assign n69 = ~n17 & ~n68 ;
  assign n70 = n69 ^ n27 ;
  assign n71 = n64 ^ n60 ;
  assign n72 = n70 & ~n71 ;
  assign n73 = n72 ^ n27 ;
  assign n74 = ~n67 & n73 ;
  assign n75 = n74 ^ n27 ;
  assign n76 = n75 ^ x9 ;
  assign n77 = n76 ^ n27 ;
  assign n78 = n22 & n77 ;
  assign n79 = ~n21 & ~n78 ;
  assign n80 = x0 & x1 ;
  assign n81 = ~n79 & n80 ;
  assign y0 = n81 ;
endmodule
