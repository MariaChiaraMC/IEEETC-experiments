module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 ;
  output y0 ;
  wire n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 ;
  assign n21 = ~x13 & ~x18 ;
  assign n22 = x2 & n21 ;
  assign n23 = x9 & x13 ;
  assign n24 = x1 & n23 ;
  assign n25 = ~n22 & ~n24 ;
  assign n27 = ~x10 & ~x12 ;
  assign n28 = ~x11 & n27 ;
  assign n26 = ~x2 & x13 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = ~x6 & ~x7 ;
  assign n32 = ~x5 & n31 ;
  assign n33 = ~x4 & n32 ;
  assign n34 = n21 & ~n33 ;
  assign n35 = n34 ^ n26 ;
  assign n36 = n30 & n35 ;
  assign n37 = n36 ^ n26 ;
  assign n38 = ~x9 & n37 ;
  assign n39 = n25 & ~n38 ;
  assign n40 = ~x0 & ~x19 ;
  assign n41 = ~n39 & n40 ;
  assign n42 = x15 & n41 ;
  assign n43 = x15 ^ x13 ;
  assign n44 = x0 & x3 ;
  assign n45 = n44 ^ n43 ;
  assign n46 = x18 ^ x15 ;
  assign n47 = n46 ^ x18 ;
  assign n48 = x18 ^ x8 ;
  assign n49 = ~n47 & ~n48 ;
  assign n50 = n49 ^ x18 ;
  assign n51 = n50 ^ n43 ;
  assign n52 = n45 & ~n51 ;
  assign n53 = n52 ^ n49 ;
  assign n54 = n53 ^ x18 ;
  assign n55 = n54 ^ n44 ;
  assign n56 = n43 & ~n55 ;
  assign n57 = n56 ^ n43 ;
  assign n58 = ~n42 & ~n57 ;
  assign n59 = ~x16 & ~x17 ;
  assign n60 = ~x14 & n59 ;
  assign n61 = ~n58 & n60 ;
  assign y0 = n61 ;
endmodule
