module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n9 = x2 ^ x1 ;
  assign n10 = n9 ^ x1 ;
  assign n11 = n10 ^ x0 ;
  assign n12 = ~x6 & ~x7 ;
  assign n13 = ~x1 & ~x3 ;
  assign n14 = ~x4 & ~x5 ;
  assign n15 = n13 & n14 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = n12 & n16 ;
  assign n18 = n17 ^ x1 ;
  assign n19 = n18 ^ n12 ;
  assign n20 = n11 & n19 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n21 ^ n12 ;
  assign n23 = ~x0 & n22 ;
  assign n24 = n23 ^ x0 ;
  assign y0 = ~n24 ;
endmodule
