module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 ;
  assign n22 = ~x0 & ~x1 ;
  assign n23 = n22 ^ x5 ;
  assign n24 = ~x1 & ~x3 ;
  assign n25 = n24 ^ x2 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = ~x1 & x3 ;
  assign n28 = x0 & ~n27 ;
  assign n29 = n28 ^ n24 ;
  assign n30 = ~n26 & ~n29 ;
  assign n31 = n30 ^ n24 ;
  assign n32 = n31 ^ n22 ;
  assign n33 = ~n23 & ~n32 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ n24 ;
  assign n36 = n35 ^ x5 ;
  assign n37 = ~n22 & n36 ;
  assign n38 = n37 ^ n22 ;
  assign n39 = ~x4 & ~n38 ;
  assign n162 = ~x19 & ~x20 ;
  assign n40 = ~x3 & n22 ;
  assign n41 = ~x10 & x11 ;
  assign n42 = x8 & n41 ;
  assign n43 = ~x6 & ~x7 ;
  assign n44 = x9 & n43 ;
  assign n45 = n42 & n44 ;
  assign n46 = ~x8 & ~x11 ;
  assign n47 = n44 & n46 ;
  assign n48 = ~n45 & ~n47 ;
  assign n49 = x3 & ~n48 ;
  assign n50 = ~x0 & n49 ;
  assign n51 = x8 & x10 ;
  assign n52 = x9 & n51 ;
  assign n53 = ~x11 & n52 ;
  assign n54 = n27 & n53 ;
  assign n55 = n43 & n46 ;
  assign n56 = x10 & n55 ;
  assign n57 = n22 & n56 ;
  assign n58 = ~n54 & ~n57 ;
  assign n59 = ~n50 & n58 ;
  assign n60 = ~x12 & ~x13 ;
  assign n61 = ~x5 & n60 ;
  assign n62 = ~n59 & n61 ;
  assign n63 = ~n40 & ~n62 ;
  assign n64 = ~x2 & ~n63 ;
  assign n65 = ~n47 & ~n53 ;
  assign n66 = ~n45 & n65 ;
  assign n67 = ~n56 & n66 ;
  assign n68 = n60 & ~n67 ;
  assign n69 = x2 & ~x3 ;
  assign n70 = x1 & n69 ;
  assign n71 = n68 & n70 ;
  assign n72 = n45 & n60 ;
  assign n73 = n27 & n72 ;
  assign n74 = n73 ^ x5 ;
  assign n75 = n74 ^ n73 ;
  assign n76 = ~x0 & x2 ;
  assign n77 = ~x9 & ~x10 ;
  assign n78 = ~x8 & x11 ;
  assign n79 = n77 & n78 ;
  assign n80 = x13 & n79 ;
  assign n81 = ~x8 & n43 ;
  assign n82 = n41 & n81 ;
  assign n83 = ~x12 & n82 ;
  assign n84 = ~x9 & n83 ;
  assign n85 = ~n80 & ~n84 ;
  assign n86 = ~n68 & n85 ;
  assign n87 = n76 & ~n86 ;
  assign n88 = ~n56 & ~n82 ;
  assign n89 = ~x9 & n88 ;
  assign n90 = n60 & ~n89 ;
  assign n91 = x3 & ~n80 ;
  assign n92 = ~n90 & n91 ;
  assign n93 = ~n27 & ~n92 ;
  assign n94 = ~n87 & ~n93 ;
  assign n95 = n94 ^ n73 ;
  assign n96 = n75 & ~n95 ;
  assign n97 = n96 ^ n73 ;
  assign n98 = ~n71 & ~n97 ;
  assign n99 = ~n64 & n98 ;
  assign n100 = ~x4 & ~n99 ;
  assign n101 = ~x1 & ~x8 ;
  assign n102 = ~x10 & ~n101 ;
  assign n103 = x11 & ~x12 ;
  assign n104 = ~n102 & n103 ;
  assign n105 = x9 & n104 ;
  assign n106 = x13 ^ x1 ;
  assign n107 = x13 ^ x0 ;
  assign n108 = n107 ^ x0 ;
  assign n109 = ~x2 & ~x12 ;
  assign n110 = x9 & n46 ;
  assign n111 = ~x10 & n110 ;
  assign n112 = ~n109 & ~n111 ;
  assign n113 = n112 ^ x0 ;
  assign n114 = n108 & ~n113 ;
  assign n115 = n114 ^ x0 ;
  assign n116 = n106 & n115 ;
  assign n117 = n116 ^ x1 ;
  assign n118 = ~n105 & ~n117 ;
  assign n119 = ~x3 & ~n118 ;
  assign n120 = n27 ^ x2 ;
  assign n121 = n27 ^ x4 ;
  assign n122 = n121 ^ x4 ;
  assign n123 = x16 & n43 ;
  assign n124 = x15 ^ x12 ;
  assign n125 = x13 & n124 ;
  assign n126 = n125 ^ x12 ;
  assign n127 = n123 & ~n126 ;
  assign n128 = ~x1 & n79 ;
  assign n129 = n127 & n128 ;
  assign n130 = ~x17 & n129 ;
  assign n131 = n130 ^ x4 ;
  assign n132 = ~n122 & ~n131 ;
  assign n133 = n132 ^ x4 ;
  assign n134 = n120 & n133 ;
  assign n135 = ~n119 & ~n134 ;
  assign n136 = x5 & ~n135 ;
  assign n137 = ~x1 & n72 ;
  assign n138 = ~n52 & ~n81 ;
  assign n139 = ~x4 & ~x11 ;
  assign n140 = ~n77 & n139 ;
  assign n141 = n60 & n140 ;
  assign n142 = ~n138 & n141 ;
  assign n143 = ~n128 & ~n142 ;
  assign n144 = ~n137 & n143 ;
  assign n145 = n69 & ~n144 ;
  assign n146 = x3 & ~x5 ;
  assign n147 = ~n24 & ~n146 ;
  assign n148 = x4 & ~n147 ;
  assign n149 = ~x2 & n27 ;
  assign n150 = n55 & n149 ;
  assign n151 = n60 & n150 ;
  assign n152 = x9 & n151 ;
  assign n153 = ~n148 & ~n152 ;
  assign n154 = ~n145 & n153 ;
  assign n155 = x0 & ~n154 ;
  assign n156 = ~n76 & ~n146 ;
  assign n157 = x4 & ~n156 ;
  assign n158 = x1 & n157 ;
  assign n159 = ~n155 & ~n158 ;
  assign n160 = ~n136 & n159 ;
  assign n161 = ~n100 & n160 ;
  assign n163 = n162 ^ n161 ;
  assign n164 = n163 ^ n161 ;
  assign n165 = n161 ^ x18 ;
  assign n166 = ~n164 & n165 ;
  assign n167 = n166 ^ n161 ;
  assign n168 = ~n39 & n167 ;
  assign n169 = x14 & ~n168 ;
  assign y0 = n169 ;
endmodule
