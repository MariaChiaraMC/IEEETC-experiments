module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 ;
  assign n12 = ~x1 & ~x6 ;
  assign n13 = ~x3 & ~x5 ;
  assign n14 = x2 & n13 ;
  assign n15 = n12 & n14 ;
  assign n10 = ~x3 & ~x4 ;
  assign n16 = x1 & x5 ;
  assign n17 = x6 & x7 ;
  assign n18 = ~x2 & n17 ;
  assign n19 = ~n16 & ~n18 ;
  assign n20 = n10 & ~n19 ;
  assign n21 = x4 ^ x2 ;
  assign n22 = n21 ^ x6 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n23 ^ x3 ;
  assign n25 = n21 ^ x4 ;
  assign n26 = n25 ^ x5 ;
  assign n27 = ~x5 & n26 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = n28 ^ x5 ;
  assign n30 = ~n24 & ~n29 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n31 ^ x5 ;
  assign n33 = ~x3 & ~n32 ;
  assign n34 = n33 ^ x2 ;
  assign n35 = x1 & n34 ;
  assign n36 = n35 ^ n20 ;
  assign n37 = ~x2 & x5 ;
  assign n38 = x3 & x7 ;
  assign n39 = ~n37 & ~n38 ;
  assign n40 = n12 & ~n39 ;
  assign n41 = ~x3 & ~x6 ;
  assign n42 = ~n13 & ~n41 ;
  assign n43 = ~x5 & ~x6 ;
  assign n44 = x2 & ~n43 ;
  assign n45 = n42 & n44 ;
  assign n46 = ~n40 & ~n45 ;
  assign n47 = n46 ^ x4 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = ~x7 & ~n42 ;
  assign n50 = n49 ^ x2 ;
  assign n51 = n49 ^ n13 ;
  assign n52 = n51 ^ n13 ;
  assign n53 = n52 ^ n50 ;
  assign n54 = x6 & ~x7 ;
  assign n55 = x6 ^ x5 ;
  assign n56 = x3 & ~n55 ;
  assign n57 = ~n54 & ~n56 ;
  assign n58 = n57 ^ x1 ;
  assign n59 = ~n57 & n58 ;
  assign n60 = n59 ^ n13 ;
  assign n61 = n60 ^ n57 ;
  assign n62 = n53 & n61 ;
  assign n63 = n62 ^ n59 ;
  assign n64 = n63 ^ n57 ;
  assign n65 = ~n50 & ~n64 ;
  assign n66 = n65 ^ n49 ;
  assign n67 = n66 ^ n46 ;
  assign n68 = n48 & ~n67 ;
  assign n69 = n68 ^ n46 ;
  assign n70 = n69 ^ n20 ;
  assign n71 = n36 & ~n70 ;
  assign n72 = n71 ^ n68 ;
  assign n73 = n72 ^ n46 ;
  assign n74 = n73 ^ n35 ;
  assign n75 = ~n20 & ~n74 ;
  assign n76 = n75 ^ n20 ;
  assign n77 = ~n15 & ~n76 ;
  assign n9 = ~x1 & ~x2 ;
  assign n11 = n9 & n10 ;
  assign n78 = n77 ^ n11 ;
  assign n79 = n78 ^ x0 ;
  assign n87 = n79 ^ n78 ;
  assign n80 = ~x6 & ~x7 ;
  assign n81 = n80 ^ n79 ;
  assign n82 = n81 ^ n78 ;
  assign n83 = n80 ^ n11 ;
  assign n84 = n83 ^ n80 ;
  assign n85 = n84 ^ n82 ;
  assign n86 = n82 & n85 ;
  assign n88 = n87 ^ n86 ;
  assign n89 = n88 ^ n82 ;
  assign n90 = n78 ^ x5 ;
  assign n91 = n86 ^ n82 ;
  assign n92 = ~n90 & n91 ;
  assign n93 = n92 ^ n78 ;
  assign n94 = ~n89 & ~n93 ;
  assign n95 = n94 ^ n78 ;
  assign n96 = n95 ^ n11 ;
  assign n97 = n96 ^ n78 ;
  assign y0 = n97 ;
endmodule
