module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 ;
  assign n20 = ~x6 & x16 ;
  assign n22 = x8 & ~x18 ;
  assign n21 = ~x7 & x17 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ n20 ;
  assign n26 = ~x8 & x18 ;
  assign n27 = x7 & ~x17 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = n26 & ~n28 ;
  assign n30 = n29 ^ n22 ;
  assign n31 = n30 ^ n26 ;
  assign n32 = n25 & n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ n26 ;
  assign n35 = ~n20 & n34 ;
  assign n36 = n35 ^ n20 ;
  assign n37 = x16 ^ x6 ;
  assign n38 = n37 ^ x6 ;
  assign n39 = ~x6 & ~n27 ;
  assign n40 = ~x6 & ~n22 ;
  assign n41 = ~n39 & ~n40 ;
  assign n42 = n41 ^ x6 ;
  assign n43 = n38 & ~n42 ;
  assign n44 = n43 ^ x6 ;
  assign n45 = ~x15 & ~n44 ;
  assign n46 = n36 & n45 ;
  assign n47 = x14 & ~n46 ;
  assign n48 = ~x0 & ~n47 ;
  assign n49 = ~x2 & x15 ;
  assign n50 = n41 & n49 ;
  assign n51 = ~n21 & ~n27 ;
  assign n52 = x9 ^ x8 ;
  assign n53 = x18 ^ x9 ;
  assign n54 = n52 & n53 ;
  assign n55 = n54 ^ x8 ;
  assign n56 = n51 & ~n55 ;
  assign n57 = x6 & ~n21 ;
  assign n58 = n22 & ~n57 ;
  assign n59 = ~n56 & ~n58 ;
  assign n60 = n50 & ~n59 ;
  assign n61 = ~x10 & n60 ;
  assign n62 = n61 ^ x16 ;
  assign n63 = n62 ^ n61 ;
  assign n64 = n63 ^ x14 ;
  assign n65 = x7 & ~x10 ;
  assign n66 = n55 & n65 ;
  assign n67 = ~x17 & ~x18 ;
  assign n68 = n67 ^ x15 ;
  assign n69 = x18 & ~n65 ;
  assign n70 = x17 & n69 ;
  assign n71 = n70 ^ n67 ;
  assign n72 = n71 ^ n70 ;
  assign n73 = n72 ^ n68 ;
  assign n74 = x12 & x13 ;
  assign n75 = x1 & ~x11 ;
  assign n76 = n75 ^ n74 ;
  assign n77 = ~n74 & ~n76 ;
  assign n78 = n77 ^ n70 ;
  assign n79 = n78 ^ n74 ;
  assign n80 = n73 & n79 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n81 ^ n74 ;
  assign n83 = n68 & ~n82 ;
  assign n84 = ~n66 & n83 ;
  assign n85 = x17 ^ x8 ;
  assign n86 = x17 ^ x7 ;
  assign n87 = n86 ^ x7 ;
  assign n88 = x9 ^ x7 ;
  assign n89 = ~n87 & ~n88 ;
  assign n90 = n89 ^ x7 ;
  assign n91 = n85 & ~n90 ;
  assign n92 = n49 & ~n91 ;
  assign n93 = n39 & n92 ;
  assign n94 = ~x10 & ~n93 ;
  assign n95 = n94 ^ n84 ;
  assign n96 = n84 & ~n95 ;
  assign n97 = n96 ^ n61 ;
  assign n98 = n97 ^ n84 ;
  assign n99 = n64 & n98 ;
  assign n100 = n99 ^ n96 ;
  assign n101 = n100 ^ n84 ;
  assign n102 = ~x14 & n101 ;
  assign n103 = n102 ^ x14 ;
  assign n104 = n48 & n103 ;
  assign y0 = n104 ;
endmodule
