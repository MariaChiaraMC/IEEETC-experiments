// Benchmark "./pla/lin.rom.pla_dbb_orig_35NonExact" written by ABC on Fri Nov 20 10:23:14 2020

module \./pla/lin.rom.pla_dbb_orig_35NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = 1'b1;
endmodule


