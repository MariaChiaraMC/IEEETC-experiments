module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 ;
  assign n11 = x2 & ~x3 ;
  assign n12 = x1 & n11 ;
  assign n13 = ~x2 & x3 ;
  assign n14 = ~x1 & n13 ;
  assign n15 = ~n12 & ~n14 ;
  assign n16 = ~x0 & x5 ;
  assign n17 = x7 ^ x6 ;
  assign n18 = n17 ^ x7 ;
  assign n19 = n14 ^ x7 ;
  assign n20 = ~n18 & n19 ;
  assign n21 = n20 ^ x7 ;
  assign n22 = n16 & n21 ;
  assign n23 = ~n15 & n22 ;
  assign n229 = ~x0 & ~n15 ;
  assign n230 = x7 & ~n229 ;
  assign n96 = ~x1 & ~x2 ;
  assign n231 = ~x0 & n96 ;
  assign n232 = n231 ^ x5 ;
  assign n233 = x6 ^ x3 ;
  assign n234 = n231 ^ x3 ;
  assign n235 = n234 ^ x3 ;
  assign n236 = n233 & ~n235 ;
  assign n237 = n236 ^ x3 ;
  assign n238 = n232 & ~n237 ;
  assign n239 = n238 ^ x5 ;
  assign n240 = ~n230 & n239 ;
  assign n24 = x0 & ~x5 ;
  assign n25 = n12 & n24 ;
  assign n31 = ~x2 & x9 ;
  assign n32 = ~x0 & n31 ;
  assign n26 = ~x1 & x2 ;
  assign n27 = x0 & x5 ;
  assign n28 = n26 & n27 ;
  assign n33 = n32 ^ n28 ;
  assign n34 = n33 ^ n28 ;
  assign n29 = n28 ^ x5 ;
  assign n30 = n29 ^ n28 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n28 ^ x1 ;
  assign n37 = n36 ^ n28 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = n34 & n38 ;
  assign n40 = n39 ^ n34 ;
  assign n41 = ~n35 & n40 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = n42 ^ n28 ;
  assign n44 = n43 ^ n34 ;
  assign n45 = ~x3 & n44 ;
  assign n46 = n45 ^ n28 ;
  assign n47 = ~n25 & ~n46 ;
  assign n48 = ~x6 & ~n47 ;
  assign n49 = x0 & ~x1 ;
  assign n50 = n11 & n49 ;
  assign n51 = ~n26 & n27 ;
  assign n52 = ~x0 & x2 ;
  assign n53 = x8 & x9 ;
  assign n54 = ~x5 & n53 ;
  assign n55 = ~x1 & ~n54 ;
  assign n56 = n52 & ~n55 ;
  assign n57 = ~x3 & n56 ;
  assign n58 = ~n51 & ~n57 ;
  assign n59 = ~x6 & ~n58 ;
  assign n60 = ~x2 & ~x5 ;
  assign n61 = x9 ^ x8 ;
  assign n62 = n61 ^ x1 ;
  assign n63 = n62 ^ n60 ;
  assign n64 = x9 ^ x0 ;
  assign n65 = ~x1 & ~n64 ;
  assign n66 = n65 ^ x0 ;
  assign n67 = ~n63 & n66 ;
  assign n68 = n67 ^ n65 ;
  assign n69 = n68 ^ x0 ;
  assign n70 = n69 ^ x1 ;
  assign n71 = n60 & ~n70 ;
  assign n72 = x3 & ~x5 ;
  assign n73 = n16 ^ x6 ;
  assign n74 = n73 ^ x6 ;
  assign n75 = n74 ^ n72 ;
  assign n76 = n14 ^ n12 ;
  assign n77 = ~n14 & n76 ;
  assign n78 = n77 ^ x6 ;
  assign n79 = n78 ^ n14 ;
  assign n80 = ~n75 & ~n79 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n81 ^ n14 ;
  assign n83 = ~n72 & ~n82 ;
  assign n84 = n83 ^ n72 ;
  assign n85 = ~n71 & ~n84 ;
  assign n86 = ~n59 & n85 ;
  assign n87 = ~n50 & n86 ;
  assign n88 = n87 ^ x7 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = ~x3 & ~x5 ;
  assign n91 = x6 & ~x9 ;
  assign n92 = x0 & x1 ;
  assign n93 = ~x2 & ~x8 ;
  assign n94 = n92 & n93 ;
  assign n95 = ~n91 & n94 ;
  assign n97 = ~x0 & ~x6 ;
  assign n98 = x0 & x9 ;
  assign n99 = ~n97 & ~n98 ;
  assign n100 = n96 & ~n99 ;
  assign n101 = x1 & ~x9 ;
  assign n102 = n101 ^ n97 ;
  assign n103 = n102 ^ n101 ;
  assign n104 = x1 & ~n91 ;
  assign n105 = ~x8 & ~n104 ;
  assign n106 = n105 ^ n101 ;
  assign n107 = ~n103 & n106 ;
  assign n108 = n107 ^ n101 ;
  assign n109 = x2 & n108 ;
  assign n110 = ~n100 & ~n109 ;
  assign n111 = ~n95 & n110 ;
  assign n112 = n90 & ~n111 ;
  assign n113 = ~x6 & x9 ;
  assign n114 = ~x1 & n113 ;
  assign n115 = ~n101 & ~n114 ;
  assign n116 = n13 & n24 ;
  assign n117 = ~n115 & n116 ;
  assign n118 = ~x2 & ~x3 ;
  assign n119 = n27 & n114 ;
  assign n120 = n118 & n119 ;
  assign n121 = n120 ^ n117 ;
  assign n147 = ~x1 & ~x9 ;
  assign n128 = x1 & x3 ;
  assign n148 = n113 & n128 ;
  assign n149 = ~n147 & ~n148 ;
  assign n122 = x1 & ~n118 ;
  assign n123 = ~x0 & x9 ;
  assign n124 = n122 & ~n123 ;
  assign n125 = x9 ^ x6 ;
  assign n126 = ~x3 & ~n125 ;
  assign n127 = ~n96 & ~n126 ;
  assign n131 = n127 ^ x6 ;
  assign n132 = n131 ^ n127 ;
  assign n129 = n128 ^ n127 ;
  assign n130 = n129 ^ n127 ;
  assign n133 = n132 ^ n130 ;
  assign n134 = x3 & ~x9 ;
  assign n135 = n134 ^ n127 ;
  assign n136 = n135 ^ n127 ;
  assign n137 = n136 ^ n132 ;
  assign n138 = ~n132 & n137 ;
  assign n139 = n138 ^ n132 ;
  assign n140 = n133 & ~n139 ;
  assign n141 = n140 ^ n138 ;
  assign n142 = n141 ^ n127 ;
  assign n143 = n142 ^ n132 ;
  assign n144 = ~x0 & n143 ;
  assign n145 = n144 ^ n127 ;
  assign n146 = ~n124 & n145 ;
  assign n150 = n149 ^ n146 ;
  assign n151 = ~n52 & ~n150 ;
  assign n152 = n151 ^ n149 ;
  assign n153 = ~x5 & ~n152 ;
  assign n154 = x5 & ~x6 ;
  assign n155 = x2 ^ x0 ;
  assign n156 = n155 ^ x3 ;
  assign n157 = n156 ^ x1 ;
  assign n158 = n157 ^ x3 ;
  assign n159 = n158 ^ x9 ;
  assign n160 = x3 ^ x1 ;
  assign n161 = n160 ^ n159 ;
  assign n162 = x9 ^ x2 ;
  assign n163 = x2 & n162 ;
  assign n164 = n163 ^ x1 ;
  assign n165 = n164 ^ x2 ;
  assign n166 = ~n161 & n165 ;
  assign n167 = n166 ^ n163 ;
  assign n168 = n167 ^ x2 ;
  assign n169 = ~n159 & n168 ;
  assign n170 = n169 ^ n156 ;
  assign n171 = n154 & ~n170 ;
  assign n172 = ~n153 & ~n171 ;
  assign n173 = n172 ^ x8 ;
  assign n174 = n173 ^ n172 ;
  assign n175 = ~n52 & ~n97 ;
  assign n176 = n72 & ~n175 ;
  assign n177 = ~x5 & x6 ;
  assign n178 = n32 & n177 ;
  assign n179 = n154 ^ x5 ;
  assign n180 = x5 ^ x2 ;
  assign n181 = n180 ^ x5 ;
  assign n182 = ~n179 & ~n181 ;
  assign n183 = n182 ^ x5 ;
  assign n184 = n98 & ~n183 ;
  assign n185 = x3 & n184 ;
  assign n186 = ~n178 & ~n185 ;
  assign n187 = ~n176 & n186 ;
  assign n188 = ~x1 & ~n187 ;
  assign n189 = n52 ^ x3 ;
  assign n190 = n189 ^ n52 ;
  assign n191 = n190 ^ n154 ;
  assign n192 = ~n31 & n92 ;
  assign n193 = n192 ^ n32 ;
  assign n194 = ~n32 & n193 ;
  assign n195 = n194 ^ n52 ;
  assign n196 = n195 ^ n32 ;
  assign n197 = ~n191 & n196 ;
  assign n198 = n197 ^ n194 ;
  assign n199 = n198 ^ n32 ;
  assign n200 = n154 & ~n199 ;
  assign n201 = n200 ^ n154 ;
  assign n202 = x6 ^ x5 ;
  assign n203 = n13 ^ n11 ;
  assign n204 = n11 ^ x6 ;
  assign n205 = n204 ^ n11 ;
  assign n206 = n203 & n205 ;
  assign n207 = n206 ^ n11 ;
  assign n208 = n202 & n207 ;
  assign n209 = x9 ^ x1 ;
  assign n210 = ~n64 & n209 ;
  assign n211 = n208 & n210 ;
  assign n212 = ~n201 & ~n211 ;
  assign n213 = ~n188 & n212 ;
  assign n214 = n213 ^ n172 ;
  assign n215 = ~n174 & n214 ;
  assign n216 = n215 ^ n172 ;
  assign n217 = n216 ^ n117 ;
  assign n218 = n121 & ~n217 ;
  assign n219 = n218 ^ n215 ;
  assign n220 = n219 ^ n172 ;
  assign n221 = n220 ^ n120 ;
  assign n222 = ~n117 & ~n221 ;
  assign n223 = n222 ^ n117 ;
  assign n224 = ~n112 & ~n223 ;
  assign n225 = n224 ^ n87 ;
  assign n226 = ~n89 & n225 ;
  assign n227 = n226 ^ n87 ;
  assign n228 = ~n48 & n227 ;
  assign n241 = n240 ^ n228 ;
  assign n242 = x4 & n241 ;
  assign n243 = n242 ^ n228 ;
  assign n244 = ~n23 & n243 ;
  assign y0 = ~n244 ;
endmodule
