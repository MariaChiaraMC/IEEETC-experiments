module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ;
  assign n15 = x2 & x5 ;
  assign n16 = ~x6 & n15 ;
  assign n17 = ~x0 & x3 ;
  assign n18 = ~n16 & n17 ;
  assign n19 = ~x9 & ~x11 ;
  assign n20 = x1 & n19 ;
  assign n21 = ~x8 & ~x12 ;
  assign n22 = x7 & ~x13 ;
  assign n23 = n21 & n22 ;
  assign n24 = ~x10 & n15 ;
  assign n25 = n23 & n24 ;
  assign n26 = n20 & n25 ;
  assign n27 = n26 ^ x4 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = n28 ^ n18 ;
  assign n30 = ~x2 & ~x5 ;
  assign n31 = n30 ^ x1 ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = n32 ^ n26 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = ~n29 & n34 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = n18 & ~n37 ;
  assign n39 = n38 ^ n18 ;
  assign y0 = n39 ;
endmodule
