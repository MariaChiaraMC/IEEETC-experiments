module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n9 = x0 & x3 ;
  assign n10 = x6 & ~n9 ;
  assign n11 = ~x4 & n10 ;
  assign n12 = ~x2 & ~x3 ;
  assign n13 = ~x0 & n12 ;
  assign n14 = x5 & x7 ;
  assign n15 = ~n13 & n14 ;
  assign n16 = n11 & n15 ;
  assign n17 = n16 ^ x1 ;
  assign n18 = n16 ^ x0 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = x3 ^ x2 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = ~n19 & ~n21 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = ~x5 & ~x6 ;
  assign n25 = ~x4 & ~n24 ;
  assign n26 = ~n16 & n25 ;
  assign n27 = n26 ^ n17 ;
  assign n28 = ~n23 & n27 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = n17 & n29 ;
  assign n31 = n30 ^ n16 ;
  assign n32 = n31 ^ n17 ;
  assign y0 = ~n32 ;
endmodule
