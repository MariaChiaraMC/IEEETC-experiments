module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 ;
  assign n15 = x2 & x6 ;
  assign n16 = ~x1 & x5 ;
  assign n17 = ~x4 & ~n16 ;
  assign n18 = ~n15 & ~n17 ;
  assign n19 = ~x0 & ~n18 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = x5 & x7 ;
  assign n22 = ~x12 & n21 ;
  assign n23 = ~x8 & ~x10 ;
  assign n24 = ~x9 & ~x13 ;
  assign n25 = n23 & n24 ;
  assign n26 = x1 & ~x11 ;
  assign n27 = n25 & n26 ;
  assign n28 = n22 & n27 ;
  assign n29 = n28 ^ x4 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = x1 & x2 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = ~n30 & ~n32 ;
  assign n34 = n33 ^ n28 ;
  assign n35 = n34 ^ n19 ;
  assign n36 = n20 & n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ n28 ;
  assign n39 = n38 ^ x3 ;
  assign n40 = n19 & n39 ;
  assign n41 = n40 ^ n19 ;
  assign y0 = n41 ;
endmodule
