// Benchmark "./pla/sqr6.pla_11" written by ABC on Mon Apr 20 15:44:26 2020

module \./pla/sqr6.pla_11  ( 
    x0, x1, x2, x3, x4, x5,
    z0  );
  input  x0, x1, x2, x3, x4, x5;
  output z0;
  assign z0 = x5;
endmodule


