module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 ;
  output y0 ;
  wire n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 ;
  assign n23 = ~x0 & ~x1 ;
  assign n24 = ~x6 & ~x7 ;
  assign n25 = x11 & n24 ;
  assign n26 = ~x10 & n25 ;
  assign n27 = x8 & n26 ;
  assign n28 = x10 & ~x11 ;
  assign n29 = x8 & n28 ;
  assign n30 = ~n27 & ~n29 ;
  assign n31 = ~n23 & ~n30 ;
  assign n32 = ~x8 & ~x10 ;
  assign n33 = x0 & n32 ;
  assign n34 = x15 & x17 ;
  assign n35 = x10 & n34 ;
  assign n36 = x1 & n35 ;
  assign n37 = ~n33 & ~n36 ;
  assign n38 = ~x11 & n24 ;
  assign n39 = ~n37 & n38 ;
  assign n40 = ~n31 & ~n39 ;
  assign n41 = x9 & ~n40 ;
  assign n42 = ~x8 & n24 ;
  assign n43 = ~x1 & x9 ;
  assign n44 = x0 & ~n43 ;
  assign n45 = n28 & n44 ;
  assign n46 = n42 & n45 ;
  assign n47 = ~n41 & ~n46 ;
  assign n48 = ~x12 & ~x13 ;
  assign n49 = ~x4 & ~x5 ;
  assign n50 = n48 & n49 ;
  assign n51 = ~n47 & n50 ;
  assign n52 = x0 & x1 ;
  assign n53 = x5 & n52 ;
  assign n54 = ~x20 & n53 ;
  assign n55 = x1 ^ x0 ;
  assign n56 = x5 ^ x1 ;
  assign n57 = ~n55 & n56 ;
  assign n58 = n57 ^ x1 ;
  assign n59 = x12 & ~x13 ;
  assign n60 = ~x8 & ~x15 ;
  assign n61 = ~n59 & ~n60 ;
  assign n62 = n61 ^ x13 ;
  assign n63 = x9 & x10 ;
  assign n64 = n63 ^ n61 ;
  assign n65 = n64 ^ n63 ;
  assign n66 = n65 ^ n62 ;
  assign n67 = x11 & x16 ;
  assign n68 = n67 ^ n28 ;
  assign n69 = ~n28 & n68 ;
  assign n70 = n69 ^ n63 ;
  assign n71 = n70 ^ n28 ;
  assign n72 = ~n66 & n71 ;
  assign n73 = n72 ^ n69 ;
  assign n74 = n73 ^ n28 ;
  assign n75 = n62 & ~n74 ;
  assign n76 = n75 ^ n61 ;
  assign n77 = ~x17 & ~n76 ;
  assign n78 = x11 & ~x12 ;
  assign n79 = x7 & x8 ;
  assign n80 = n78 & n79 ;
  assign n81 = ~x9 & x13 ;
  assign n82 = ~x11 & ~x15 ;
  assign n83 = n42 & ~n82 ;
  assign n84 = ~n81 & ~n83 ;
  assign n85 = ~n80 & n84 ;
  assign n86 = x10 & ~n85 ;
  assign n88 = x16 ^ x13 ;
  assign n87 = x16 ^ x6 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = n89 ^ x7 ;
  assign n91 = n90 ^ n89 ;
  assign n92 = n91 ^ x6 ;
  assign n93 = x12 ^ x6 ;
  assign n94 = n93 ^ n89 ;
  assign n95 = n94 ^ n89 ;
  assign n96 = ~n92 & ~n95 ;
  assign n97 = n96 ^ x6 ;
  assign n98 = n89 ^ n88 ;
  assign n99 = n98 ^ x6 ;
  assign n100 = n99 ^ n92 ;
  assign n101 = n100 ^ n95 ;
  assign n103 = n88 ^ x11 ;
  assign n104 = n103 ^ n88 ;
  assign n105 = n101 & n104 ;
  assign n102 = ~n95 & n101 ;
  assign n106 = n105 ^ n102 ;
  assign n107 = n106 ^ n89 ;
  assign n108 = n107 ^ n104 ;
  assign n109 = n108 ^ n98 ;
  assign n110 = n109 ^ n92 ;
  assign n111 = x6 & n110 ;
  assign n112 = n111 ^ n105 ;
  assign n113 = n112 ^ n104 ;
  assign n114 = n113 ^ n92 ;
  assign n115 = n97 & ~n114 ;
  assign n116 = n115 ^ n102 ;
  assign n117 = n116 ^ n89 ;
  assign n118 = n117 ^ n98 ;
  assign n119 = n118 ^ x13 ;
  assign n120 = ~n86 & n119 ;
  assign n121 = n77 & n120 ;
  assign n122 = x10 ^ x8 ;
  assign n123 = x10 ^ x9 ;
  assign n124 = n123 ^ x9 ;
  assign n125 = ~x11 & x16 ;
  assign n126 = n125 ^ x9 ;
  assign n127 = n124 & ~n126 ;
  assign n128 = n127 ^ x9 ;
  assign n129 = ~n122 & n128 ;
  assign n130 = n129 ^ x8 ;
  assign n132 = n130 ^ n24 ;
  assign n142 = n132 ^ n130 ;
  assign n143 = n142 ^ n130 ;
  assign n144 = n142 & n143 ;
  assign n134 = ~x8 & n78 ;
  assign n135 = n134 ^ x12 ;
  assign n131 = n130 ^ x9 ;
  assign n133 = n132 ^ n131 ;
  assign n136 = n135 ^ n133 ;
  assign n137 = n136 ^ n133 ;
  assign n138 = n133 ^ n132 ;
  assign n139 = n138 ^ n130 ;
  assign n140 = n137 & n139 ;
  assign n147 = n144 ^ n140 ;
  assign n141 = n140 ^ n59 ;
  assign n145 = n144 ^ n142 ;
  assign n146 = n141 & n145 ;
  assign n148 = n147 ^ n146 ;
  assign n149 = n59 & n148 ;
  assign n150 = n149 ^ n140 ;
  assign n151 = n150 ^ n144 ;
  assign n152 = n151 ^ n146 ;
  assign n153 = n152 ^ n24 ;
  assign n154 = n121 & ~n153 ;
  assign n155 = ~x1 & n154 ;
  assign n156 = n155 ^ x4 ;
  assign n157 = ~n58 & n156 ;
  assign n158 = n157 ^ n155 ;
  assign n159 = x4 & n158 ;
  assign n160 = n159 ^ x4 ;
  assign n161 = ~n54 & ~n160 ;
  assign n162 = ~n51 & n161 ;
  assign n163 = x2 & ~n162 ;
  assign n168 = x4 & x5 ;
  assign n164 = ~x8 & ~x9 ;
  assign n165 = ~x10 & x11 ;
  assign n166 = n164 & n165 ;
  assign n167 = n49 & n166 ;
  assign n169 = n168 ^ n167 ;
  assign n170 = x2 & n169 ;
  assign n171 = n170 ^ n168 ;
  assign n172 = x0 & n171 ;
  assign n173 = ~x0 & ~x2 ;
  assign n174 = n49 & n173 ;
  assign n175 = x20 & x21 ;
  assign n176 = n174 & n175 ;
  assign n177 = x15 & n176 ;
  assign n178 = ~n172 & ~n177 ;
  assign n179 = n178 ^ x1 ;
  assign n180 = n179 ^ n178 ;
  assign n181 = n180 ^ x3 ;
  assign n182 = x0 & ~x13 ;
  assign n183 = n63 & n78 ;
  assign n184 = n182 & ~n183 ;
  assign n185 = n184 ^ n168 ;
  assign n186 = n168 & ~n185 ;
  assign n187 = n186 ^ n178 ;
  assign n188 = n187 ^ n168 ;
  assign n189 = ~n181 & ~n188 ;
  assign n190 = n189 ^ n186 ;
  assign n191 = n190 ^ n168 ;
  assign n192 = ~x3 & n191 ;
  assign n193 = n192 ^ x3 ;
  assign n194 = ~n163 & ~n193 ;
  assign n195 = ~x2 & n168 ;
  assign n196 = n23 & n195 ;
  assign n197 = ~x2 & n53 ;
  assign n198 = n24 & n32 ;
  assign n199 = x11 & n198 ;
  assign n200 = ~x9 & ~n199 ;
  assign n201 = n197 & ~n200 ;
  assign n209 = x8 & x10 ;
  assign n216 = ~n198 & ~n209 ;
  assign n217 = x5 & ~x11 ;
  assign n218 = ~n216 & n217 ;
  assign n219 = ~n27 & ~n218 ;
  assign n220 = n43 & ~n219 ;
  assign n202 = ~x5 & ~x11 ;
  assign n203 = ~x1 & x10 ;
  assign n204 = ~x9 & ~n203 ;
  assign n205 = n42 & ~n204 ;
  assign n206 = n205 ^ n43 ;
  assign n207 = n205 ^ x0 ;
  assign n208 = n207 ^ x0 ;
  assign n210 = n209 ^ x0 ;
  assign n211 = ~n208 & n210 ;
  assign n212 = n211 ^ x0 ;
  assign n213 = n206 & ~n212 ;
  assign n214 = n213 ^ n43 ;
  assign n215 = n202 & n214 ;
  assign n221 = n220 ^ n215 ;
  assign n222 = n221 ^ x2 ;
  assign n229 = n222 ^ n221 ;
  assign n223 = n222 ^ x5 ;
  assign n224 = n223 ^ n221 ;
  assign n225 = n222 ^ n215 ;
  assign n226 = n225 ^ x5 ;
  assign n227 = n226 ^ n224 ;
  assign n228 = ~n224 & ~n227 ;
  assign n230 = n229 ^ n228 ;
  assign n231 = n230 ^ n224 ;
  assign n232 = n221 ^ x0 ;
  assign n233 = n228 ^ n224 ;
  assign n234 = n232 & ~n233 ;
  assign n235 = n234 ^ n221 ;
  assign n236 = n231 & n235 ;
  assign n237 = n236 ^ n221 ;
  assign n238 = n237 ^ n220 ;
  assign n239 = n238 ^ n221 ;
  assign n240 = ~n201 & ~n239 ;
  assign n241 = n48 & ~n240 ;
  assign n242 = ~x8 & n165 ;
  assign n243 = n197 & n242 ;
  assign n244 = n81 & n243 ;
  assign n245 = ~n241 & ~n244 ;
  assign n246 = ~x4 & ~n245 ;
  assign n247 = x2 & x21 ;
  assign n248 = x4 & ~x5 ;
  assign n249 = n52 & n248 ;
  assign n250 = ~n247 & n249 ;
  assign n251 = x3 & ~n250 ;
  assign n252 = ~n246 & n251 ;
  assign n253 = ~n196 & n252 ;
  assign n254 = ~x18 & ~x19 ;
  assign n255 = x14 & n254 ;
  assign n256 = ~n253 & n255 ;
  assign n257 = ~n194 & n256 ;
  assign y0 = n257 ;
endmodule
