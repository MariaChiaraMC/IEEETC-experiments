module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 ;
  assign n8 = ~x3 & ~x4 ;
  assign n9 = x5 & x6 ;
  assign n10 = n8 & n9 ;
  assign n11 = x1 & n10 ;
  assign n12 = x0 & n11 ;
  assign n13 = x3 & x4 ;
  assign n14 = ~x5 & ~x6 ;
  assign n15 = n13 & ~n14 ;
  assign n16 = n15 ^ x0 ;
  assign n20 = n16 ^ n15 ;
  assign n17 = ~x3 & ~x5 ;
  assign n21 = n20 ^ n17 ;
  assign n18 = n17 ^ n16 ;
  assign n22 = n21 ^ n18 ;
  assign n19 = n18 ^ n16 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n23 ^ x2 ;
  assign n25 = n18 ^ x2 ;
  assign n26 = n24 & ~n25 ;
  assign n27 = n26 ^ n22 ;
  assign n28 = ~x3 & ~x6 ;
  assign n29 = x1 & ~n28 ;
  assign n30 = n29 ^ n16 ;
  assign n31 = n30 ^ n22 ;
  assign n32 = n31 ^ n23 ;
  assign n33 = n30 & n32 ;
  assign n34 = n30 ^ n18 ;
  assign n35 = n34 ^ n23 ;
  assign n36 = n35 ^ x2 ;
  assign n37 = n8 & ~n36 ;
  assign n38 = n37 ^ n8 ;
  assign n39 = n38 ^ n30 ;
  assign n40 = n39 ^ n23 ;
  assign n41 = n40 ^ x2 ;
  assign n42 = n33 & n41 ;
  assign n43 = n42 ^ x2 ;
  assign n44 = n27 & n43 ;
  assign n45 = n44 ^ n26 ;
  assign n46 = n45 ^ n42 ;
  assign n47 = n46 ^ n22 ;
  assign n48 = n47 ^ x2 ;
  assign n49 = n48 ^ x2 ;
  assign n50 = ~n12 & ~n49 ;
  assign n51 = x3 & x5 ;
  assign n52 = ~x1 & ~n51 ;
  assign n53 = ~n13 & n52 ;
  assign n54 = n53 ^ x0 ;
  assign n55 = n54 ^ n53 ;
  assign n56 = n55 ^ n54 ;
  assign n57 = n54 ^ n8 ;
  assign n58 = n57 ^ n54 ;
  assign n59 = ~n56 & n58 ;
  assign n60 = n59 ^ n54 ;
  assign n61 = n9 & ~n54 ;
  assign n62 = n61 ^ x2 ;
  assign n63 = ~n60 & n62 ;
  assign n64 = n63 ^ n61 ;
  assign n65 = x2 & n64 ;
  assign n66 = n65 ^ x2 ;
  assign n67 = n50 & ~n66 ;
  assign y0 = ~n67 ;
endmodule
