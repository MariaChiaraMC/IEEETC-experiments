module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n15 = ~x11 & ~x12 ;
  assign n16 = ~x13 & ~n15 ;
  assign n17 = x9 & ~n16 ;
  assign n18 = ~x9 & ~x13 ;
  assign n19 = ~x5 & ~x10 ;
  assign n20 = ~n18 & n19 ;
  assign n21 = x0 & x6 ;
  assign n22 = n21 ^ x11 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n21 ^ x12 ;
  assign n25 = n23 & ~n24 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = ~x9 & ~n21 ;
  assign n28 = n27 ^ n20 ;
  assign n29 = ~n26 & n28 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n20 & n30 ;
  assign n32 = n31 ^ n20 ;
  assign n33 = ~n17 & n32 ;
  assign y0 = n33 ;
endmodule
