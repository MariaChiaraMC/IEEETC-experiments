module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 ;
  assign n17 = ~x0 & ~x1 ;
  assign n18 = ~x6 & n17 ;
  assign n19 = ~x4 & ~x13 ;
  assign n20 = ~x8 & n19 ;
  assign n21 = n18 & n20 ;
  assign n22 = x14 ^ x2 ;
  assign n23 = x7 & x10 ;
  assign n24 = x3 & n23 ;
  assign n25 = n24 ^ x14 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n26 ^ n22 ;
  assign n28 = ~x3 & ~x7 ;
  assign n29 = ~x9 & ~x10 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = n28 & n30 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = n32 ^ n28 ;
  assign n34 = n27 & n33 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = n35 ^ n28 ;
  assign n37 = n22 & n36 ;
  assign n38 = n21 & n37 ;
  assign n39 = x2 & x13 ;
  assign n40 = ~x3 & n39 ;
  assign n41 = ~x1 & n40 ;
  assign n42 = x6 & ~n41 ;
  assign n71 = x3 & ~n39 ;
  assign n43 = x0 & x7 ;
  assign n44 = ~x13 & ~x14 ;
  assign n45 = n43 & n44 ;
  assign n46 = x1 & x4 ;
  assign n47 = ~x2 & x3 ;
  assign n48 = n46 & n47 ;
  assign n49 = n45 & n48 ;
  assign n72 = n71 ^ n49 ;
  assign n73 = n72 ^ n49 ;
  assign n50 = ~x7 & x8 ;
  assign n51 = x11 & n17 ;
  assign n52 = n50 & n51 ;
  assign n53 = ~x2 & x10 ;
  assign n54 = x9 & ~x13 ;
  assign n55 = n53 & n54 ;
  assign n56 = n52 & n55 ;
  assign n57 = x14 & n56 ;
  assign n58 = ~x8 & n29 ;
  assign n59 = ~x14 & n58 ;
  assign n60 = n43 ^ x13 ;
  assign n61 = n60 ^ n43 ;
  assign n62 = x2 & ~x7 ;
  assign n63 = n17 & n62 ;
  assign n64 = n63 ^ n43 ;
  assign n65 = ~n61 & n64 ;
  assign n66 = n65 ^ n43 ;
  assign n67 = n59 & n66 ;
  assign n68 = ~n57 & ~n67 ;
  assign n69 = n68 ^ n49 ;
  assign n70 = n69 ^ n49 ;
  assign n74 = n73 ^ n70 ;
  assign n75 = n49 ^ x4 ;
  assign n76 = n75 ^ n49 ;
  assign n77 = n76 ^ n73 ;
  assign n78 = ~n73 & n77 ;
  assign n79 = n78 ^ n73 ;
  assign n80 = n74 & ~n79 ;
  assign n81 = n80 ^ n78 ;
  assign n82 = n81 ^ n49 ;
  assign n83 = n82 ^ n73 ;
  assign n84 = ~x15 & ~n83 ;
  assign n85 = n84 ^ n49 ;
  assign n86 = n42 & n85 ;
  assign n87 = ~n38 & ~n86 ;
  assign n88 = ~x5 & ~n87 ;
  assign n89 = x5 & x10 ;
  assign n90 = x2 & x4 ;
  assign n91 = n18 & n90 ;
  assign n92 = n89 & n91 ;
  assign n93 = ~x9 & ~x15 ;
  assign n94 = n44 & n50 ;
  assign n95 = n93 & n94 ;
  assign n96 = n95 ^ x3 ;
  assign n97 = n96 ^ n95 ;
  assign n98 = x9 & x15 ;
  assign n99 = ~x8 & n98 ;
  assign n100 = x14 ^ x13 ;
  assign n101 = n99 & n100 ;
  assign n102 = n101 ^ n95 ;
  assign n103 = ~n97 & n102 ;
  assign n104 = n103 ^ n95 ;
  assign n105 = n92 & n104 ;
  assign n106 = ~n88 & ~n105 ;
  assign n107 = ~x12 & ~n106 ;
  assign y0 = n107 ;
endmodule
