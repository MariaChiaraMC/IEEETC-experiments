module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 ;
  output y0 ;
  wire n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 ;
  assign n19 = ~x16 & ~x17 ;
  assign n20 = ~x13 & n19 ;
  assign n21 = x10 & ~x14 ;
  assign n22 = n20 & n21 ;
  assign n23 = x12 ^ x11 ;
  assign n24 = n22 & n23 ;
  assign n25 = x1 & n24 ;
  assign n26 = ~x15 & ~n25 ;
  assign n27 = ~x0 & ~n26 ;
  assign n28 = ~x2 & ~x9 ;
  assign n29 = n28 ^ n19 ;
  assign n30 = x6 & x7 ;
  assign n31 = ~x5 & n30 ;
  assign n32 = x5 & ~x6 ;
  assign n33 = ~x7 & ~x8 ;
  assign n34 = n32 & n33 ;
  assign n35 = ~n31 & ~n34 ;
  assign n36 = n35 ^ n20 ;
  assign n37 = n29 & n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = n20 & n38 ;
  assign n40 = n39 ^ x13 ;
  assign n41 = n40 ^ x14 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = n42 ^ n27 ;
  assign n44 = x7 & x8 ;
  assign n45 = x17 & ~n44 ;
  assign n46 = x4 & n32 ;
  assign n47 = n45 & n46 ;
  assign n48 = x15 & ~n47 ;
  assign n49 = ~x16 & ~n48 ;
  assign n50 = n19 ^ x13 ;
  assign n51 = n19 ^ x3 ;
  assign n52 = n51 ^ x3 ;
  assign n53 = n31 ^ x3 ;
  assign n54 = n52 & ~n53 ;
  assign n55 = n54 ^ x3 ;
  assign n56 = ~n50 & n55 ;
  assign n57 = n56 ^ x13 ;
  assign n58 = ~n49 & ~n57 ;
  assign n59 = x7 ^ x6 ;
  assign n60 = n59 ^ x7 ;
  assign n61 = n60 ^ x17 ;
  assign n62 = n61 ^ n59 ;
  assign n63 = n62 ^ x5 ;
  assign n64 = n59 ^ x17 ;
  assign n65 = n64 ^ x8 ;
  assign n66 = ~x8 & ~n65 ;
  assign n67 = n66 ^ n59 ;
  assign n68 = n67 ^ x8 ;
  assign n69 = ~n63 & ~n68 ;
  assign n70 = n69 ^ n66 ;
  assign n71 = n70 ^ x8 ;
  assign n72 = x5 & ~n71 ;
  assign n73 = x4 & n72 ;
  assign n74 = x16 & n73 ;
  assign n75 = n74 ^ n58 ;
  assign n76 = n58 & ~n75 ;
  assign n77 = n76 ^ n40 ;
  assign n78 = n77 ^ n58 ;
  assign n79 = ~n43 & n78 ;
  assign n80 = n79 ^ n76 ;
  assign n81 = n80 ^ n58 ;
  assign n82 = n27 & n81 ;
  assign n83 = n82 ^ n27 ;
  assign y0 = n83 ;
endmodule
