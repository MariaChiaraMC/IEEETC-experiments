module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 ;
  output y0 ;
  wire n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 ;
  assign n24 = ~x0 & x1 ;
  assign n25 = ~x2 & n24 ;
  assign n26 = x0 & ~x1 ;
  assign n27 = x5 & n26 ;
  assign n28 = ~n25 & ~n27 ;
  assign n29 = x5 ^ x3 ;
  assign n30 = ~x4 & ~n29 ;
  assign n31 = ~n28 & n30 ;
  assign n249 = ~x19 & ~x20 ;
  assign n32 = ~x1 & x4 ;
  assign n33 = x8 & x10 ;
  assign n34 = x6 & x9 ;
  assign n35 = ~n33 & ~n34 ;
  assign n36 = x7 & ~n35 ;
  assign n37 = ~x6 & ~x7 ;
  assign n38 = ~x12 & n37 ;
  assign n39 = x15 & ~x16 ;
  assign n40 = ~x10 & ~n39 ;
  assign n41 = n38 & ~n40 ;
  assign n42 = ~n36 & ~n41 ;
  assign n43 = x11 & ~n42 ;
  assign n44 = x9 & x10 ;
  assign n45 = ~x12 & n44 ;
  assign n46 = ~n38 & ~n45 ;
  assign n47 = x10 & x15 ;
  assign n48 = ~x8 & ~n47 ;
  assign n49 = ~n46 & ~n48 ;
  assign n50 = ~x17 & ~n49 ;
  assign n63 = ~x10 & x11 ;
  assign n64 = x12 & ~n63 ;
  assign n65 = x11 & ~x16 ;
  assign n66 = x9 & ~x10 ;
  assign n67 = ~n65 & ~n66 ;
  assign n68 = ~x6 & ~x8 ;
  assign n69 = ~x15 & n68 ;
  assign n70 = n67 & n69 ;
  assign n71 = ~n64 & n70 ;
  assign n51 = x12 ^ x6 ;
  assign n52 = n51 ^ x12 ;
  assign n53 = n52 ^ x7 ;
  assign n54 = n44 ^ x16 ;
  assign n55 = x12 & n54 ;
  assign n56 = n55 ^ n44 ;
  assign n57 = n53 & n56 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = n58 ^ n44 ;
  assign n60 = n59 ^ x12 ;
  assign n61 = ~x7 & n60 ;
  assign n62 = n61 ^ x12 ;
  assign n72 = n71 ^ n62 ;
  assign n73 = ~x13 & ~n72 ;
  assign n74 = n73 ^ n71 ;
  assign n75 = n50 & n74 ;
  assign n76 = ~n43 & n75 ;
  assign n77 = x2 & ~n76 ;
  assign n78 = x11 & ~x12 ;
  assign n79 = ~x8 & n78 ;
  assign n80 = n79 ^ x13 ;
  assign n81 = n80 ^ x9 ;
  assign n88 = n81 ^ n80 ;
  assign n83 = x7 & n78 ;
  assign n82 = n81 ^ n79 ;
  assign n84 = n83 ^ n82 ;
  assign n85 = n83 ^ n81 ;
  assign n86 = n85 ^ n80 ;
  assign n87 = n84 & ~n86 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = x10 & ~x12 ;
  assign n91 = n90 ^ n81 ;
  assign n92 = n88 & n91 ;
  assign n93 = n92 ^ n90 ;
  assign n94 = n89 & n93 ;
  assign n95 = n94 ^ n87 ;
  assign n96 = n95 ^ n81 ;
  assign n97 = n96 ^ x13 ;
  assign n98 = n97 ^ n80 ;
  assign n99 = ~n77 & ~n98 ;
  assign n100 = n32 & ~n99 ;
  assign n101 = ~x11 & n66 ;
  assign n102 = ~x8 & n101 ;
  assign n103 = x12 & ~n102 ;
  assign n104 = ~x1 & ~x2 ;
  assign n105 = x13 & n104 ;
  assign n106 = ~n103 & n105 ;
  assign n110 = x2 & x4 ;
  assign n107 = ~x2 & ~x4 ;
  assign n108 = ~n32 & ~n107 ;
  assign n109 = n108 ^ x0 ;
  assign n111 = n110 ^ n109 ;
  assign n112 = n111 ^ n106 ;
  assign n113 = x1 & x13 ;
  assign n114 = n44 & n78 ;
  assign n115 = ~n113 & ~n114 ;
  assign n116 = x4 & ~n115 ;
  assign n117 = n116 ^ x0 ;
  assign n118 = n110 & ~n117 ;
  assign n119 = n118 ^ n116 ;
  assign n120 = n112 & ~n119 ;
  assign n121 = n120 ^ n118 ;
  assign n122 = n121 ^ n116 ;
  assign n123 = n122 ^ n110 ;
  assign n124 = ~n106 & ~n123 ;
  assign n125 = ~n100 & n124 ;
  assign n126 = ~x3 & ~n125 ;
  assign n127 = x1 & x2 ;
  assign n128 = n127 ^ x4 ;
  assign n129 = n128 ^ x4 ;
  assign n130 = x4 ^ x0 ;
  assign n131 = n130 ^ n128 ;
  assign n136 = n131 ^ n128 ;
  assign n137 = n136 ^ x4 ;
  assign n132 = n131 ^ x21 ;
  assign n133 = n132 ^ n131 ;
  assign n134 = n133 ^ x4 ;
  assign n135 = n134 ^ n129 ;
  assign n138 = n137 ^ n135 ;
  assign n139 = n129 & ~n138 ;
  assign n140 = n139 ^ n133 ;
  assign n141 = n140 ^ n137 ;
  assign n142 = n131 ^ n104 ;
  assign n143 = n142 ^ n131 ;
  assign n144 = n143 ^ n133 ;
  assign n145 = n144 ^ n129 ;
  assign n146 = n143 ^ x16 ;
  assign n147 = n146 ^ n133 ;
  assign n148 = n147 ^ x4 ;
  assign n149 = ~n145 & n148 ;
  assign n150 = n149 ^ x16 ;
  assign n151 = n150 ^ x4 ;
  assign n152 = n151 ^ n129 ;
  assign n153 = n152 ^ n137 ;
  assign n154 = n146 ^ x4 ;
  assign n155 = n154 ^ n129 ;
  assign n156 = n155 ^ n137 ;
  assign n157 = n148 ^ n129 ;
  assign n158 = n157 ^ n137 ;
  assign n159 = ~n156 & ~n158 ;
  assign n160 = n159 ^ x16 ;
  assign n161 = n160 ^ x4 ;
  assign n162 = n161 ^ n129 ;
  assign n163 = n153 & ~n162 ;
  assign n164 = n163 ^ n129 ;
  assign n165 = n164 ^ n137 ;
  assign n166 = ~n141 & ~n165 ;
  assign n167 = n166 ^ n139 ;
  assign n168 = n167 ^ n163 ;
  assign n169 = n168 ^ n133 ;
  assign n170 = n169 ^ n129 ;
  assign n171 = n170 ^ n127 ;
  assign n172 = ~n126 & n171 ;
  assign n173 = x5 & ~n172 ;
  assign n174 = x3 & x5 ;
  assign n175 = ~x0 & n104 ;
  assign n176 = ~x12 & ~x13 ;
  assign n177 = ~x7 & n68 ;
  assign n178 = n176 & n177 ;
  assign n179 = ~x9 & n107 ;
  assign n180 = x11 ^ x10 ;
  assign n181 = n179 & n180 ;
  assign n182 = n178 & n181 ;
  assign n183 = ~n175 & ~n182 ;
  assign n184 = ~n127 & n183 ;
  assign n185 = n174 & ~n184 ;
  assign n186 = ~x3 & n175 ;
  assign n187 = x10 & ~x11 ;
  assign n188 = n177 ^ n175 ;
  assign n189 = x8 & x9 ;
  assign n190 = n189 ^ n177 ;
  assign n191 = n190 ^ n189 ;
  assign n192 = ~x3 & ~x5 ;
  assign n193 = n24 & n192 ;
  assign n194 = n193 ^ n189 ;
  assign n195 = n191 & ~n194 ;
  assign n196 = n195 ^ n189 ;
  assign n197 = n188 & ~n196 ;
  assign n198 = n197 ^ n175 ;
  assign n199 = n187 & n198 ;
  assign n200 = ~x1 & n33 ;
  assign n201 = ~n177 & ~n200 ;
  assign n202 = x0 & ~x11 ;
  assign n203 = x9 & n202 ;
  assign n204 = x2 & n192 ;
  assign n205 = n203 & n204 ;
  assign n206 = ~n201 & n205 ;
  assign n207 = n37 & n189 ;
  assign n208 = n63 & n207 ;
  assign n209 = n193 & n208 ;
  assign n210 = ~n206 & ~n209 ;
  assign n211 = ~n199 & n210 ;
  assign n212 = n176 & ~n211 ;
  assign n213 = ~n186 & ~n212 ;
  assign n214 = n213 ^ x4 ;
  assign n215 = n214 ^ n213 ;
  assign n216 = x1 ^ x0 ;
  assign n217 = n216 ^ x3 ;
  assign n218 = x3 ^ x2 ;
  assign n219 = n218 ^ x3 ;
  assign n220 = n217 & n219 ;
  assign n221 = n220 ^ n216 ;
  assign n222 = n216 ^ x0 ;
  assign n223 = n222 ^ x3 ;
  assign n224 = n223 ^ n218 ;
  assign n225 = n216 ^ x22 ;
  assign n226 = n225 ^ x5 ;
  assign n227 = n224 & ~n226 ;
  assign n228 = n227 ^ x22 ;
  assign n229 = n228 ^ x5 ;
  assign n230 = n229 ^ x3 ;
  assign n231 = n216 ^ x5 ;
  assign n232 = n231 ^ n223 ;
  assign n233 = n223 ^ n217 ;
  assign n234 = n232 & ~n233 ;
  assign n235 = n234 ^ x3 ;
  assign n236 = n235 ^ n223 ;
  assign n237 = ~n230 & n236 ;
  assign n238 = n237 ^ x5 ;
  assign n239 = ~n221 & n238 ;
  assign n240 = n239 ^ n220 ;
  assign n241 = n240 ^ n237 ;
  assign n242 = n241 ^ n216 ;
  assign n243 = n242 ^ x5 ;
  assign n244 = n243 ^ n213 ;
  assign n245 = n215 & ~n244 ;
  assign n246 = n245 ^ n213 ;
  assign n247 = ~n185 & n246 ;
  assign n248 = ~n173 & n247 ;
  assign n250 = n249 ^ n248 ;
  assign n251 = n250 ^ n248 ;
  assign n252 = n248 ^ x18 ;
  assign n253 = ~n251 & n252 ;
  assign n254 = n253 ^ n248 ;
  assign n255 = ~n31 & n254 ;
  assign n256 = x14 & ~n255 ;
  assign y0 = n256 ;
endmodule
