module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 ;
  assign n11 = ~x6 & ~x7 ;
  assign n12 = x8 & ~x9 ;
  assign n13 = n11 & n12 ;
  assign n14 = ~x2 & ~x3 ;
  assign n15 = ~x4 & n14 ;
  assign n16 = ~x0 & x1 ;
  assign n17 = n15 & n16 ;
  assign n18 = n13 & n17 ;
  assign n19 = x6 & ~x9 ;
  assign n20 = ~x8 & n19 ;
  assign n21 = ~x2 & ~x7 ;
  assign n22 = x3 & n21 ;
  assign n23 = n20 & n22 ;
  assign n24 = ~x6 & x7 ;
  assign n25 = ~x8 & x9 ;
  assign n26 = n14 & ~n25 ;
  assign n27 = n24 & n26 ;
  assign n28 = ~n23 & ~n27 ;
  assign n29 = x4 & ~n28 ;
  assign n30 = x0 & x1 ;
  assign n31 = x8 & x9 ;
  assign n32 = n15 & n31 ;
  assign n33 = x7 ^ x6 ;
  assign n34 = n32 & ~n33 ;
  assign n35 = n30 & ~n34 ;
  assign n36 = ~n29 & n35 ;
  assign n37 = x3 & ~n31 ;
  assign n38 = x4 & ~n37 ;
  assign n39 = n11 & n38 ;
  assign n40 = x8 ^ x2 ;
  assign n41 = n40 ^ x9 ;
  assign n42 = x9 ^ x3 ;
  assign n43 = x8 ^ x3 ;
  assign n44 = ~n42 & n43 ;
  assign n45 = n44 ^ x3 ;
  assign n46 = n41 & ~n45 ;
  assign n47 = n46 ^ x2 ;
  assign n48 = n39 & n47 ;
  assign n49 = x3 & ~x4 ;
  assign n50 = n24 & n31 ;
  assign n51 = n50 ^ x7 ;
  assign n52 = n51 ^ n50 ;
  assign n53 = n50 ^ n19 ;
  assign n54 = n53 ^ n50 ;
  assign n55 = ~n52 & n54 ;
  assign n56 = n55 ^ n50 ;
  assign n57 = x2 & n56 ;
  assign n58 = n57 ^ n50 ;
  assign n59 = n49 & n58 ;
  assign n60 = ~n48 & ~n59 ;
  assign n61 = n36 & n60 ;
  assign n62 = x7 & ~x8 ;
  assign n63 = x9 ^ x6 ;
  assign n64 = x9 ^ x4 ;
  assign n65 = x4 ^ x3 ;
  assign n66 = n65 ^ x9 ;
  assign n67 = ~x9 & ~n66 ;
  assign n68 = n67 ^ x9 ;
  assign n69 = ~n64 & ~n68 ;
  assign n70 = n69 ^ n67 ;
  assign n71 = n70 ^ x9 ;
  assign n72 = n71 ^ n65 ;
  assign n73 = ~n63 & ~n72 ;
  assign n74 = n62 & n73 ;
  assign n75 = ~x4 & ~x6 ;
  assign n76 = n31 & n75 ;
  assign n77 = ~n20 & ~n76 ;
  assign n78 = ~x7 & ~n77 ;
  assign n79 = ~x3 & n78 ;
  assign n80 = ~n74 & ~n79 ;
  assign n81 = x2 & ~n80 ;
  assign n82 = x4 & ~x7 ;
  assign n83 = n12 & n82 ;
  assign n84 = n14 ^ x3 ;
  assign n85 = x6 & n84 ;
  assign n86 = n85 ^ x3 ;
  assign n87 = n83 & n86 ;
  assign n88 = n16 & ~n87 ;
  assign n89 = ~n81 & n88 ;
  assign n90 = ~n61 & ~n89 ;
  assign n91 = x4 & x8 ;
  assign n92 = ~x7 & x8 ;
  assign n93 = ~n91 & ~n92 ;
  assign n94 = x2 & n19 ;
  assign n95 = ~n82 & n94 ;
  assign n96 = ~n93 & n95 ;
  assign n97 = n19 & n21 ;
  assign n98 = x6 & x7 ;
  assign n99 = ~x2 & ~x9 ;
  assign n100 = ~n98 & n99 ;
  assign n101 = ~n92 & n100 ;
  assign n102 = ~n97 & ~n101 ;
  assign n103 = x4 & ~n102 ;
  assign n104 = ~x2 & ~x8 ;
  assign n105 = ~x4 & x6 ;
  assign n106 = n104 & n105 ;
  assign n107 = ~x7 & n106 ;
  assign n108 = ~x0 & ~n107 ;
  assign n109 = ~n103 & n108 ;
  assign n110 = ~n96 & n109 ;
  assign n111 = n110 ^ x7 ;
  assign n112 = x8 & n98 ;
  assign n113 = ~x2 & ~x4 ;
  assign n114 = n112 & n113 ;
  assign n115 = x0 & ~n114 ;
  assign n116 = n115 ^ n111 ;
  assign n117 = n116 ^ n110 ;
  assign n118 = n117 ^ n116 ;
  assign n119 = n25 & n75 ;
  assign n120 = x2 & n119 ;
  assign n121 = n120 ^ n116 ;
  assign n122 = n121 ^ n111 ;
  assign n123 = ~n118 & n122 ;
  assign n124 = n123 ^ n120 ;
  assign n125 = ~x9 & ~n104 ;
  assign n126 = n75 & ~n125 ;
  assign n127 = x2 & ~n91 ;
  assign n128 = ~n19 & n127 ;
  assign n129 = x8 ^ x4 ;
  assign n130 = x9 & n129 ;
  assign n131 = n130 ^ x4 ;
  assign n132 = n128 & n131 ;
  assign n133 = ~n126 & ~n132 ;
  assign n134 = ~n120 & n133 ;
  assign n135 = n134 ^ n111 ;
  assign n136 = ~n124 & ~n135 ;
  assign n137 = n136 ^ n134 ;
  assign n138 = ~n111 & n137 ;
  assign n139 = n138 ^ n123 ;
  assign n140 = n139 ^ x7 ;
  assign n141 = n140 ^ n120 ;
  assign n142 = n141 ^ x3 ;
  assign n143 = n142 ^ n141 ;
  assign n144 = x0 & ~x9 ;
  assign n145 = n24 & n144 ;
  assign n146 = ~x4 & ~x8 ;
  assign n147 = n146 ^ n91 ;
  assign n148 = ~x2 & n147 ;
  assign n149 = n148 ^ n91 ;
  assign n150 = n145 & n149 ;
  assign n151 = x4 ^ x2 ;
  assign n152 = n50 ^ x4 ;
  assign n153 = n152 ^ n50 ;
  assign n156 = n13 ^ x6 ;
  assign n157 = n156 ^ n13 ;
  assign n154 = n13 ^ x9 ;
  assign n155 = n154 ^ n13 ;
  assign n158 = n157 ^ n155 ;
  assign n159 = ~n62 & ~n92 ;
  assign n160 = n159 ^ n13 ;
  assign n161 = n160 ^ n13 ;
  assign n162 = n161 ^ n157 ;
  assign n163 = n157 & ~n162 ;
  assign n164 = n163 ^ n157 ;
  assign n165 = ~n158 & n164 ;
  assign n166 = n165 ^ n163 ;
  assign n167 = n166 ^ n13 ;
  assign n168 = n167 ^ n157 ;
  assign n169 = x0 & n168 ;
  assign n170 = n169 ^ n13 ;
  assign n171 = n170 ^ n50 ;
  assign n172 = n153 & n171 ;
  assign n173 = n172 ^ n50 ;
  assign n174 = ~n151 & n173 ;
  assign n175 = ~n150 & ~n174 ;
  assign n176 = n175 ^ n141 ;
  assign n177 = ~n143 & ~n176 ;
  assign n178 = n177 ^ n141 ;
  assign n179 = ~x1 & ~n178 ;
  assign n180 = n90 & ~n179 ;
  assign n181 = n180 ^ x5 ;
  assign n182 = n181 ^ n180 ;
  assign n183 = ~x1 & ~x4 ;
  assign n184 = ~x0 & n21 ;
  assign n185 = ~n183 & n184 ;
  assign n186 = ~x6 & x9 ;
  assign n187 = ~n129 & n186 ;
  assign n188 = n185 & n187 ;
  assign n265 = x8 ^ x7 ;
  assign n271 = n265 ^ x1 ;
  assign n272 = n271 ^ n265 ;
  assign n266 = x9 ^ x8 ;
  assign n267 = n266 ^ n265 ;
  assign n268 = n267 ^ n40 ;
  assign n269 = n268 ^ x8 ;
  assign n270 = n269 ^ n265 ;
  assign n273 = n272 ^ n270 ;
  assign n276 = n269 ^ x8 ;
  assign n274 = n40 ^ x8 ;
  assign n275 = n274 ^ n270 ;
  assign n277 = n276 ^ n275 ;
  assign n278 = ~n273 & n277 ;
  assign n279 = n278 ^ n269 ;
  assign n280 = n279 ^ n274 ;
  assign n281 = n280 ^ n276 ;
  assign n282 = n275 ^ n272 ;
  assign n283 = n279 & n282 ;
  assign n284 = n283 ^ n269 ;
  assign n285 = n284 ^ n270 ;
  assign n286 = n285 ^ n272 ;
  assign n287 = n281 & ~n286 ;
  assign n288 = n105 & n287 ;
  assign n289 = x0 & n288 ;
  assign n189 = n16 & n94 ;
  assign n190 = n146 & n189 ;
  assign n191 = ~x2 & x8 ;
  assign n192 = x1 & x9 ;
  assign n193 = ~x1 & ~x9 ;
  assign n194 = ~n192 & ~n193 ;
  assign n195 = n75 & ~n194 ;
  assign n196 = n191 & n195 ;
  assign n197 = x6 & n31 ;
  assign n198 = n197 ^ x0 ;
  assign n199 = n198 ^ x0 ;
  assign n200 = x4 ^ x0 ;
  assign n201 = n200 ^ x0 ;
  assign n202 = n199 & ~n201 ;
  assign n203 = n202 ^ x0 ;
  assign n204 = x2 & n203 ;
  assign n205 = n204 ^ x0 ;
  assign n206 = ~n196 & ~n205 ;
  assign n207 = x1 & n19 ;
  assign n208 = n183 & n186 ;
  assign n209 = ~n207 & ~n208 ;
  assign n210 = n104 & ~n209 ;
  assign n211 = x0 & ~n210 ;
  assign n212 = x7 & ~n211 ;
  assign n213 = ~n206 & n212 ;
  assign n214 = ~n190 & ~n213 ;
  assign n215 = x7 & n99 ;
  assign n216 = ~x1 & x8 ;
  assign n217 = n215 & n216 ;
  assign n218 = x1 & ~x6 ;
  assign n219 = ~x8 & n218 ;
  assign n220 = ~x7 & x9 ;
  assign n221 = x2 & x6 ;
  assign n222 = ~x1 & ~x2 ;
  assign n223 = ~n221 & ~n222 ;
  assign n224 = ~n191 & ~n216 ;
  assign n225 = n223 & n224 ;
  assign n226 = n220 & n225 ;
  assign n227 = ~n219 & n226 ;
  assign n228 = ~n217 & ~n227 ;
  assign n229 = n228 ^ x0 ;
  assign n230 = n229 ^ n228 ;
  assign n231 = n197 & n222 ;
  assign n232 = x7 & n221 ;
  assign n233 = n216 & n232 ;
  assign n234 = ~n191 & n218 ;
  assign n235 = ~n159 & n234 ;
  assign n236 = ~n233 & ~n235 ;
  assign n237 = ~x9 & ~n236 ;
  assign n238 = ~n231 & ~n237 ;
  assign n239 = n238 ^ n228 ;
  assign n240 = ~n230 & n239 ;
  assign n241 = n240 ^ n228 ;
  assign n242 = x4 & ~n241 ;
  assign n243 = n214 & ~n242 ;
  assign n290 = n289 ^ n243 ;
  assign n291 = n290 ^ n243 ;
  assign n244 = ~x0 & ~x1 ;
  assign n245 = x2 & ~x4 ;
  assign n246 = n50 & n245 ;
  assign n247 = n99 & n112 ;
  assign n248 = ~n246 & ~n247 ;
  assign n249 = n244 & ~n248 ;
  assign n250 = x6 ^ x1 ;
  assign n251 = n31 ^ x6 ;
  assign n252 = n251 ^ n250 ;
  assign n253 = n146 ^ x4 ;
  assign n254 = ~x6 & n253 ;
  assign n255 = n254 ^ x4 ;
  assign n256 = ~n252 & ~n255 ;
  assign n257 = n256 ^ n254 ;
  assign n258 = n257 ^ x4 ;
  assign n259 = n258 ^ x6 ;
  assign n260 = n250 & n259 ;
  assign n261 = n184 & n260 ;
  assign n262 = ~n249 & ~n261 ;
  assign n263 = n262 ^ n243 ;
  assign n264 = n263 ^ n243 ;
  assign n292 = n291 ^ n264 ;
  assign n293 = n219 & n220 ;
  assign n294 = n21 & n197 ;
  assign n295 = x6 & ~x8 ;
  assign n296 = x2 & x7 ;
  assign n297 = ~n186 & n296 ;
  assign n298 = ~n295 & n297 ;
  assign n299 = ~n294 & ~n298 ;
  assign n300 = ~x1 & ~n299 ;
  assign n301 = ~n293 & ~n300 ;
  assign n302 = x0 & ~n301 ;
  assign n303 = ~n184 & ~n232 ;
  assign n304 = n192 & ~n303 ;
  assign n305 = n11 ^ x7 ;
  assign n306 = n305 ^ x1 ;
  assign n313 = n306 ^ n305 ;
  assign n307 = n306 ^ n99 ;
  assign n308 = n307 ^ n305 ;
  assign n309 = n306 ^ n11 ;
  assign n310 = n309 ^ n99 ;
  assign n311 = n310 ^ n308 ;
  assign n312 = n308 & ~n311 ;
  assign n314 = n313 ^ n312 ;
  assign n315 = n314 ^ n308 ;
  assign n316 = n305 ^ n19 ;
  assign n317 = n312 ^ n308 ;
  assign n318 = ~n316 & n317 ;
  assign n319 = n318 ^ n305 ;
  assign n320 = ~n315 & n319 ;
  assign n321 = n320 ^ n305 ;
  assign n322 = n321 ^ x7 ;
  assign n323 = n322 ^ n305 ;
  assign n324 = ~x0 & n323 ;
  assign n325 = ~n304 & ~n324 ;
  assign n326 = x8 & ~n325 ;
  assign n327 = x7 ^ x2 ;
  assign n328 = n327 ^ n25 ;
  assign n329 = ~n11 & n328 ;
  assign n330 = n329 ^ n11 ;
  assign n331 = n329 ^ n244 ;
  assign n332 = n327 & n331 ;
  assign n333 = n332 ^ n327 ;
  assign n334 = n333 ^ n25 ;
  assign n335 = ~n330 & n334 ;
  assign n336 = ~n326 & ~n335 ;
  assign n337 = ~n302 & n336 ;
  assign n338 = x4 & ~n337 ;
  assign n339 = n338 ^ n243 ;
  assign n340 = n339 ^ n243 ;
  assign n341 = n340 ^ n291 ;
  assign n342 = ~n291 & n341 ;
  assign n343 = n342 ^ n291 ;
  assign n344 = ~n292 & ~n343 ;
  assign n345 = n344 ^ n342 ;
  assign n346 = n345 ^ n243 ;
  assign n347 = n346 ^ n291 ;
  assign n348 = x3 & ~n347 ;
  assign n349 = n348 ^ n243 ;
  assign n350 = ~n188 & n349 ;
  assign n351 = n350 ^ n180 ;
  assign n352 = n182 & ~n351 ;
  assign n353 = n352 ^ n180 ;
  assign n354 = ~n18 & ~n353 ;
  assign y0 = ~n354 ;
endmodule
