module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 ;
  assign n16 = x5 & ~x7 ;
  assign n17 = ~x11 & ~n16 ;
  assign n18 = x9 & x14 ;
  assign n19 = x3 & ~n18 ;
  assign n20 = x14 ^ x13 ;
  assign n21 = n19 & ~n20 ;
  assign n22 = n17 & n21 ;
  assign n23 = x5 & x14 ;
  assign n24 = ~x7 & n23 ;
  assign n25 = x13 & x14 ;
  assign n26 = x9 & ~x11 ;
  assign n27 = ~n25 & n26 ;
  assign n28 = ~n24 & n27 ;
  assign n29 = ~x1 & ~x6 ;
  assign n30 = x1 & x7 ;
  assign n31 = ~x11 & ~x14 ;
  assign n32 = ~x5 & n31 ;
  assign n33 = n30 & n32 ;
  assign n34 = ~x13 & x14 ;
  assign n35 = x5 & ~x9 ;
  assign n36 = n34 & n35 ;
  assign n37 = ~n33 & ~n36 ;
  assign n38 = ~n29 & ~n37 ;
  assign n39 = x3 & n38 ;
  assign n40 = ~n28 & ~n39 ;
  assign n41 = ~n22 & n40 ;
  assign n42 = ~x0 & ~n41 ;
  assign n43 = x9 & ~x14 ;
  assign n44 = x9 & ~x13 ;
  assign n45 = ~n21 & ~n44 ;
  assign n46 = x7 & ~n45 ;
  assign n47 = ~n43 & ~n46 ;
  assign n48 = x6 & ~x11 ;
  assign n49 = ~n47 & n48 ;
  assign n50 = x5 & n49 ;
  assign n51 = ~n42 & ~n50 ;
  assign n52 = x4 & ~n51 ;
  assign n53 = ~x0 & x9 ;
  assign n54 = x8 ^ x6 ;
  assign n55 = n54 ^ x8 ;
  assign n56 = x13 ^ x8 ;
  assign n57 = n55 & n56 ;
  assign n58 = n57 ^ x8 ;
  assign n59 = ~x7 & ~n58 ;
  assign n60 = n59 ^ x6 ;
  assign n61 = n32 & ~n60 ;
  assign n62 = n53 & n61 ;
  assign n63 = ~n52 & ~n62 ;
  assign n64 = x10 & ~n63 ;
  assign n65 = x11 & ~x13 ;
  assign n66 = ~x4 & ~x5 ;
  assign n67 = ~x6 & n66 ;
  assign n68 = ~x9 & ~x14 ;
  assign n69 = x7 & x8 ;
  assign n70 = n68 & n69 ;
  assign n71 = n67 & n70 ;
  assign n72 = x14 & n35 ;
  assign n73 = ~x6 & ~x8 ;
  assign n74 = ~x7 & n66 ;
  assign n75 = ~n73 & n74 ;
  assign n76 = ~n72 & ~n75 ;
  assign n77 = ~x4 & ~x9 ;
  assign n78 = ~x0 & x10 ;
  assign n79 = ~n77 & n78 ;
  assign n80 = ~n76 & n79 ;
  assign n81 = ~n71 & ~n80 ;
  assign n82 = x3 & ~n81 ;
  assign n83 = n65 & n82 ;
  assign n84 = x4 & ~x5 ;
  assign n85 = x7 & ~x11 ;
  assign n86 = n84 & n85 ;
  assign n87 = x10 & ~n86 ;
  assign n88 = x13 & n53 ;
  assign n89 = ~n87 & n88 ;
  assign n90 = ~x10 & ~x13 ;
  assign n91 = n77 & n90 ;
  assign n92 = ~x3 & n91 ;
  assign n93 = ~n89 & ~n92 ;
  assign n94 = x3 & n23 ;
  assign n95 = n94 ^ x9 ;
  assign n96 = n95 ^ n94 ;
  assign n104 = n96 ^ x13 ;
  assign n105 = n94 ^ x1 ;
  assign n106 = ~n104 & n105 ;
  assign n97 = x14 ^ x0 ;
  assign n98 = n97 ^ n96 ;
  assign n99 = n97 ^ x14 ;
  assign n100 = n99 ^ n98 ;
  assign n101 = n98 & n100 ;
  assign n112 = n106 ^ n101 ;
  assign n102 = n101 ^ n96 ;
  assign n103 = n102 ^ n98 ;
  assign n107 = n97 ^ n94 ;
  assign n108 = n107 ^ n106 ;
  assign n109 = n108 ^ n105 ;
  assign n110 = n109 ^ x13 ;
  assign n111 = n103 & n110 ;
  assign n113 = n112 ^ n111 ;
  assign n114 = n113 ^ n107 ;
  assign n115 = n114 ^ n105 ;
  assign n116 = n115 ^ x13 ;
  assign n117 = ~x13 & n116 ;
  assign n118 = n117 ^ x13 ;
  assign n119 = n118 ^ x13 ;
  assign n120 = ~x10 & ~n119 ;
  assign n121 = x11 & n120 ;
  assign n122 = n93 & ~n121 ;
  assign n123 = ~x12 & n122 ;
  assign n124 = ~n83 & n123 ;
  assign n125 = ~n64 & n124 ;
  assign n126 = x8 & ~x11 ;
  assign n127 = ~x7 & n126 ;
  assign n128 = x10 & n25 ;
  assign n129 = n127 & n128 ;
  assign n130 = n67 & n129 ;
  assign n131 = n90 ^ x9 ;
  assign n132 = n131 ^ n90 ;
  assign n133 = n34 & n67 ;
  assign n134 = x7 & ~x8 ;
  assign n135 = ~x11 & n134 ;
  assign n136 = n133 & n135 ;
  assign n137 = x11 ^ x10 ;
  assign n138 = n137 ^ x10 ;
  assign n139 = n138 ^ n136 ;
  assign n140 = x13 & ~x14 ;
  assign n141 = n30 & n84 ;
  assign n142 = n140 & n141 ;
  assign n143 = x5 & ~x13 ;
  assign n144 = ~x2 & n143 ;
  assign n145 = ~n29 & n144 ;
  assign n146 = ~n142 & ~n145 ;
  assign n147 = n146 ^ n78 ;
  assign n148 = ~n146 & ~n147 ;
  assign n149 = n148 ^ x10 ;
  assign n150 = n149 ^ n146 ;
  assign n151 = ~n139 & n150 ;
  assign n152 = n151 ^ n148 ;
  assign n153 = n152 ^ n146 ;
  assign n154 = ~n136 & ~n153 ;
  assign n155 = n154 ^ n136 ;
  assign n156 = n155 ^ n90 ;
  assign n157 = ~n132 & n156 ;
  assign n158 = n157 ^ n90 ;
  assign n159 = ~n130 & ~n158 ;
  assign n160 = x3 & ~n159 ;
  assign n161 = x12 & ~n160 ;
  assign n163 = x11 & n44 ;
  assign n164 = x8 ^ x7 ;
  assign n165 = n164 ^ n44 ;
  assign n166 = n163 ^ n16 ;
  assign n167 = n165 & n166 ;
  assign n168 = n167 ^ n16 ;
  assign n169 = n163 & n168 ;
  assign n170 = n169 ^ n44 ;
  assign n172 = x14 ^ x9 ;
  assign n173 = n172 ^ x7 ;
  assign n171 = x14 ^ x11 ;
  assign n174 = n173 ^ n171 ;
  assign n175 = n174 ^ n173 ;
  assign n176 = n175 ^ x11 ;
  assign n177 = n176 ^ n172 ;
  assign n178 = x6 & n127 ;
  assign n179 = n178 ^ x11 ;
  assign n180 = ~n177 & n179 ;
  assign n181 = n180 ^ n178 ;
  assign n187 = n177 ^ n172 ;
  assign n182 = x6 & ~x13 ;
  assign n183 = n182 ^ n173 ;
  assign n184 = n173 & ~n183 ;
  assign n185 = n184 ^ n173 ;
  assign n186 = n185 ^ n177 ;
  assign n188 = n187 ^ n186 ;
  assign n189 = n183 ^ x11 ;
  assign n190 = n189 ^ n177 ;
  assign n191 = n190 ^ n187 ;
  assign n192 = n190 & n191 ;
  assign n193 = n192 ^ n182 ;
  assign n194 = n193 ^ n187 ;
  assign n195 = ~n188 & ~n194 ;
  assign n196 = n195 ^ n177 ;
  assign n197 = n196 ^ n187 ;
  assign n198 = n181 & ~n197 ;
  assign n199 = n198 ^ n195 ;
  assign n200 = n199 ^ n177 ;
  assign n201 = n200 ^ n187 ;
  assign n202 = n201 ^ x9 ;
  assign n203 = ~n170 & n202 ;
  assign n162 = n65 & n77 ;
  assign n204 = n203 ^ n162 ;
  assign n205 = x10 & ~n204 ;
  assign n206 = n205 ^ n203 ;
  assign n207 = n161 & n206 ;
  assign n208 = ~n125 & ~n207 ;
  assign n209 = ~x10 & ~x11 ;
  assign n210 = ~n43 & ~n53 ;
  assign n211 = ~x7 & ~x8 ;
  assign n212 = n182 & ~n211 ;
  assign n213 = n66 & n212 ;
  assign n214 = ~n210 & n213 ;
  assign n215 = n214 ^ x3 ;
  assign n216 = n215 ^ n214 ;
  assign n217 = n214 ^ n68 ;
  assign n218 = ~n216 & n217 ;
  assign n219 = n218 ^ n214 ;
  assign n220 = n209 & n219 ;
  assign n221 = ~n208 & ~n220 ;
  assign y0 = ~n221 ;
endmodule
