// Benchmark "./pla/p1.pla_dbb_orig_4NonExact" written by ABC on Fri Nov 20 10:27:46 2020

module \./pla/p1.pla_dbb_orig_4NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = 1'b1;
endmodule


