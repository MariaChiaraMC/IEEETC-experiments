module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n9 = x2 & ~x5 ;
  assign n10 = ~x6 & n9 ;
  assign n11 = x2 & ~x3 ;
  assign n12 = x4 & ~n11 ;
  assign n13 = ~n10 & n12 ;
  assign n14 = x6 ^ x5 ;
  assign n15 = n14 ^ x7 ;
  assign n16 = ~x3 & n15 ;
  assign n17 = n13 & ~n16 ;
  assign n18 = x5 ^ x3 ;
  assign n19 = x7 ^ x5 ;
  assign n20 = x3 ^ x2 ;
  assign n21 = n20 ^ x3 ;
  assign n22 = n21 ^ x7 ;
  assign n23 = ~x7 & n22 ;
  assign n24 = n23 ^ x7 ;
  assign n25 = ~n19 & ~n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n26 ^ x7 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = n18 & n28 ;
  assign n30 = n29 ^ n20 ;
  assign n31 = ~x4 & n30 ;
  assign n32 = ~x0 & ~n31 ;
  assign n33 = ~x1 & n32 ;
  assign n34 = ~n17 & n33 ;
  assign y0 = n34 ;
endmodule
