module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n19 = ~x13 & ~x15 ;
  assign n18 = x12 ^ x11 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = n20 ^ x12 ;
  assign n22 = n19 ^ x14 ;
  assign n23 = n22 ^ x14 ;
  assign n24 = x1 & ~x3 ;
  assign n25 = x4 & x5 ;
  assign n26 = n24 & n25 ;
  assign n27 = ~x14 & n26 ;
  assign n28 = n27 ^ x14 ;
  assign n29 = n23 & n28 ;
  assign n30 = n29 ^ x14 ;
  assign n31 = n30 ^ n20 ;
  assign n32 = ~n21 & n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ x14 ;
  assign n35 = n34 ^ x12 ;
  assign n36 = n20 & ~n35 ;
  assign n37 = n36 ^ n20 ;
  assign n38 = n37 ^ n18 ;
  assign y0 = n38 ;
endmodule
