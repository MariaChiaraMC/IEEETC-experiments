module top( x0 , x1 , x2 , x3 , x4 , y0 );
  input x0 , x1 , x2 , x3 , x4 ;
  output y0 ;
  wire n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n6 = x4 ^ x1 ;
  assign n7 = n6 ^ x2 ;
  assign n8 = n7 ^ n6 ;
  assign n9 = n8 ^ x0 ;
  assign n10 = n9 ^ x0 ;
  assign n11 = x4 ^ x0 ;
  assign n12 = n11 ^ n6 ;
  assign n13 = n12 ^ x3 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n14 ^ x0 ;
  assign n16 = n15 ^ n10 ;
  assign n20 = n10 ^ n9 ;
  assign n21 = n6 & ~n20 ;
  assign n17 = n12 ^ n6 ;
  assign n18 = n17 ^ n6 ;
  assign n19 = ~n9 & n18 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ n6 ;
  assign n24 = n23 ^ n17 ;
  assign n25 = n16 & n24 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = n10 & n26 ;
  assign n28 = n27 ^ n19 ;
  assign n29 = n28 ^ n25 ;
  assign y0 = n29 ;
endmodule
