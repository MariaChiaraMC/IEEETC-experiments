module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 ;
  assign n79 = ~x1 & ~x2 ;
  assign n83 = x0 & ~x3 ;
  assign n9 = x5 & ~x7 ;
  assign n80 = ~x3 & ~n9 ;
  assign n81 = n80 ^ x6 ;
  assign n82 = n81 ^ n80 ;
  assign n84 = n83 ^ n82 ;
  assign n85 = n84 ^ n83 ;
  assign n20 = x5 & x7 ;
  assign n26 = x0 & x7 ;
  assign n86 = ~n26 & ~n83 ;
  assign n87 = ~n20 & n86 ;
  assign n88 = n85 ^ n81 ;
  assign n89 = n88 ^ n85 ;
  assign n90 = ~n87 & ~n89 ;
  assign n91 = n90 ^ n83 ;
  assign n92 = ~x5 & x7 ;
  assign n93 = n92 ^ n83 ;
  assign n94 = ~n88 & n93 ;
  assign n95 = n94 ^ n85 ;
  assign n96 = n95 ^ n88 ;
  assign n97 = ~n91 & ~n96 ;
  assign n98 = n85 & n97 ;
  assign n99 = n98 ^ n90 ;
  assign n100 = n79 & n99 ;
  assign n101 = x5 ^ x3 ;
  assign n102 = ~x3 & ~x6 ;
  assign n103 = x0 & ~n102 ;
  assign n104 = ~x7 & n103 ;
  assign n105 = ~x2 & ~x3 ;
  assign n106 = x6 & ~n105 ;
  assign n107 = n104 & ~n106 ;
  assign n108 = n107 ^ n101 ;
  assign n109 = n108 ^ x5 ;
  assign n110 = n109 ^ n108 ;
  assign n111 = x2 & x6 ;
  assign n112 = n9 & n111 ;
  assign n113 = n112 ^ n108 ;
  assign n114 = n113 ^ n101 ;
  assign n115 = ~n110 & ~n114 ;
  assign n116 = n115 ^ n112 ;
  assign n14 = ~x0 & ~x6 ;
  assign n117 = ~x2 & n14 ;
  assign n118 = ~n112 & ~n117 ;
  assign n119 = n118 ^ n101 ;
  assign n120 = ~n116 & n119 ;
  assign n121 = n120 ^ n118 ;
  assign n122 = n101 & n121 ;
  assign n123 = n122 ^ n115 ;
  assign n124 = n123 ^ x3 ;
  assign n125 = n124 ^ n112 ;
  assign n126 = x1 & ~n125 ;
  assign n127 = ~x1 & x2 ;
  assign n128 = x5 & n127 ;
  assign n129 = n104 & n128 ;
  assign n130 = ~n126 & ~n129 ;
  assign n131 = ~n100 & n130 ;
  assign n10 = x2 & ~x6 ;
  assign n11 = ~x0 & x1 ;
  assign n12 = n10 & n11 ;
  assign n13 = n9 & n12 ;
  assign n15 = x2 & ~x5 ;
  assign n16 = n14 & ~n15 ;
  assign n17 = ~x5 & ~x7 ;
  assign n18 = x2 ^ x1 ;
  assign n19 = n18 ^ x2 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = n19 & ~n21 ;
  assign n23 = n22 ^ x2 ;
  assign n24 = ~n17 & ~n23 ;
  assign n25 = n16 & ~n24 ;
  assign n27 = ~x2 & x5 ;
  assign n28 = x1 & n27 ;
  assign n29 = ~x1 & ~x6 ;
  assign n30 = n15 & n29 ;
  assign n31 = ~n28 & ~n30 ;
  assign n32 = n26 & ~n31 ;
  assign n33 = x1 & ~x6 ;
  assign n34 = ~x2 & n17 ;
  assign n35 = n33 & n34 ;
  assign n36 = ~n32 & ~n35 ;
  assign n37 = x1 ^ x0 ;
  assign n38 = n37 ^ n18 ;
  assign n39 = x5 ^ x2 ;
  assign n40 = n39 ^ x5 ;
  assign n41 = n20 ^ x5 ;
  assign n42 = n40 & ~n41 ;
  assign n43 = n42 ^ x5 ;
  assign n44 = n43 ^ n18 ;
  assign n45 = ~n38 & n44 ;
  assign n46 = n45 ^ n42 ;
  assign n47 = n46 ^ x5 ;
  assign n48 = n47 ^ n37 ;
  assign n49 = ~n18 & ~n48 ;
  assign n50 = n49 ^ n18 ;
  assign n51 = x6 & ~n50 ;
  assign n52 = n36 & ~n51 ;
  assign n53 = ~n25 & n52 ;
  assign n54 = ~x3 & ~n53 ;
  assign n55 = ~x7 & n30 ;
  assign n56 = n55 ^ x3 ;
  assign n57 = n56 ^ n55 ;
  assign n58 = x7 ^ x5 ;
  assign n61 = n39 ^ x6 ;
  assign n59 = n39 ^ x1 ;
  assign n60 = n59 ^ x7 ;
  assign n62 = n61 ^ n60 ;
  assign n63 = n62 ^ n58 ;
  assign n64 = n58 & ~n63 ;
  assign n65 = n64 ^ n39 ;
  assign n66 = n65 ^ n58 ;
  assign n67 = n59 & ~n61 ;
  assign n68 = n67 ^ n39 ;
  assign n69 = n66 & n68 ;
  assign n70 = n69 ^ n39 ;
  assign n71 = n70 ^ n55 ;
  assign n72 = n71 ^ n55 ;
  assign n73 = n57 & n72 ;
  assign n74 = n73 ^ n55 ;
  assign n75 = x0 & n74 ;
  assign n76 = n75 ^ n55 ;
  assign n77 = ~n54 & ~n76 ;
  assign n78 = ~n13 & n77 ;
  assign n132 = n131 ^ n78 ;
  assign n133 = n132 ^ n78 ;
  assign n134 = ~x0 & ~x5 ;
  assign n135 = n105 & n134 ;
  assign n136 = n135 ^ x6 ;
  assign n137 = n136 ^ x3 ;
  assign n138 = n137 ^ n136 ;
  assign n139 = n138 ^ x6 ;
  assign n140 = n139 ^ x6 ;
  assign n141 = n137 ^ n28 ;
  assign n142 = n141 ^ n136 ;
  assign n143 = n142 ^ x6 ;
  assign n144 = ~n140 & ~n143 ;
  assign n145 = n144 ^ n136 ;
  assign n146 = n145 ^ x6 ;
  assign n147 = n146 ^ n139 ;
  assign n148 = n136 ^ x0 ;
  assign n149 = n148 ^ x6 ;
  assign n150 = ~x0 & ~n149 ;
  assign n151 = n142 ^ x0 ;
  assign n152 = n151 ^ x6 ;
  assign n153 = n152 ^ n139 ;
  assign n154 = ~n128 & n153 ;
  assign n155 = n154 ^ n128 ;
  assign n156 = n155 ^ x0 ;
  assign n157 = n156 ^ x6 ;
  assign n158 = n157 ^ n139 ;
  assign n159 = n150 & ~n158 ;
  assign n160 = n159 ^ x6 ;
  assign n161 = n147 & ~n160 ;
  assign n162 = n161 ^ n159 ;
  assign n163 = n162 ^ n136 ;
  assign n164 = n163 ^ x6 ;
  assign n165 = n164 ^ n135 ;
  assign n166 = n165 ^ n136 ;
  assign n167 = x7 & ~n166 ;
  assign n168 = n167 ^ n78 ;
  assign n169 = n168 ^ n78 ;
  assign n170 = n133 & ~n169 ;
  assign n171 = n170 ^ n78 ;
  assign n172 = ~x4 & n171 ;
  assign n173 = n172 ^ n78 ;
  assign y0 = ~n173 ;
endmodule
