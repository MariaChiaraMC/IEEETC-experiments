module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 ;
  assign n17 = ~x3 & ~x4 ;
  assign n18 = ~x5 & x7 ;
  assign n19 = x7 & x9 ;
  assign n20 = x10 & n19 ;
  assign n21 = ~x12 & ~n20 ;
  assign n22 = x13 & x15 ;
  assign n23 = ~x8 & ~x11 ;
  assign n24 = ~n22 & n23 ;
  assign n25 = ~x9 & ~x10 ;
  assign n26 = x5 & ~x6 ;
  assign n27 = ~x13 & ~x15 ;
  assign n28 = n27 ^ x14 ;
  assign n29 = ~n26 & ~n28 ;
  assign n30 = ~n25 & n29 ;
  assign n31 = n24 & n30 ;
  assign n32 = n21 & n31 ;
  assign n33 = ~n18 & ~n32 ;
  assign n34 = ~x0 & ~x2 ;
  assign n35 = ~n33 & n34 ;
  assign n36 = n35 ^ x1 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = n35 ^ x0 ;
  assign n39 = ~n37 & n38 ;
  assign n40 = n39 ^ n35 ;
  assign n41 = n17 & n40 ;
  assign y0 = n41 ;
endmodule
