module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 ;
  assign n18 = ~x2 & x4 ;
  assign n19 = x0 & ~x1 ;
  assign n20 = x3 & n19 ;
  assign n21 = ~x10 & n20 ;
  assign n22 = ~x13 & ~n21 ;
  assign n23 = ~n18 & ~n22 ;
  assign n26 = x3 ^ x0 ;
  assign n27 = n26 ^ x3 ;
  assign n24 = x3 ^ x2 ;
  assign n25 = n24 ^ x3 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = x1 & ~x10 ;
  assign n30 = n29 ^ x3 ;
  assign n31 = n30 ^ x3 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = ~n27 & ~n32 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = n28 & ~n34 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = n36 ^ x3 ;
  assign n38 = n37 ^ n27 ;
  assign n39 = ~x13 & ~n38 ;
  assign n40 = n39 ^ x3 ;
  assign n41 = ~n23 & ~n40 ;
  assign n42 = ~x9 & ~n41 ;
  assign n43 = ~x2 & ~x3 ;
  assign n44 = n19 & ~n43 ;
  assign n45 = x14 & ~n44 ;
  assign n46 = ~x13 & ~n45 ;
  assign n47 = x10 & ~n46 ;
  assign n48 = ~n42 & ~n47 ;
  assign n16 = x9 & x10 ;
  assign n17 = ~x13 & n16 ;
  assign n49 = n48 ^ n17 ;
  assign n50 = n17 ^ x14 ;
  assign n51 = n17 ^ x11 ;
  assign n52 = n17 & ~n51 ;
  assign n53 = n52 ^ n17 ;
  assign n54 = ~n50 & n53 ;
  assign n55 = n54 ^ n52 ;
  assign n56 = n55 ^ n17 ;
  assign n57 = n56 ^ x11 ;
  assign n58 = ~n49 & ~n57 ;
  assign n59 = n58 ^ n17 ;
  assign y0 = n59 ;
endmodule
