module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 ;
  assign n9 = x6 ^ x5 ;
  assign n10 = x7 ^ x6 ;
  assign n11 = ~n9 & ~n10 ;
  assign n12 = n11 ^ x4 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n13 ^ x3 ;
  assign n15 = ~x5 & ~x6 ;
  assign n16 = n15 ^ x2 ;
  assign n17 = ~n15 & n16 ;
  assign n18 = n17 ^ n11 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = ~n14 & ~n19 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n21 ^ n15 ;
  assign n23 = ~x3 & ~n22 ;
  assign n24 = n23 ^ x3 ;
  assign n25 = n24 ^ x2 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = ~x7 & ~n15 ;
  assign n28 = x5 & x6 ;
  assign n29 = ~x3 & x4 ;
  assign n30 = ~n28 & n29 ;
  assign n31 = ~n27 & n30 ;
  assign n32 = n31 ^ n25 ;
  assign n33 = n26 & ~n32 ;
  assign n34 = n33 ^ n25 ;
  assign n35 = x4 & ~x5 ;
  assign n36 = ~n25 & ~n35 ;
  assign n37 = n36 ^ x1 ;
  assign n38 = ~n34 & ~n37 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = ~x1 & n39 ;
  assign n41 = n40 ^ x2 ;
  assign n42 = n41 ^ x1 ;
  assign y0 = n42 ;
endmodule
