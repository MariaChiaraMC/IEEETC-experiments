// Benchmark "./newxcpla1.pla" written by ABC on Thu Apr 23 10:59:58 2020

module \./newxcpla1.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8,
    z10  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8;
  output z10;
  assign z10 = ~x0 | x2;
endmodule


