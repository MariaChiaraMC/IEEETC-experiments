module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 ;
  assign n9 = x2 & x3 ;
  assign n10 = n9 ^ x5 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = ~x0 & ~x7 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = n13 ^ n9 ;
  assign n15 = n11 & n14 ;
  assign n16 = n15 ^ n9 ;
  assign n17 = x6 & n16 ;
  assign n18 = n17 ^ n9 ;
  assign n19 = ~x1 & n18 ;
  assign n20 = ~x2 & ~x3 ;
  assign n21 = x1 & ~x3 ;
  assign n22 = ~n20 & ~n21 ;
  assign n23 = ~x6 & n12 ;
  assign n24 = n22 & n23 ;
  assign n25 = x6 & x7 ;
  assign n26 = n25 ^ x1 ;
  assign n27 = n26 ^ x1 ;
  assign n28 = ~x0 & x3 ;
  assign n29 = n28 ^ x1 ;
  assign n30 = n27 & n29 ;
  assign n31 = n30 ^ x1 ;
  assign n32 = ~x2 & n31 ;
  assign n33 = ~n24 & ~n32 ;
  assign n34 = ~x5 & ~n33 ;
  assign n42 = x7 ^ x6 ;
  assign n36 = x7 ^ x1 ;
  assign n43 = n42 ^ n36 ;
  assign n44 = n43 ^ n36 ;
  assign n38 = x5 ^ x2 ;
  assign n35 = x7 ^ x5 ;
  assign n37 = n36 ^ n35 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = n39 ^ x7 ;
  assign n41 = n40 ^ n36 ;
  assign n45 = n44 ^ n41 ;
  assign n48 = n40 ^ x7 ;
  assign n46 = n38 ^ x7 ;
  assign n47 = n46 ^ n41 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = n45 & n49 ;
  assign n51 = n50 ^ n40 ;
  assign n52 = n51 ^ n46 ;
  assign n53 = n52 ^ n48 ;
  assign n54 = n47 ^ n44 ;
  assign n55 = ~n51 & n54 ;
  assign n56 = n55 ^ n40 ;
  assign n57 = n56 ^ n41 ;
  assign n58 = n57 ^ n44 ;
  assign n59 = n53 & ~n58 ;
  assign n60 = ~x0 & ~n59 ;
  assign n61 = x5 & x6 ;
  assign n62 = ~x0 & x6 ;
  assign n63 = ~n61 & ~n62 ;
  assign n64 = x2 & n63 ;
  assign n65 = ~n60 & ~n64 ;
  assign n66 = ~x3 & n65 ;
  assign n67 = ~n34 & ~n66 ;
  assign n68 = ~n19 & n67 ;
  assign n69 = x4 & ~n68 ;
  assign n70 = x5 & x7 ;
  assign n71 = n20 & n70 ;
  assign n72 = x0 & n71 ;
  assign n84 = ~x2 & x6 ;
  assign n85 = n28 & ~n84 ;
  assign n86 = ~x5 & ~x7 ;
  assign n87 = ~x6 & ~n86 ;
  assign n88 = n85 & ~n87 ;
  assign n89 = ~x4 & ~n88 ;
  assign n90 = x3 ^ x0 ;
  assign n91 = n61 ^ x3 ;
  assign n92 = n91 ^ n61 ;
  assign n93 = ~x7 & ~n84 ;
  assign n94 = n93 ^ n61 ;
  assign n95 = ~n92 & n94 ;
  assign n96 = n95 ^ n61 ;
  assign n97 = ~n90 & ~n96 ;
  assign n98 = n97 ^ x0 ;
  assign n99 = n89 & ~n98 ;
  assign n100 = x0 & n9 ;
  assign n101 = ~x7 & n61 ;
  assign n102 = n20 & n101 ;
  assign n103 = ~n100 & ~n102 ;
  assign n104 = ~n99 & n103 ;
  assign n73 = ~x2 & ~n25 ;
  assign n75 = n73 ^ x6 ;
  assign n74 = n73 ^ n62 ;
  assign n76 = n75 ^ n74 ;
  assign n77 = n75 ^ x3 ;
  assign n78 = n77 ^ n75 ;
  assign n79 = ~n76 & n78 ;
  assign n80 = n79 ^ n75 ;
  assign n81 = ~x5 & ~n80 ;
  assign n82 = n81 ^ n73 ;
  assign n83 = ~x4 & ~n82 ;
  assign n105 = n104 ^ n83 ;
  assign n106 = n105 ^ n104 ;
  assign n107 = n104 ^ x0 ;
  assign n108 = n107 ^ n9 ;
  assign n109 = n108 ^ n104 ;
  assign n110 = ~n106 & ~n109 ;
  assign n111 = n110 ^ n104 ;
  assign n112 = x1 & n111 ;
  assign n113 = n112 ^ n104 ;
  assign n114 = ~n72 & n113 ;
  assign n115 = ~n69 & n114 ;
  assign y0 = ~n115 ;
endmodule
