// Benchmark "./bench.pla" written by ABC on Thu Apr 23 10:59:48 2020

module \./bench.pla  ( 
    x0, x1, x2, x3, x4, x5,
    z4  );
  input  x0, x1, x2, x3, x4, x5;
  output z4;
  assign z4 = ~x1 | ~x3;
endmodule


