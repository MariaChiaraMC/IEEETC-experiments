module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 ;
  assign n13 = x7 ^ x4 ;
  assign n9 = x4 ^ x3 ;
  assign n10 = n9 ^ x5 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = n11 ^ x4 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n9 ^ x7 ;
  assign n16 = n15 ^ x4 ;
  assign n17 = n16 ^ x4 ;
  assign n18 = ~n11 & ~n17 ;
  assign n19 = n18 ^ n11 ;
  assign n20 = n16 & ~n19 ;
  assign n21 = n20 ^ x4 ;
  assign n22 = n14 & ~n21 ;
  assign n23 = n22 ^ n18 ;
  assign n24 = n23 ^ x4 ;
  assign n25 = n24 ^ x3 ;
  assign n26 = n25 ^ n13 ;
  assign n27 = ~x2 & ~n26 ;
  assign n28 = ~x3 & ~x5 ;
  assign n29 = x4 & n28 ;
  assign n30 = ~x4 & x5 ;
  assign n31 = n30 ^ x7 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = x2 & ~x5 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = ~n32 & n34 ;
  assign n36 = n35 ^ n30 ;
  assign n37 = ~n29 & ~n36 ;
  assign n38 = ~x1 & ~n37 ;
  assign n39 = ~n27 & ~n38 ;
  assign n40 = ~x6 & ~n39 ;
  assign n41 = x5 & x6 ;
  assign n42 = ~x2 & n41 ;
  assign n43 = x4 & ~n42 ;
  assign n44 = ~x1 & ~n43 ;
  assign n45 = ~x4 & ~n28 ;
  assign n46 = n45 ^ n41 ;
  assign n47 = n46 ^ n45 ;
  assign n48 = n45 ^ x3 ;
  assign n49 = n48 ^ n45 ;
  assign n50 = ~n47 & ~n49 ;
  assign n51 = n50 ^ n45 ;
  assign n52 = x2 & n51 ;
  assign n53 = n52 ^ n45 ;
  assign n54 = n44 & ~n53 ;
  assign n55 = ~x3 & ~x7 ;
  assign n56 = x1 & ~x4 ;
  assign n57 = ~n55 & ~n56 ;
  assign n58 = n42 & ~n57 ;
  assign n59 = x5 ^ x4 ;
  assign n60 = x7 ^ x5 ;
  assign n61 = x7 ^ x3 ;
  assign n62 = ~x7 & ~n61 ;
  assign n63 = n62 ^ x7 ;
  assign n64 = ~n60 & ~n63 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = n65 ^ x7 ;
  assign n67 = n66 ^ x3 ;
  assign n68 = ~n59 & ~n67 ;
  assign n69 = n68 ^ x4 ;
  assign n70 = x1 & n69 ;
  assign n71 = ~x2 & n70 ;
  assign n72 = ~n58 & ~n71 ;
  assign n73 = ~n54 & n72 ;
  assign n74 = ~n40 & n73 ;
  assign n75 = ~x0 & ~n74 ;
  assign y0 = n75 ;
endmodule
