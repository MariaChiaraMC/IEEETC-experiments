module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n18 = x12 ^ x0 ;
  assign n19 = x3 & x6 ;
  assign n20 = x1 & n19 ;
  assign n21 = ~x14 & ~n20 ;
  assign n22 = ~x15 & ~x16 ;
  assign n23 = ~n21 & n22 ;
  assign n24 = ~x13 & n23 ;
  assign n25 = n24 ^ x11 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = x13 & ~x14 ;
  assign n28 = n27 ^ n24 ;
  assign n29 = n26 & n28 ;
  assign n30 = n29 ^ n24 ;
  assign n31 = n30 ^ x12 ;
  assign n32 = n18 & ~n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ n24 ;
  assign n35 = n34 ^ x0 ;
  assign n36 = ~x12 & ~n35 ;
  assign n37 = n36 ^ x12 ;
  assign y0 = ~n37 ;
endmodule
