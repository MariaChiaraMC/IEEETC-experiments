module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 ;
  assign n25 = x1 ^ x0 ;
  assign n26 = x2 ^ x1 ;
  assign n27 = n26 ^ x5 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = x5 ^ x3 ;
  assign n30 = x5 ^ x1 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = ~n29 & ~n31 ;
  assign n33 = n32 ^ x5 ;
  assign n34 = n33 ^ n29 ;
  assign n35 = n28 & ~n34 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ n29 ;
  assign n38 = n25 & ~n37 ;
  assign n39 = ~x4 & n38 ;
  assign n40 = ~x20 & ~x21 ;
  assign n41 = n40 ^ x19 ;
  assign n42 = n41 ^ x19 ;
  assign n43 = ~x8 & ~x9 ;
  assign n44 = x10 & ~x11 ;
  assign n45 = n43 & n44 ;
  assign n46 = x12 & x16 ;
  assign n47 = x0 & x1 ;
  assign n48 = x6 & x13 ;
  assign n49 = n47 & n48 ;
  assign n50 = n46 & n49 ;
  assign n51 = n45 & n50 ;
  assign n52 = x7 & n51 ;
  assign n53 = x12 & n44 ;
  assign n54 = x8 & n53 ;
  assign n55 = x13 & ~n54 ;
  assign n56 = x7 & ~n55 ;
  assign n57 = x13 ^ x11 ;
  assign n58 = x16 ^ x13 ;
  assign n59 = n58 ^ x16 ;
  assign n60 = n59 ^ n57 ;
  assign n61 = n46 ^ x6 ;
  assign n62 = x6 & n61 ;
  assign n63 = n62 ^ x16 ;
  assign n64 = n63 ^ x6 ;
  assign n65 = n60 & ~n64 ;
  assign n66 = n65 ^ n62 ;
  assign n67 = n66 ^ x6 ;
  assign n68 = n57 & n67 ;
  assign n69 = n68 ^ x13 ;
  assign n70 = x10 & ~n69 ;
  assign n71 = ~n56 & ~n70 ;
  assign n72 = ~x9 & ~n71 ;
  assign n73 = x9 & x10 ;
  assign n74 = n73 ^ x12 ;
  assign n75 = n74 ^ x13 ;
  assign n76 = ~x9 & ~x10 ;
  assign n77 = n76 ^ x7 ;
  assign n78 = x12 & ~n77 ;
  assign n79 = n78 ^ n76 ;
  assign n80 = ~n75 & ~n79 ;
  assign n81 = n80 ^ n78 ;
  assign n82 = n81 ^ n76 ;
  assign n83 = n82 ^ x12 ;
  assign n84 = x13 & ~n83 ;
  assign n85 = ~x11 & ~n84 ;
  assign n86 = ~x8 & n85 ;
  assign n87 = x7 & ~x10 ;
  assign n88 = n87 ^ x16 ;
  assign n89 = n87 ^ x13 ;
  assign n90 = n89 ^ x13 ;
  assign n91 = n90 ^ n88 ;
  assign n92 = x12 ^ x6 ;
  assign n93 = x6 & ~n92 ;
  assign n94 = n93 ^ x13 ;
  assign n95 = n94 ^ x6 ;
  assign n96 = ~n91 & ~n95 ;
  assign n97 = n96 ^ n93 ;
  assign n98 = n97 ^ x6 ;
  assign n99 = ~n88 & n98 ;
  assign n100 = n99 ^ n87 ;
  assign n101 = n43 & n100 ;
  assign n102 = x6 & ~x7 ;
  assign n103 = x15 ^ x13 ;
  assign n104 = n103 ^ x15 ;
  assign n105 = x8 & n87 ;
  assign n106 = ~x12 & ~n105 ;
  assign n107 = n106 ^ x15 ;
  assign n108 = ~n104 & ~n107 ;
  assign n109 = n108 ^ x15 ;
  assign n110 = x15 & ~n43 ;
  assign n111 = n110 ^ n102 ;
  assign n112 = n109 & ~n111 ;
  assign n113 = n112 ^ n110 ;
  assign n114 = ~n102 & n113 ;
  assign n115 = n114 ^ n102 ;
  assign n116 = ~n101 & ~n115 ;
  assign n117 = ~n86 & n116 ;
  assign n118 = ~n72 & n117 ;
  assign n119 = ~x17 & ~n118 ;
  assign n120 = x11 & ~x12 ;
  assign n121 = ~x6 & ~x7 ;
  assign n122 = x17 & n121 ;
  assign n123 = ~x13 & ~x18 ;
  assign n124 = ~x15 & ~n123 ;
  assign n125 = ~x10 & n43 ;
  assign n126 = x16 & n125 ;
  assign n127 = ~n124 & n126 ;
  assign n128 = n122 & n127 ;
  assign n129 = n120 & n128 ;
  assign n130 = ~x0 & ~n129 ;
  assign n131 = ~n119 & n130 ;
  assign n132 = x2 & ~n131 ;
  assign n133 = ~x2 & n73 ;
  assign n134 = x13 & n126 ;
  assign n135 = ~n133 & ~n134 ;
  assign n136 = n120 & ~n135 ;
  assign n137 = ~x0 & ~x1 ;
  assign n138 = ~x13 & n47 ;
  assign n139 = ~n137 & ~n138 ;
  assign n140 = ~n136 & ~n139 ;
  assign n141 = x15 & ~n140 ;
  assign n142 = x4 & ~n141 ;
  assign n143 = ~n132 & n142 ;
  assign n144 = ~n52 & n143 ;
  assign n145 = ~x3 & ~n144 ;
  assign n165 = ~x12 & ~x13 ;
  assign n166 = ~x4 & n165 ;
  assign n167 = x9 & n166 ;
  assign n168 = n44 & n167 ;
  assign n146 = x11 & n76 ;
  assign n147 = x13 & n146 ;
  assign n148 = n76 ^ x11 ;
  assign n149 = ~x2 & ~x15 ;
  assign n150 = n149 ^ n76 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = n151 ^ n148 ;
  assign n153 = ~x2 & ~x9 ;
  assign n154 = n153 ^ x13 ;
  assign n155 = ~x13 & n154 ;
  assign n156 = n155 ^ n149 ;
  assign n157 = n156 ^ x13 ;
  assign n158 = n152 & n157 ;
  assign n159 = n158 ^ n155 ;
  assign n160 = n159 ^ x13 ;
  assign n161 = ~n148 & ~n160 ;
  assign n162 = n121 & n161 ;
  assign n163 = ~x12 & n162 ;
  assign n164 = ~n147 & ~n163 ;
  assign n169 = n168 ^ n164 ;
  assign n170 = n164 ^ x4 ;
  assign n171 = n164 ^ x8 ;
  assign n172 = ~n164 & n171 ;
  assign n173 = n172 ^ n164 ;
  assign n174 = ~n170 & ~n173 ;
  assign n175 = n174 ^ n172 ;
  assign n176 = n175 ^ n164 ;
  assign n177 = n176 ^ x8 ;
  assign n178 = ~n169 & n177 ;
  assign n179 = n178 ^ n168 ;
  assign n180 = ~x0 & ~x15 ;
  assign n181 = x3 & ~n180 ;
  assign n182 = x4 & ~n181 ;
  assign n183 = x1 & ~n167 ;
  assign n184 = ~n182 & ~n183 ;
  assign n185 = n184 ^ x1 ;
  assign n186 = ~x2 & n185 ;
  assign n187 = n186 ^ x1 ;
  assign n188 = ~n179 & ~n187 ;
  assign n189 = ~n145 & n188 ;
  assign n190 = x5 & ~n189 ;
  assign n191 = x2 & ~n137 ;
  assign n192 = x15 & x17 ;
  assign n193 = ~x0 & ~x8 ;
  assign n194 = n73 & n193 ;
  assign n195 = ~n192 & n194 ;
  assign n196 = n191 & ~n195 ;
  assign n211 = ~x11 & n121 ;
  assign n212 = n166 & n211 ;
  assign n197 = n180 ^ n121 ;
  assign n198 = x11 ^ x10 ;
  assign n199 = n198 ^ n180 ;
  assign n200 = ~n180 & ~n199 ;
  assign n201 = n200 ^ n180 ;
  assign n202 = ~n197 & ~n201 ;
  assign n203 = n202 ^ n200 ;
  assign n204 = n203 ^ n180 ;
  assign n205 = n204 ^ n198 ;
  assign n206 = x11 & ~n205 ;
  assign n207 = n206 ^ n198 ;
  assign n208 = n167 & n207 ;
  assign n213 = n212 ^ n208 ;
  assign n209 = ~x1 & x11 ;
  assign n210 = n209 ^ n208 ;
  assign n214 = n213 ^ n210 ;
  assign n215 = n213 ^ n76 ;
  assign n216 = n215 ^ n213 ;
  assign n217 = n214 & n216 ;
  assign n218 = n217 ^ n213 ;
  assign n219 = ~x8 & n218 ;
  assign n220 = n219 ^ n208 ;
  assign n221 = n196 & n220 ;
  assign n222 = ~x0 & ~x2 ;
  assign n223 = x22 & x23 ;
  assign n224 = ~x15 & n223 ;
  assign n225 = ~x4 & ~n224 ;
  assign n226 = x13 ^ x12 ;
  assign n231 = x13 ^ x8 ;
  assign n232 = ~x10 & n231 ;
  assign n227 = x13 ^ x9 ;
  assign n228 = n227 ^ x13 ;
  assign n229 = n57 & n228 ;
  assign n236 = n232 ^ n229 ;
  assign n230 = n229 ^ n226 ;
  assign n233 = n232 ^ x13 ;
  assign n234 = n233 ^ n226 ;
  assign n235 = ~n230 & n234 ;
  assign n237 = n236 ^ n235 ;
  assign n238 = ~n226 & n237 ;
  assign n239 = n238 ^ n226 ;
  assign n240 = n239 ^ x12 ;
  assign n241 = x5 & n240 ;
  assign n242 = ~x1 & n241 ;
  assign n243 = ~n225 & ~n242 ;
  assign n244 = n222 & ~n243 ;
  assign n245 = ~n221 & ~n244 ;
  assign n246 = ~x3 & ~n245 ;
  assign n270 = x0 & ~x1 ;
  assign n271 = ~x5 & n270 ;
  assign n272 = x3 & ~x5 ;
  assign n273 = x1 & n272 ;
  assign n263 = x1 & x2 ;
  assign n274 = ~x0 & n263 ;
  assign n275 = ~n273 & ~n274 ;
  assign n276 = ~n271 & n275 ;
  assign n247 = ~x9 & ~n193 ;
  assign n248 = x3 & ~n47 ;
  assign n249 = ~n247 & n248 ;
  assign n250 = x8 & ~x11 ;
  assign n251 = ~n121 & ~n250 ;
  assign n252 = n165 & ~n251 ;
  assign n253 = n249 & n252 ;
  assign n254 = x9 & ~n250 ;
  assign n255 = ~x1 & x10 ;
  assign n256 = ~n254 & ~n255 ;
  assign n257 = x8 & ~x10 ;
  assign n258 = n257 ^ x2 ;
  assign n259 = x11 ^ x2 ;
  assign n260 = n259 ^ x2 ;
  assign n261 = ~n258 & n260 ;
  assign n262 = n261 ^ x2 ;
  assign n264 = n263 ^ n256 ;
  assign n265 = n262 & ~n264 ;
  assign n266 = n265 ^ n263 ;
  assign n267 = ~n256 & n266 ;
  assign n268 = n267 ^ n256 ;
  assign n269 = n253 & ~n268 ;
  assign n277 = n276 ^ n269 ;
  assign n278 = ~x4 & ~n277 ;
  assign n279 = n278 ^ n276 ;
  assign n280 = ~n246 & n279 ;
  assign n281 = ~n190 & n280 ;
  assign n282 = n281 ^ x19 ;
  assign n283 = n42 & n282 ;
  assign n284 = n283 ^ x19 ;
  assign n285 = x14 & n284 ;
  assign n286 = ~n39 & n285 ;
  assign y0 = ~n286 ;
endmodule
