module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 ;
  assign n13 = ~x8 & ~x11 ;
  assign n14 = ~x7 & ~n13 ;
  assign n15 = x0 & x1 ;
  assign n16 = ~x4 & x7 ;
  assign n17 = n15 & ~n16 ;
  assign n18 = x6 ^ x5 ;
  assign n19 = n17 & n18 ;
  assign n20 = n18 ^ x9 ;
  assign n21 = x3 & ~x8 ;
  assign n22 = x5 & n21 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = ~n20 & n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n19 & n25 ;
  assign n27 = ~n14 & n26 ;
  assign n28 = x2 & x7 ;
  assign n29 = ~x11 & n28 ;
  assign n30 = n29 ^ x9 ;
  assign n31 = n30 ^ n29 ;
  assign n44 = x8 & ~x10 ;
  assign n34 = ~x4 & ~x10 ;
  assign n35 = x3 & ~n34 ;
  assign n32 = x7 ^ x2 ;
  assign n36 = n35 ^ n32 ;
  assign n33 = n32 ^ x7 ;
  assign n37 = n36 ^ n33 ;
  assign n45 = n44 ^ n37 ;
  assign n49 = n45 ^ n36 ;
  assign n50 = n49 ^ n32 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = n38 ^ n32 ;
  assign n40 = n39 ^ n32 ;
  assign n41 = n36 ^ x11 ;
  assign n42 = n41 ^ n32 ;
  assign n43 = ~n40 & ~n42 ;
  assign n46 = n45 ^ n43 ;
  assign n47 = n46 ^ n32 ;
  assign n48 = ~n39 & ~n47 ;
  assign n51 = n50 ^ n48 ;
  assign n52 = n51 ^ n39 ;
  assign n53 = n32 ^ x5 ;
  assign n54 = n50 ^ n47 ;
  assign n55 = n54 ^ n39 ;
  assign n56 = ~n53 & n55 ;
  assign n57 = n56 ^ n32 ;
  assign n58 = ~n52 & n57 ;
  assign n59 = n58 ^ n56 ;
  assign n60 = n59 ^ n32 ;
  assign n61 = n60 ^ x7 ;
  assign n62 = n61 ^ n29 ;
  assign n63 = n31 & ~n62 ;
  assign n64 = n63 ^ n29 ;
  assign n65 = ~x5 & ~n29 ;
  assign n66 = n65 ^ n27 ;
  assign n67 = ~n64 & n66 ;
  assign n68 = n67 ^ n65 ;
  assign n69 = n27 & n68 ;
  assign n70 = n69 ^ n27 ;
  assign y0 = n70 ;
endmodule
