module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n15 = x1 & x5 ;
  assign n16 = x2 & n15 ;
  assign n17 = x3 & x4 ;
  assign n18 = x0 & n17 ;
  assign n19 = n16 & n18 ;
  assign n20 = x9 ^ x8 ;
  assign n21 = x9 & ~n20 ;
  assign n22 = x7 & n21 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = x6 & ~n23 ;
  assign n25 = ~x11 & ~x12 ;
  assign n26 = x10 & n25 ;
  assign n27 = n26 ^ x13 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = ~x8 & ~x9 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n30 ^ n26 ;
  assign n32 = n28 & ~n31 ;
  assign n33 = n32 ^ n26 ;
  assign n34 = x7 & n33 ;
  assign n35 = n34 ^ n26 ;
  assign n36 = ~n24 & ~n35 ;
  assign n37 = n19 & ~n36 ;
  assign y0 = n37 ;
endmodule
