module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n12 = x8 ^ x3 ;
  assign n13 = x7 ^ x2 ;
  assign n15 = x7 ^ x1 ;
  assign n14 = x7 ^ x6 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n16 ^ n13 ;
  assign n23 = n15 ^ x7 ;
  assign n18 = x7 ^ x5 ;
  assign n19 = n18 ^ x7 ;
  assign n20 = x7 ^ x0 ;
  assign n21 = n20 ^ x7 ;
  assign n22 = n19 & n21 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n17 & n24 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = n26 ^ n15 ;
  assign n28 = n27 ^ n23 ;
  assign n29 = n13 & ~n28 ;
  assign n30 = n29 ^ x2 ;
  assign n31 = n30 ^ x8 ;
  assign n32 = n12 & ~n31 ;
  assign n33 = n32 ^ x3 ;
  assign n11 = x9 ^ x4 ;
  assign n34 = n33 ^ n11 ;
  assign y0 = n34 ;
endmodule
