module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 ;
  output y0 ;
  wire n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 ;
  assign n35 = x3 & x5 ;
  assign n36 = x20 & x21 ;
  assign n37 = x25 & x26 ;
  assign n38 = x17 & ~n37 ;
  assign n39 = x13 & x24 ;
  assign n40 = n38 & n39 ;
  assign n41 = ~n36 & n40 ;
  assign n42 = ~x4 & x13 ;
  assign n43 = x4 & ~x13 ;
  assign n44 = x15 & ~x18 ;
  assign n45 = x19 & ~n44 ;
  assign n46 = n43 & ~n45 ;
  assign n47 = ~n42 & ~n46 ;
  assign n48 = ~n41 & n47 ;
  assign n49 = x3 & ~n48 ;
  assign n50 = ~x0 & ~n49 ;
  assign n51 = ~n35 & ~n50 ;
  assign n52 = ~x2 & n51 ;
  assign n53 = x29 & x31 ;
  assign n54 = x27 & x28 ;
  assign n55 = n53 & n54 ;
  assign n56 = ~x2 & ~x30 ;
  assign n57 = ~n55 & n56 ;
  assign n58 = ~x13 & ~n57 ;
  assign n59 = x15 ^ x14 ;
  assign n60 = x17 ^ x15 ;
  assign n61 = ~n59 & ~n60 ;
  assign n62 = x23 & n61 ;
  assign n63 = n62 ^ x2 ;
  assign n64 = n63 ^ n62 ;
  assign n65 = n64 ^ n58 ;
  assign n66 = x6 & x7 ;
  assign n67 = x9 ^ x8 ;
  assign n68 = n67 ^ x10 ;
  assign n69 = n68 ^ x11 ;
  assign n70 = x11 ^ x10 ;
  assign n71 = n70 ^ x11 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = x12 ^ x9 ;
  assign n74 = x11 & ~n73 ;
  assign n75 = n74 ^ x12 ;
  assign n76 = n72 & ~n75 ;
  assign n77 = n76 ^ n74 ;
  assign n78 = n77 ^ x12 ;
  assign n79 = n78 ^ x11 ;
  assign n80 = n69 & ~n79 ;
  assign n81 = n80 ^ n67 ;
  assign n82 = n81 ^ n66 ;
  assign n83 = n66 & n82 ;
  assign n84 = n83 ^ n62 ;
  assign n85 = n84 ^ n66 ;
  assign n86 = n65 & ~n85 ;
  assign n87 = n86 ^ n83 ;
  assign n88 = n87 ^ n66 ;
  assign n89 = ~n58 & n88 ;
  assign n90 = n89 ^ n58 ;
  assign n91 = ~x4 & n90 ;
  assign n92 = x4 & x14 ;
  assign n98 = n92 ^ x12 ;
  assign n93 = x16 & x17 ;
  assign n94 = ~x18 & n93 ;
  assign n95 = x19 & ~n94 ;
  assign n96 = ~n36 & ~n95 ;
  assign n97 = n96 ^ n92 ;
  assign n99 = n98 ^ n97 ;
  assign n100 = n98 ^ x15 ;
  assign n101 = n100 ^ n98 ;
  assign n102 = ~n99 & ~n101 ;
  assign n103 = n102 ^ n98 ;
  assign n104 = x2 & ~n103 ;
  assign n105 = n104 ^ n92 ;
  assign n106 = ~x13 & n105 ;
  assign n107 = ~n91 & ~n106 ;
  assign n108 = ~x5 & ~n107 ;
  assign n109 = ~x4 & ~x13 ;
  assign n110 = x33 & n109 ;
  assign n111 = n110 ^ x2 ;
  assign n112 = n111 ^ n110 ;
  assign n113 = n112 ^ x5 ;
  assign n114 = ~x32 & n42 ;
  assign n115 = x15 & n114 ;
  assign n116 = x21 & n43 ;
  assign n117 = ~x22 & n116 ;
  assign n118 = n117 ^ n115 ;
  assign n119 = ~n115 & n118 ;
  assign n120 = n119 ^ n110 ;
  assign n121 = n120 ^ n115 ;
  assign n122 = n113 & n121 ;
  assign n123 = n122 ^ n119 ;
  assign n124 = n123 ^ n115 ;
  assign n125 = x5 & ~n124 ;
  assign n126 = n125 ^ x5 ;
  assign n127 = ~n108 & ~n126 ;
  assign n128 = ~x3 & ~n127 ;
  assign n134 = x3 ^ x0 ;
  assign n133 = x2 ^ x0 ;
  assign n135 = n134 ^ n133 ;
  assign n130 = x13 ^ x0 ;
  assign n136 = n135 ^ n130 ;
  assign n137 = n136 ^ n133 ;
  assign n129 = x4 ^ x0 ;
  assign n131 = n130 ^ n129 ;
  assign n138 = n137 ^ n131 ;
  assign n139 = n138 ^ x0 ;
  assign n132 = n131 ^ n130 ;
  assign n140 = n139 ^ n132 ;
  assign n141 = n132 ^ n130 ;
  assign n142 = n140 & n141 ;
  assign n143 = n142 ^ n139 ;
  assign n144 = n139 ^ n136 ;
  assign n145 = n144 ^ n130 ;
  assign n146 = n145 ^ n132 ;
  assign n149 = x5 ^ x0 ;
  assign n150 = n149 ^ x0 ;
  assign n151 = n150 ^ x0 ;
  assign n152 = n145 & n151 ;
  assign n147 = n130 ^ x0 ;
  assign n148 = ~n130 & ~n147 ;
  assign n153 = n152 ^ n148 ;
  assign n154 = n153 ^ n130 ;
  assign n155 = ~n146 & ~n154 ;
  assign n156 = n155 ^ n152 ;
  assign n157 = n156 ^ x0 ;
  assign n158 = ~n143 & n157 ;
  assign n159 = n158 ^ n152 ;
  assign n160 = n159 ^ n148 ;
  assign n161 = n160 ^ n155 ;
  assign n162 = n161 ^ x0 ;
  assign n163 = n162 ^ n130 ;
  assign n164 = n163 ^ x0 ;
  assign n165 = ~n128 & n164 ;
  assign n166 = ~n52 & n165 ;
  assign n167 = x1 & ~n166 ;
  assign y0 = n167 ;
endmodule
