// Benchmark "./pla/newcwp.pla_res_2NonExact" written by ABC on Fri Nov 20 10:27:08 2020

module \./pla/newcwp.pla_res_2NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = ~x0;
endmodule


