module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 ;
  assign n9 = x1 & x6 ;
  assign n10 = x0 & n9 ;
  assign n11 = ~x3 & x4 ;
  assign n12 = n11 ^ x2 ;
  assign n13 = n11 ^ x5 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = x7 ^ x5 ;
  assign n16 = ~n14 & ~n15 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = ~n12 & n17 ;
  assign n19 = n10 & n18 ;
  assign y0 = n19 ;
endmodule
