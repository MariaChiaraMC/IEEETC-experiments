module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 ;
  assign n44 = ~x0 & ~x2 ;
  assign n40 = x0 & ~x3 ;
  assign n41 = x7 & n40 ;
  assign n45 = n44 ^ n41 ;
  assign n46 = n45 ^ n41 ;
  assign n17 = x5 ^ x3 ;
  assign n18 = n17 ^ x3 ;
  assign n19 = n18 ^ x7 ;
  assign n20 = n19 ^ x7 ;
  assign n22 = x4 ^ x3 ;
  assign n21 = x6 ^ x3 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n23 ^ x7 ;
  assign n25 = n24 ^ n20 ;
  assign n29 = n20 ^ n19 ;
  assign n30 = ~x3 & n29 ;
  assign n26 = n22 ^ x3 ;
  assign n27 = n26 ^ x3 ;
  assign n28 = ~n19 & ~n27 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n31 ^ x3 ;
  assign n33 = n32 ^ n26 ;
  assign n34 = n25 & ~n33 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = ~n20 & n35 ;
  assign n37 = n36 ^ n28 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = n38 ^ x3 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = n42 ^ n41 ;
  assign n47 = n46 ^ n43 ;
  assign n48 = x9 & ~x11 ;
  assign n49 = ~x8 & n48 ;
  assign n50 = ~x12 & n49 ;
  assign n51 = n50 ^ x10 ;
  assign n52 = ~x14 & ~x15 ;
  assign n53 = n52 ^ x13 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = x15 ^ x14 ;
  assign n56 = n55 ^ n52 ;
  assign n57 = ~n54 & n56 ;
  assign n58 = n57 ^ n52 ;
  assign n59 = n58 ^ n50 ;
  assign n60 = ~n51 & n59 ;
  assign n61 = n60 ^ n57 ;
  assign n62 = n61 ^ n52 ;
  assign n63 = n62 ^ x10 ;
  assign n64 = n50 & ~n63 ;
  assign n65 = n64 ^ n50 ;
  assign n66 = ~x3 & ~n65 ;
  assign n67 = n66 ^ n41 ;
  assign n68 = n67 ^ n41 ;
  assign n69 = n68 ^ n46 ;
  assign n70 = n46 & ~n69 ;
  assign n71 = n70 ^ n46 ;
  assign n72 = ~n47 & n71 ;
  assign n73 = n72 ^ n70 ;
  assign n74 = n73 ^ n41 ;
  assign n75 = n74 ^ n46 ;
  assign n76 = x1 & n75 ;
  assign n77 = n76 ^ n41 ;
  assign y0 = n77 ;
endmodule
