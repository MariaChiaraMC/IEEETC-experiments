module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n16 = x13 & x14 ;
  assign n17 = x4 & x9 ;
  assign n18 = n16 & n17 ;
  assign n19 = x2 & x3 ;
  assign n20 = x11 & n19 ;
  assign n21 = n18 & n20 ;
  assign n22 = x0 & ~x1 ;
  assign n23 = x10 & x12 ;
  assign n24 = n22 & n23 ;
  assign n25 = x6 ^ x5 ;
  assign n26 = n25 ^ x5 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = x8 ^ x5 ;
  assign n29 = n28 ^ x7 ;
  assign n30 = x7 & ~n29 ;
  assign n31 = n30 ^ x5 ;
  assign n32 = n31 ^ x7 ;
  assign n33 = n27 & ~n32 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ x7 ;
  assign n36 = n24 & n35 ;
  assign n37 = n21 & n36 ;
  assign y0 = n37 ;
endmodule
