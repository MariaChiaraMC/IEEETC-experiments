// Benchmark "./pla/sqr6.pla_res_8NonExact" written by ABC on Fri Nov 20 10:29:19 2020

module \./pla/sqr6.pla_res_8NonExact  ( 
    x0, x1,
    z0  );
  input  x0, x1;
  output z0;
  assign z0 = x0 & x1;
endmodule


