module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 ;
  output y0 ;
  wire n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 ;
  assign n26 = ~x12 & ~x17 ;
  assign n27 = ~x18 & n26 ;
  assign n28 = ~x16 & ~x19 ;
  assign n29 = ~x15 & n28 ;
  assign n30 = n27 & n29 ;
  assign n31 = x10 & ~x11 ;
  assign n32 = n30 & n31 ;
  assign n33 = x12 & x17 ;
  assign n34 = x18 & n33 ;
  assign n35 = x16 & x19 ;
  assign n36 = x15 & n35 ;
  assign n37 = n34 & n36 ;
  assign n38 = x11 & n37 ;
  assign n39 = x7 & n38 ;
  assign n40 = ~n32 & ~n39 ;
  assign n41 = x1 ^ x0 ;
  assign n42 = x1 & x2 ;
  assign n43 = ~n41 & n42 ;
  assign n44 = n43 ^ n41 ;
  assign n45 = ~n40 & ~n44 ;
  assign n46 = ~x2 & ~x9 ;
  assign n47 = n30 & ~n46 ;
  assign n48 = n47 ^ n37 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = x6 ^ x3 ;
  assign n51 = ~x2 & n50 ;
  assign n52 = n51 ^ x3 ;
  assign n53 = n52 ^ n47 ;
  assign n54 = n53 ^ n47 ;
  assign n55 = n49 & n54 ;
  assign n56 = n55 ^ n47 ;
  assign n57 = x11 & n56 ;
  assign n58 = n57 ^ n47 ;
  assign n59 = ~x0 & ~x1 ;
  assign n60 = ~x8 & ~x11 ;
  assign n61 = ~n59 & ~n60 ;
  assign n62 = n61 ^ x2 ;
  assign n63 = n62 ^ n61 ;
  assign n64 = ~x4 & ~x5 ;
  assign n65 = n64 ^ n61 ;
  assign n66 = ~n63 & n65 ;
  assign n67 = n66 ^ n61 ;
  assign n68 = n58 & n67 ;
  assign n69 = ~n45 & ~n68 ;
  assign y0 = ~n69 ;
endmodule
