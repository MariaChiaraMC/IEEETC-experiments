module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 ;
  output y0 ;
  wire n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 ;
  assign n26 = x10 ^ x8 ;
  assign n27 = n26 ^ x8 ;
  assign n28 = x8 ^ x1 ;
  assign n29 = n28 ^ x8 ;
  assign n30 = n27 & n29 ;
  assign n31 = n30 ^ x8 ;
  assign n32 = ~x2 & n31 ;
  assign n33 = n32 ^ x8 ;
  assign n34 = x0 & n33 ;
  assign n35 = ~x2 & ~x4 ;
  assign n36 = ~x5 & x9 ;
  assign n37 = n35 & n36 ;
  assign n39 = x2 & x8 ;
  assign n38 = ~x0 & x10 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = ~x1 & n40 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = ~n37 & ~n42 ;
  assign n44 = ~n34 & n43 ;
  assign n45 = ~x16 & ~x19 ;
  assign n46 = ~x11 & ~x17 ;
  assign n47 = ~x18 & n46 ;
  assign n48 = ~x12 & n47 ;
  assign n49 = n45 & n48 ;
  assign n50 = ~n44 & n49 ;
  assign y0 = n50 ;
endmodule
