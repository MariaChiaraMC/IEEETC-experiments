module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 ;
  assign n16 = ~x0 & ~x11 ;
  assign n17 = ~x13 & ~x14 ;
  assign n64 = ~x3 & n17 ;
  assign n18 = ~x10 & n17 ;
  assign n19 = ~x1 & ~x4 ;
  assign n20 = n18 & n19 ;
  assign n21 = x5 & n20 ;
  assign n22 = x8 ^ x7 ;
  assign n23 = x8 ^ x3 ;
  assign n24 = n23 ^ x3 ;
  assign n25 = x3 & x9 ;
  assign n26 = n25 ^ x3 ;
  assign n27 = ~n24 & ~n26 ;
  assign n28 = n27 ^ x3 ;
  assign n29 = ~n22 & ~n28 ;
  assign n30 = ~x2 & n29 ;
  assign n31 = n21 & n30 ;
  assign n32 = x1 & n25 ;
  assign n33 = x4 & n32 ;
  assign n34 = x2 & ~x8 ;
  assign n35 = x5 & x7 ;
  assign n36 = n34 & ~n35 ;
  assign n37 = n33 & n36 ;
  assign n38 = x5 & ~x13 ;
  assign n39 = ~n17 & ~n38 ;
  assign n40 = n37 & n39 ;
  assign n41 = ~n31 & ~n40 ;
  assign n42 = ~x6 & ~n41 ;
  assign n43 = x10 ^ x7 ;
  assign n44 = x13 ^ x5 ;
  assign n45 = n44 ^ n43 ;
  assign n46 = x14 ^ x10 ;
  assign n47 = ~x5 & n46 ;
  assign n48 = n47 ^ x10 ;
  assign n49 = n45 & ~n48 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = n50 ^ x10 ;
  assign n52 = n51 ^ x5 ;
  assign n53 = ~n43 & n52 ;
  assign n54 = n33 & n53 ;
  assign n55 = ~x3 & ~x7 ;
  assign n56 = x6 & n55 ;
  assign n57 = n20 & n56 ;
  assign n58 = ~x5 & n57 ;
  assign n59 = ~n54 & ~n58 ;
  assign n60 = n34 & ~n59 ;
  assign n61 = ~n42 & ~n60 ;
  assign n65 = n64 ^ n61 ;
  assign n66 = n65 ^ n61 ;
  assign n62 = n61 ^ x10 ;
  assign n63 = n62 ^ n61 ;
  assign n67 = n66 ^ n63 ;
  assign n68 = x4 & n34 ;
  assign n69 = ~x1 & x5 ;
  assign n70 = ~x6 & n69 ;
  assign n71 = n68 & n70 ;
  assign n72 = x9 & n71 ;
  assign n73 = n72 ^ n61 ;
  assign n74 = n73 ^ n61 ;
  assign n75 = n74 ^ n66 ;
  assign n76 = n66 & n75 ;
  assign n77 = n76 ^ n66 ;
  assign n78 = n67 & n77 ;
  assign n79 = n78 ^ n76 ;
  assign n80 = n79 ^ n61 ;
  assign n81 = n80 ^ n66 ;
  assign n82 = x12 & ~n81 ;
  assign n83 = n82 ^ n61 ;
  assign n84 = n16 & ~n83 ;
  assign y0 = n84 ;
endmodule
