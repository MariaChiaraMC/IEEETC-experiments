module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 ;
  assign n8 = x4 ^ x1 ;
  assign n11 = x3 ^ x0 ;
  assign n12 = x6 ^ x3 ;
  assign n13 = n11 & ~n12 ;
  assign n14 = n13 ^ x0 ;
  assign n9 = x4 ^ x2 ;
  assign n10 = n9 ^ x5 ;
  assign n15 = n14 ^ n10 ;
  assign n16 = n15 ^ n9 ;
  assign n17 = x5 ^ x4 ;
  assign n18 = n17 ^ n9 ;
  assign n19 = ~n16 & n18 ;
  assign n20 = n19 ^ n9 ;
  assign n21 = n8 & ~n20 ;
  assign n22 = n21 ^ x1 ;
  assign y0 = n22 ;
endmodule
