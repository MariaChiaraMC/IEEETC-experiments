module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 ;
  assign n16 = x7 & ~x11 ;
  assign n17 = x13 & n16 ;
  assign n18 = ~x5 & x9 ;
  assign n19 = x4 & n18 ;
  assign n20 = n17 & n19 ;
  assign n21 = ~x13 & ~x14 ;
  assign n22 = ~x11 & ~x13 ;
  assign n23 = ~x10 & ~n22 ;
  assign n24 = ~n21 & n23 ;
  assign n25 = ~x7 & ~x8 ;
  assign n26 = ~x13 & x14 ;
  assign n27 = x11 & n26 ;
  assign n28 = ~x4 & ~x5 ;
  assign n29 = x6 & n28 ;
  assign n30 = n27 & n29 ;
  assign n31 = n25 & n30 ;
  assign n32 = ~n24 & ~n31 ;
  assign n35 = n32 ^ x5 ;
  assign n36 = n35 ^ n32 ;
  assign n33 = n32 ^ n27 ;
  assign n34 = n33 ^ n32 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = ~x3 & x4 ;
  assign n39 = n38 ^ n32 ;
  assign n40 = n39 ^ n32 ;
  assign n41 = n40 ^ n36 ;
  assign n42 = n36 & n41 ;
  assign n43 = n42 ^ n36 ;
  assign n44 = n37 & n43 ;
  assign n45 = n44 ^ n42 ;
  assign n46 = n45 ^ n32 ;
  assign n47 = n46 ^ n36 ;
  assign n48 = ~x9 & ~n47 ;
  assign n49 = n48 ^ n32 ;
  assign n50 = ~n20 & n49 ;
  assign n51 = ~x0 & ~n50 ;
  assign n52 = ~x10 & x11 ;
  assign n53 = x14 & n52 ;
  assign n54 = x13 & n53 ;
  assign n55 = ~x11 & ~x14 ;
  assign n56 = ~x3 & n55 ;
  assign n57 = x13 & n56 ;
  assign n58 = ~x6 & x7 ;
  assign n59 = n28 & n58 ;
  assign n60 = x11 & n21 ;
  assign n61 = x8 & n60 ;
  assign n62 = n59 & n61 ;
  assign n63 = x5 & x14 ;
  assign n64 = x3 & ~n63 ;
  assign n65 = n52 & ~n64 ;
  assign n66 = ~x3 & ~x13 ;
  assign n67 = ~x4 & n66 ;
  assign n68 = ~n60 & ~n67 ;
  assign n69 = ~x10 & ~n68 ;
  assign n70 = ~n65 & ~n69 ;
  assign n71 = ~n62 & n70 ;
  assign n72 = ~n57 & n71 ;
  assign n73 = n72 ^ x1 ;
  assign n74 = n73 ^ x9 ;
  assign n84 = n74 ^ n73 ;
  assign n75 = ~x9 & x13 ;
  assign n76 = x10 & n75 ;
  assign n77 = n55 & n76 ;
  assign n78 = n77 ^ n74 ;
  assign n79 = n78 ^ n73 ;
  assign n80 = n74 ^ n72 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n81 ^ n79 ;
  assign n83 = n79 & n82 ;
  assign n85 = n84 ^ n83 ;
  assign n86 = n85 ^ n79 ;
  assign n87 = n73 ^ n53 ;
  assign n88 = n83 ^ n79 ;
  assign n89 = ~n87 & n88 ;
  assign n90 = n89 ^ n73 ;
  assign n91 = ~n86 & n90 ;
  assign n92 = n91 ^ n73 ;
  assign n93 = n92 ^ x1 ;
  assign n94 = n93 ^ n73 ;
  assign n95 = ~n54 & n94 ;
  assign n96 = ~n51 & n95 ;
  assign n97 = ~x12 & ~n96 ;
  assign n98 = n21 ^ x13 ;
  assign n99 = n98 ^ x13 ;
  assign n100 = x13 ^ x3 ;
  assign n101 = n100 ^ x13 ;
  assign n102 = ~n99 & n101 ;
  assign n103 = n102 ^ x13 ;
  assign n104 = ~x9 & ~n103 ;
  assign n105 = n104 ^ x13 ;
  assign n106 = x12 & ~n105 ;
  assign n107 = ~x11 & n106 ;
  assign n108 = x13 & ~x14 ;
  assign n109 = ~x7 & n108 ;
  assign n110 = n109 ^ x14 ;
  assign n111 = ~n25 & n66 ;
  assign n112 = ~x7 & x8 ;
  assign n113 = ~x5 & n112 ;
  assign n114 = n113 ^ x8 ;
  assign n115 = n111 & ~n114 ;
  assign n116 = n115 ^ x6 ;
  assign n117 = n116 ^ n115 ;
  assign n118 = n117 ^ n110 ;
  assign n119 = n112 ^ x13 ;
  assign n120 = n112 & n119 ;
  assign n121 = n120 ^ n115 ;
  assign n122 = n121 ^ n112 ;
  assign n123 = n118 & n122 ;
  assign n124 = n123 ^ n120 ;
  assign n125 = n124 ^ n112 ;
  assign n126 = n110 & n125 ;
  assign n127 = n126 ^ n110 ;
  assign n128 = x12 & ~n127 ;
  assign n129 = n22 & ~n25 ;
  assign n130 = n29 & n129 ;
  assign n131 = x8 ^ x0 ;
  assign n132 = x14 ^ x3 ;
  assign n133 = x8 ^ x3 ;
  assign n134 = n133 ^ x3 ;
  assign n135 = ~n132 & ~n134 ;
  assign n136 = n135 ^ x3 ;
  assign n137 = n131 & n136 ;
  assign n138 = n137 ^ x0 ;
  assign n139 = n130 & ~n138 ;
  assign n140 = ~x0 & ~x13 ;
  assign n141 = x11 & ~n26 ;
  assign n142 = ~n140 & n141 ;
  assign n143 = ~n139 & ~n142 ;
  assign n144 = ~n128 & n143 ;
  assign n145 = n144 ^ n56 ;
  assign n146 = x8 & n29 ;
  assign n147 = ~x13 & n146 ;
  assign n148 = n147 ^ n144 ;
  assign n149 = n144 ^ x9 ;
  assign n150 = n144 & n149 ;
  assign n151 = n150 ^ n144 ;
  assign n152 = n148 & n151 ;
  assign n153 = n152 ^ n150 ;
  assign n154 = n153 ^ n144 ;
  assign n155 = n154 ^ x9 ;
  assign n156 = ~n145 & n155 ;
  assign n157 = n156 ^ n56 ;
  assign n158 = ~n107 & ~n157 ;
  assign n159 = ~x10 & ~n158 ;
  assign n160 = ~x0 & n38 ;
  assign n161 = ~x5 & x7 ;
  assign n162 = x1 & n108 ;
  assign n163 = n161 & n162 ;
  assign n164 = ~x2 & ~x13 ;
  assign n165 = x5 & ~x6 ;
  assign n166 = ~x1 & n165 ;
  assign n167 = n166 ^ x5 ;
  assign n168 = n164 & n167 ;
  assign n169 = ~n163 & ~n168 ;
  assign n170 = n160 & ~n169 ;
  assign n171 = x11 & n170 ;
  assign n172 = ~x8 & ~x11 ;
  assign n173 = n26 & n172 ;
  assign n174 = n59 & n173 ;
  assign n175 = ~x4 & n60 ;
  assign n176 = ~n174 & ~n175 ;
  assign n177 = ~n171 & n176 ;
  assign n178 = ~x9 & ~n177 ;
  assign n179 = x3 & ~x9 ;
  assign n180 = x13 & x14 ;
  assign n181 = ~x6 & ~x11 ;
  assign n182 = n28 & n181 ;
  assign n183 = n180 & n182 ;
  assign n184 = n112 & n183 ;
  assign n185 = ~n179 & n184 ;
  assign n186 = ~n178 & ~n185 ;
  assign n187 = n186 ^ x12 ;
  assign n188 = n187 ^ n186 ;
  assign n189 = n188 ^ x10 ;
  assign n190 = n16 ^ x9 ;
  assign n191 = n190 ^ n16 ;
  assign n192 = n191 ^ x14 ;
  assign n193 = n167 ^ n16 ;
  assign n194 = n193 ^ x13 ;
  assign n195 = ~x13 & ~n194 ;
  assign n196 = n195 ^ n16 ;
  assign n197 = n196 ^ x13 ;
  assign n198 = ~n192 & ~n197 ;
  assign n199 = n198 ^ n195 ;
  assign n200 = n199 ^ x13 ;
  assign n201 = x14 & ~n200 ;
  assign n202 = n201 ^ n16 ;
  assign n203 = n160 & n202 ;
  assign n204 = x5 & x6 ;
  assign n205 = x0 & ~n204 ;
  assign n206 = x4 & ~n205 ;
  assign n207 = x14 ^ x9 ;
  assign n218 = n207 ^ x14 ;
  assign n208 = x5 & ~x7 ;
  assign n209 = n208 ^ n207 ;
  assign n210 = n209 ^ x14 ;
  assign n211 = n210 ^ x14 ;
  assign n212 = n211 ^ n207 ;
  assign n213 = n212 ^ x14 ;
  assign n214 = n165 ^ x13 ;
  assign n215 = ~n213 & n214 ;
  assign n216 = n215 ^ x13 ;
  assign n217 = n216 ^ x14 ;
  assign n219 = n218 ^ n217 ;
  assign n220 = n219 ^ n212 ;
  assign n221 = n218 ^ x14 ;
  assign n222 = ~n218 & n221 ;
  assign n223 = n222 ^ x14 ;
  assign n224 = n223 ^ n212 ;
  assign n225 = n165 ^ x14 ;
  assign n226 = n225 ^ x3 ;
  assign n227 = ~n165 & n226 ;
  assign n228 = n227 ^ x14 ;
  assign n229 = n228 ^ n218 ;
  assign n230 = ~n224 & n229 ;
  assign n231 = n230 ^ n212 ;
  assign n232 = ~n220 & n231 ;
  assign n233 = n232 ^ n222 ;
  assign n234 = n233 ^ n215 ;
  assign n235 = n234 ^ x13 ;
  assign n236 = n235 ^ x14 ;
  assign n237 = n236 ^ n218 ;
  assign n238 = n237 ^ n212 ;
  assign n239 = n238 ^ x9 ;
  assign n240 = n239 ^ x14 ;
  assign n241 = n206 & ~n240 ;
  assign n242 = x4 & n161 ;
  assign n243 = n108 & ~n242 ;
  assign n244 = ~x9 & n243 ;
  assign n245 = ~n241 & ~n244 ;
  assign n246 = ~x11 & ~n245 ;
  assign n247 = x6 & n55 ;
  assign n248 = x8 ^ x6 ;
  assign n249 = n248 ^ x8 ;
  assign n250 = ~n133 & n249 ;
  assign n251 = n250 ^ x8 ;
  assign n252 = x11 & n251 ;
  assign n253 = ~x4 & n252 ;
  assign n254 = ~n247 & ~n253 ;
  assign n255 = ~x7 & ~x13 ;
  assign n256 = ~n254 & n255 ;
  assign n257 = ~x14 & n181 ;
  assign n258 = ~n25 & n257 ;
  assign n259 = ~n256 & ~n258 ;
  assign n260 = n18 & ~n259 ;
  assign n261 = ~x0 & n260 ;
  assign n262 = ~n246 & ~n261 ;
  assign n263 = n262 ^ n203 ;
  assign n264 = ~n203 & ~n263 ;
  assign n265 = n264 ^ n186 ;
  assign n266 = n265 ^ n203 ;
  assign n267 = ~n189 & ~n266 ;
  assign n268 = n267 ^ n264 ;
  assign n269 = n268 ^ n203 ;
  assign n270 = x10 & ~n269 ;
  assign n271 = n270 ^ x10 ;
  assign n272 = ~n159 & ~n271 ;
  assign n273 = ~n97 & n272 ;
  assign y0 = ~n273 ;
endmodule
