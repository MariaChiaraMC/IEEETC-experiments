// Benchmark "./f51m.pla" written by ABC on Thu Apr 23 10:59:51 2020

module \./f51m.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z6  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z6;
  assign z6 = 1'b1;
endmodule


