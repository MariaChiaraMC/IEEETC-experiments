module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n20 = ~x7 & ~x9 ;
  assign n21 = x16 & x18 ;
  assign n22 = ~x3 & n21 ;
  assign n23 = n20 & n22 ;
  assign n24 = x0 & x14 ;
  assign n25 = n23 & n24 ;
  assign n26 = ~x4 & x10 ;
  assign n27 = x11 & n26 ;
  assign n28 = ~x1 & ~x5 ;
  assign n29 = n27 & n28 ;
  assign n30 = x15 & x17 ;
  assign n31 = x12 & x13 ;
  assign n32 = n30 & n31 ;
  assign n33 = x2 & x8 ;
  assign n34 = ~x6 & n33 ;
  assign n35 = n32 & n34 ;
  assign n36 = n29 & n35 ;
  assign n37 = n25 & n36 ;
  assign y0 = n37 ;
endmodule
