module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 ;
  assign n10 = ~x3 & ~x4 ;
  assign n11 = ~x2 & x6 ;
  assign n12 = n10 & n11 ;
  assign n13 = x1 & n12 ;
  assign n27 = x4 & x8 ;
  assign n111 = x3 & x7 ;
  assign n112 = ~n27 & ~n111 ;
  assign n67 = x2 & ~x7 ;
  assign n107 = x8 & ~n10 ;
  assign n108 = n67 & ~n107 ;
  assign n113 = n112 ^ n108 ;
  assign n114 = n113 ^ n108 ;
  assign n60 = ~x3 & ~x7 ;
  assign n109 = n108 ^ n60 ;
  assign n110 = n109 ^ n108 ;
  assign n115 = n114 ^ n110 ;
  assign n116 = n108 ^ x2 ;
  assign n117 = n116 ^ n108 ;
  assign n118 = n117 ^ n114 ;
  assign n119 = ~n114 & ~n118 ;
  assign n120 = n119 ^ n114 ;
  assign n121 = n115 & ~n120 ;
  assign n122 = n121 ^ n119 ;
  assign n123 = n122 ^ n108 ;
  assign n124 = n123 ^ n114 ;
  assign n125 = ~x1 & ~n124 ;
  assign n126 = n125 ^ n108 ;
  assign n127 = x6 & n126 ;
  assign n128 = x8 ^ x2 ;
  assign n135 = n128 ^ x8 ;
  assign n129 = n128 ^ x3 ;
  assign n130 = n129 ^ x8 ;
  assign n131 = x8 ^ x6 ;
  assign n132 = n131 ^ x3 ;
  assign n133 = n132 ^ n130 ;
  assign n134 = n130 & ~n133 ;
  assign n136 = n135 ^ n134 ;
  assign n137 = n136 ^ n130 ;
  assign n138 = x8 ^ x4 ;
  assign n139 = n138 ^ x8 ;
  assign n140 = n134 ^ n130 ;
  assign n141 = ~n139 & n140 ;
  assign n142 = n141 ^ x8 ;
  assign n143 = n137 & n142 ;
  assign n144 = n143 ^ x8 ;
  assign n145 = n144 ^ x8 ;
  assign n146 = x7 & n145 ;
  assign n147 = n11 & ~n111 ;
  assign n148 = ~n10 & n147 ;
  assign n149 = ~n146 & ~n148 ;
  assign n150 = x1 & ~n149 ;
  assign n151 = ~n127 & ~n150 ;
  assign n15 = x6 & ~x8 ;
  assign n16 = ~x7 & n15 ;
  assign n48 = ~x4 & n16 ;
  assign n20 = ~x4 & ~x8 ;
  assign n49 = ~x7 & ~n27 ;
  assign n50 = ~n20 & n49 ;
  assign n51 = x6 & ~n50 ;
  assign n52 = x7 ^ x2 ;
  assign n53 = n52 ^ n27 ;
  assign n54 = ~n51 & n53 ;
  assign n55 = ~n48 & ~n54 ;
  assign n56 = x3 & ~n55 ;
  assign n14 = x2 & ~x3 ;
  assign n17 = x4 & x6 ;
  assign n18 = ~n16 & n17 ;
  assign n19 = n14 & ~n18 ;
  assign n23 = x7 & ~x8 ;
  assign n24 = x2 & ~n23 ;
  assign n21 = x7 & ~n20 ;
  assign n22 = x2 & ~n21 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n25 ^ x6 ;
  assign n35 = n26 ^ n25 ;
  assign n28 = x7 & n27 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = n26 ^ n22 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n30 & n33 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = n25 ^ x4 ;
  assign n39 = n34 ^ n30 ;
  assign n40 = n38 & n39 ;
  assign n41 = n40 ^ n25 ;
  assign n42 = ~n37 & ~n41 ;
  assign n43 = n42 ^ n25 ;
  assign n44 = n43 ^ n24 ;
  assign n45 = n44 ^ n25 ;
  assign n46 = x3 & ~n45 ;
  assign n47 = ~n19 & ~n46 ;
  assign n57 = n56 ^ n47 ;
  assign n58 = n57 ^ n47 ;
  assign n59 = ~x6 & x8 ;
  assign n61 = ~n59 & ~n60 ;
  assign n62 = ~x2 & ~n61 ;
  assign n63 = n62 ^ x6 ;
  assign n64 = n62 ^ x7 ;
  assign n65 = n64 ^ x7 ;
  assign n66 = n65 ^ n63 ;
  assign n68 = n67 ^ x7 ;
  assign n69 = x8 & n68 ;
  assign n70 = n69 ^ x7 ;
  assign n71 = n70 ^ x3 ;
  assign n72 = ~x3 & ~n71 ;
  assign n73 = n72 ^ x7 ;
  assign n74 = n73 ^ x3 ;
  assign n75 = ~n66 & n74 ;
  assign n76 = n75 ^ n72 ;
  assign n77 = n76 ^ x3 ;
  assign n78 = n63 & ~n77 ;
  assign n79 = n78 ^ n62 ;
  assign n80 = n79 ^ n14 ;
  assign n81 = n80 ^ x4 ;
  assign n89 = n81 ^ n80 ;
  assign n82 = ~x6 & ~x7 ;
  assign n83 = n82 ^ n81 ;
  assign n84 = n83 ^ n80 ;
  assign n85 = n81 ^ n79 ;
  assign n86 = n85 ^ n82 ;
  assign n87 = n86 ^ n84 ;
  assign n88 = ~n84 & ~n87 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = n90 ^ n84 ;
  assign n92 = x7 & ~n59 ;
  assign n93 = n92 ^ n80 ;
  assign n94 = n88 ^ n84 ;
  assign n95 = ~n93 & ~n94 ;
  assign n96 = n95 ^ n80 ;
  assign n97 = ~n91 & n96 ;
  assign n98 = n97 ^ n80 ;
  assign n99 = n98 ^ n14 ;
  assign n100 = n99 ^ n80 ;
  assign n101 = n100 ^ n47 ;
  assign n102 = n101 ^ n47 ;
  assign n103 = ~n58 & ~n102 ;
  assign n104 = n103 ^ n47 ;
  assign n105 = x1 & n104 ;
  assign n106 = n105 ^ n47 ;
  assign n152 = n151 ^ n106 ;
  assign n153 = n152 ^ n151 ;
  assign n154 = n17 & n111 ;
  assign n155 = x8 & n154 ;
  assign n156 = n155 ^ n151 ;
  assign n157 = n156 ^ n151 ;
  assign n158 = n153 & ~n157 ;
  assign n159 = n158 ^ n151 ;
  assign n160 = x5 & n159 ;
  assign n161 = n160 ^ n151 ;
  assign n162 = ~n13 & n161 ;
  assign n163 = x0 & ~n162 ;
  assign y0 = n163 ;
endmodule
