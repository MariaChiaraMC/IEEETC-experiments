module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 ;
  assign n9 = x0 & ~x3 ;
  assign n10 = x5 ^ x4 ;
  assign n11 = n10 ^ x1 ;
  assign n13 = x6 ^ x5 ;
  assign n14 = n13 ^ x6 ;
  assign n12 = x2 ^ x1 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n16 ^ n10 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = n18 ^ x1 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = ~n11 & ~n20 ;
  assign n22 = n21 ^ n11 ;
  assign n23 = n22 ^ n10 ;
  assign n24 = n13 ^ x1 ;
  assign n25 = n24 ^ n10 ;
  assign n26 = n25 ^ n17 ;
  assign n27 = n25 ^ n10 ;
  assign n28 = ~n26 & ~n27 ;
  assign n29 = n28 ^ n10 ;
  assign n30 = n14 ^ x7 ;
  assign n31 = n30 ^ n14 ;
  assign n32 = n31 ^ n19 ;
  assign n33 = n32 ^ n10 ;
  assign n34 = ~n25 & ~n33 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = n35 ^ n10 ;
  assign n37 = n36 ^ n25 ;
  assign n38 = n29 & ~n37 ;
  assign n39 = n38 ^ n11 ;
  assign n40 = n39 ^ n19 ;
  assign n41 = ~n23 & n40 ;
  assign n42 = n41 ^ n10 ;
  assign n43 = n42 ^ n10 ;
  assign n44 = n9 & n43 ;
  assign y0 = n44 ;
endmodule
