module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 ;
  assign n13 = x2 & x3 ;
  assign n14 = n13 ^ x6 ;
  assign n15 = n13 ^ x5 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = n15 ^ x11 ;
  assign n18 = n16 & ~n17 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = ~x10 & ~n15 ;
  assign n21 = n20 ^ n14 ;
  assign n22 = ~n19 & ~n21 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = ~n14 & n23 ;
  assign n25 = n24 ^ n14 ;
  assign n28 = n25 ^ x2 ;
  assign n29 = n28 ^ n25 ;
  assign n26 = n25 ^ x6 ;
  assign n27 = n26 ^ n25 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = ~x3 & x5 ;
  assign n32 = n31 ^ n25 ;
  assign n33 = n32 ^ n25 ;
  assign n34 = n33 ^ n29 ;
  assign n35 = n29 & n34 ;
  assign n36 = n35 ^ n29 ;
  assign n37 = n30 & n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = n38 ^ n25 ;
  assign n40 = n39 ^ n29 ;
  assign n41 = ~x4 & ~n40 ;
  assign n42 = n41 ^ n25 ;
  assign y0 = ~n42 ;
endmodule
