module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 ;
  assign n11 = ~x4 & x8 ;
  assign n12 = ~x5 & x9 ;
  assign n13 = ~n11 & ~n12 ;
  assign n15 = ~x0 & ~x6 ;
  assign n16 = x2 & ~n15 ;
  assign n17 = ~x1 & n16 ;
  assign n14 = x3 & ~x7 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = n18 ^ n14 ;
  assign n20 = ~x2 & x6 ;
  assign n21 = x7 ^ x3 ;
  assign n22 = ~n20 & ~n21 ;
  assign n23 = n22 ^ n14 ;
  assign n24 = ~n19 & n23 ;
  assign n25 = n24 ^ n14 ;
  assign n26 = n13 & n25 ;
  assign y0 = n26 ;
endmodule
