module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 ;
  assign n10 = ~x4 & ~x8 ;
  assign n11 = ~x0 & n10 ;
  assign n12 = x2 & ~x3 ;
  assign n13 = ~x1 & ~x6 ;
  assign n14 = n12 & n13 ;
  assign n15 = n11 & n14 ;
  assign n79 = x2 & ~x6 ;
  assign n20 = x1 & x3 ;
  assign n80 = n11 & n20 ;
  assign n81 = ~n79 & n80 ;
  assign n51 = x1 & x2 ;
  assign n82 = x4 & ~x8 ;
  assign n83 = ~x4 & x8 ;
  assign n84 = n83 ^ x6 ;
  assign n85 = n84 ^ x6 ;
  assign n86 = x3 & ~x6 ;
  assign n87 = n86 ^ x6 ;
  assign n88 = n87 ^ x6 ;
  assign n89 = ~n85 & n88 ;
  assign n90 = n89 ^ x6 ;
  assign n91 = ~n82 & n90 ;
  assign n92 = n91 ^ x6 ;
  assign n93 = n51 & n92 ;
  assign n44 = ~x2 & ~x3 ;
  assign n94 = x1 & n44 ;
  assign n95 = n82 & n94 ;
  assign n96 = ~x1 & ~x4 ;
  assign n97 = x8 ^ x6 ;
  assign n98 = x8 ^ x2 ;
  assign n99 = ~n97 & ~n98 ;
  assign n100 = n96 & n99 ;
  assign n101 = ~x3 & n100 ;
  assign n102 = ~n95 & ~n101 ;
  assign n103 = ~n93 & n102 ;
  assign n104 = x0 & ~n103 ;
  assign n105 = x6 & ~x8 ;
  assign n106 = n94 & n105 ;
  assign n107 = x2 ^ x1 ;
  assign n108 = ~x0 & x8 ;
  assign n109 = n108 ^ n107 ;
  assign n110 = n86 ^ x3 ;
  assign n111 = x3 ^ x1 ;
  assign n112 = n111 ^ x3 ;
  assign n113 = ~n110 & n112 ;
  assign n114 = n113 ^ x3 ;
  assign n115 = n114 ^ n107 ;
  assign n116 = n109 & ~n115 ;
  assign n117 = n116 ^ n113 ;
  assign n118 = n117 ^ x3 ;
  assign n119 = n118 ^ n108 ;
  assign n120 = n107 & ~n119 ;
  assign n121 = n120 ^ n107 ;
  assign n122 = ~n106 & ~n121 ;
  assign n123 = x4 & ~n122 ;
  assign n124 = ~n104 & ~n123 ;
  assign n125 = ~n81 & n124 ;
  assign n64 = ~x2 & x3 ;
  assign n21 = n20 ^ x6 ;
  assign n22 = n20 ^ x4 ;
  assign n23 = n22 ^ x4 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = ~x3 & ~x4 ;
  assign n26 = ~x1 & x4 ;
  assign n27 = x0 & ~n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = ~n25 & ~n28 ;
  assign n30 = n29 ^ x4 ;
  assign n31 = n30 ^ n25 ;
  assign n32 = n24 & ~n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ n25 ;
  assign n35 = ~n21 & ~n34 ;
  assign n36 = x2 & n35 ;
  assign n37 = x3 ^ x0 ;
  assign n16 = ~x4 & x6 ;
  assign n38 = x0 & ~x2 ;
  assign n39 = ~x1 & n38 ;
  assign n40 = n16 & n39 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n41 ^ x3 ;
  assign n43 = n42 ^ n41 ;
  assign n45 = n26 & n44 ;
  assign n46 = x6 & n45 ;
  assign n47 = n46 ^ n41 ;
  assign n48 = n47 ^ n37 ;
  assign n49 = n43 & ~n48 ;
  assign n50 = n49 ^ n46 ;
  assign n52 = ~x4 & n51 ;
  assign n53 = ~n46 & ~n52 ;
  assign n54 = n53 ^ n37 ;
  assign n55 = ~n50 & n54 ;
  assign n56 = n55 ^ n53 ;
  assign n57 = n37 & n56 ;
  assign n58 = n57 ^ n49 ;
  assign n59 = n58 ^ x0 ;
  assign n60 = n59 ^ n46 ;
  assign n61 = ~n36 & ~n60 ;
  assign n65 = n64 ^ n61 ;
  assign n66 = n65 ^ n61 ;
  assign n17 = n16 ^ x6 ;
  assign n18 = x1 & ~n17 ;
  assign n19 = n18 ^ x6 ;
  assign n62 = n61 ^ n19 ;
  assign n63 = n62 ^ n61 ;
  assign n67 = n66 ^ n63 ;
  assign n68 = n61 ^ x0 ;
  assign n69 = n68 ^ n61 ;
  assign n70 = n69 ^ n66 ;
  assign n71 = n66 & ~n70 ;
  assign n72 = n71 ^ n66 ;
  assign n73 = ~n67 & n72 ;
  assign n74 = n73 ^ n71 ;
  assign n75 = n74 ^ n61 ;
  assign n76 = n75 ^ n66 ;
  assign n77 = x8 & ~n76 ;
  assign n78 = n77 ^ n61 ;
  assign n126 = n125 ^ n78 ;
  assign n127 = ~x5 & n126 ;
  assign n128 = n127 ^ n125 ;
  assign n129 = ~n15 & n128 ;
  assign n130 = x7 & ~n129 ;
  assign n131 = x0 & x3 ;
  assign n132 = ~x0 & x2 ;
  assign n133 = ~n131 & ~n132 ;
  assign n134 = ~n44 & n133 ;
  assign n135 = x5 & n10 ;
  assign n136 = n134 & n135 ;
  assign n137 = x2 & ~x7 ;
  assign n138 = n131 & n137 ;
  assign n139 = ~x5 & x8 ;
  assign n140 = ~n83 & ~n139 ;
  assign n141 = n138 & ~n140 ;
  assign n142 = ~x5 & ~x7 ;
  assign n143 = x0 & n142 ;
  assign n144 = n44 & n82 ;
  assign n145 = n143 & n144 ;
  assign n146 = ~n141 & ~n145 ;
  assign n147 = ~x0 & x5 ;
  assign n148 = n12 & n147 ;
  assign n149 = ~x7 & x8 ;
  assign n150 = x4 & n149 ;
  assign n151 = n148 & n150 ;
  assign n152 = x1 & ~n151 ;
  assign n153 = n146 & n152 ;
  assign n154 = ~n136 & n153 ;
  assign n155 = x6 & ~n154 ;
  assign n156 = x4 ^ x3 ;
  assign n157 = n156 ^ x8 ;
  assign n158 = x2 ^ x0 ;
  assign n159 = n158 ^ n157 ;
  assign n160 = x8 ^ x4 ;
  assign n161 = x4 ^ x2 ;
  assign n162 = n161 ^ x4 ;
  assign n163 = n160 & ~n162 ;
  assign n164 = n163 ^ x4 ;
  assign n165 = n164 ^ n157 ;
  assign n166 = ~n159 & n165 ;
  assign n167 = n166 ^ n163 ;
  assign n168 = n167 ^ x4 ;
  assign n169 = n168 ^ n158 ;
  assign n170 = ~n157 & ~n169 ;
  assign n171 = n170 ^ n157 ;
  assign n172 = n142 & ~n171 ;
  assign n173 = x5 & ~x8 ;
  assign n174 = x4 & n38 ;
  assign n175 = ~x3 & n174 ;
  assign n176 = ~n138 & ~n175 ;
  assign n177 = n173 & ~n176 ;
  assign n178 = ~x1 & ~n177 ;
  assign n179 = ~n172 & n178 ;
  assign n180 = n155 & ~n179 ;
  assign n181 = ~n143 & ~n147 ;
  assign n182 = n52 & ~n181 ;
  assign n183 = ~x4 & ~n142 ;
  assign n184 = n39 & ~n183 ;
  assign n185 = ~n182 & ~n184 ;
  assign n186 = x8 & ~n185 ;
  assign n187 = ~x2 & ~x4 ;
  assign n188 = ~x7 & n173 ;
  assign n189 = ~x0 & x1 ;
  assign n190 = n188 & n189 ;
  assign n191 = ~n187 & n190 ;
  assign n192 = ~n186 & ~n191 ;
  assign n193 = ~x6 & ~n192 ;
  assign n194 = x0 & n26 ;
  assign n195 = x8 ^ x5 ;
  assign n196 = x5 ^ x2 ;
  assign n197 = n195 & n196 ;
  assign n198 = n194 & n197 ;
  assign n199 = ~x7 & n198 ;
  assign n200 = ~n193 & ~n199 ;
  assign n201 = ~x3 & ~n200 ;
  assign n202 = x4 ^ x1 ;
  assign n203 = n131 ^ x4 ;
  assign n204 = n203 ^ n131 ;
  assign n205 = n204 ^ n202 ;
  assign n206 = x6 ^ x0 ;
  assign n207 = ~x6 & n206 ;
  assign n208 = n207 ^ n131 ;
  assign n209 = n208 ^ x6 ;
  assign n210 = ~n205 & ~n209 ;
  assign n211 = n210 ^ n207 ;
  assign n212 = n211 ^ x6 ;
  assign n213 = ~n202 & ~n212 ;
  assign n214 = n188 & n213 ;
  assign n215 = x2 & n214 ;
  assign n216 = ~n201 & ~n215 ;
  assign n217 = ~n180 & n216 ;
  assign n218 = ~n130 & n217 ;
  assign y0 = ~n218 ;
endmodule
