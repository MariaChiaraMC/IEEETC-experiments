module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 ;
  assign n59 = x6 ^ x3 ;
  assign n60 = n59 ^ x6 ;
  assign n61 = ~x6 & ~x7 ;
  assign n62 = n61 ^ x6 ;
  assign n63 = ~n60 & ~n62 ;
  assign n64 = n63 ^ x6 ;
  assign n65 = ~x5 & ~n64 ;
  assign n66 = n65 ^ x3 ;
  assign n67 = x4 & n66 ;
  assign n39 = ~x3 & x6 ;
  assign n68 = x2 & ~n39 ;
  assign n69 = n68 ^ x5 ;
  assign n70 = n69 ^ n68 ;
  assign n71 = x6 & x7 ;
  assign n72 = x3 & ~x4 ;
  assign n73 = ~n71 & n72 ;
  assign n74 = n73 ^ n68 ;
  assign n75 = ~n70 & ~n74 ;
  assign n76 = n75 ^ n68 ;
  assign n77 = ~n67 & n76 ;
  assign n78 = ~x1 & ~n77 ;
  assign n9 = ~x1 & x5 ;
  assign n15 = ~x4 & x7 ;
  assign n16 = ~x6 & n15 ;
  assign n17 = n9 & n16 ;
  assign n20 = x5 ^ x3 ;
  assign n21 = n20 ^ x6 ;
  assign n22 = n21 ^ x4 ;
  assign n18 = x7 ^ x5 ;
  assign n19 = n18 ^ x6 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n23 ^ n22 ;
  assign n27 = n18 ^ x7 ;
  assign n28 = n27 ^ n22 ;
  assign n29 = ~n22 & ~n28 ;
  assign n25 = ~n18 & ~n21 ;
  assign n32 = n29 ^ n25 ;
  assign n26 = n25 ^ n24 ;
  assign n30 = n29 ^ n22 ;
  assign n31 = ~n26 & ~n30 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = ~n24 & n33 ;
  assign n35 = n34 ^ n29 ;
  assign n36 = n35 ^ n31 ;
  assign n37 = n36 ^ n21 ;
  assign n38 = ~x1 & ~n37 ;
  assign n40 = n39 ^ x4 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = n41 ^ x1 ;
  assign n43 = ~x3 & ~x5 ;
  assign n44 = x3 & x5 ;
  assign n45 = x7 & n44 ;
  assign n46 = n45 ^ n43 ;
  assign n47 = ~n43 & n46 ;
  assign n48 = n47 ^ n39 ;
  assign n49 = n48 ^ n43 ;
  assign n50 = n42 & n49 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = n51 ^ n43 ;
  assign n53 = x1 & ~n52 ;
  assign n54 = n53 ^ x1 ;
  assign n55 = ~n38 & ~n54 ;
  assign n56 = ~n17 & n55 ;
  assign n57 = n56 ^ x2 ;
  assign n10 = ~x3 & n9 ;
  assign n11 = ~x2 & x4 ;
  assign n12 = ~n10 & ~n11 ;
  assign n13 = x7 & ~n12 ;
  assign n14 = n13 ^ x2 ;
  assign n58 = n57 ^ n14 ;
  assign n79 = n78 ^ n58 ;
  assign n80 = n79 ^ n58 ;
  assign n81 = n58 ^ n57 ;
  assign n82 = n81 ^ x2 ;
  assign n83 = ~n80 & ~n82 ;
  assign n84 = n83 ^ n57 ;
  assign n85 = x3 & ~x6 ;
  assign n86 = x1 & ~x5 ;
  assign n87 = ~n72 & ~n86 ;
  assign n88 = ~n39 & n87 ;
  assign n89 = ~n85 & n88 ;
  assign n90 = n57 & n89 ;
  assign n91 = n90 ^ x2 ;
  assign n92 = n84 & ~n91 ;
  assign n93 = n92 ^ n90 ;
  assign n94 = ~x2 & n93 ;
  assign n95 = n94 ^ n83 ;
  assign n96 = n95 ^ n56 ;
  assign n97 = n96 ^ n57 ;
  assign n98 = ~x0 & ~n97 ;
  assign y0 = n98 ;
endmodule
