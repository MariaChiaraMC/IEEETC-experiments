module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n7 = x0 & ~x3 ;
  assign n8 = x1 & ~x5 ;
  assign n9 = n7 & n8 ;
  assign n10 = ~x2 & n9 ;
  assign n11 = ~x3 & ~x4 ;
  assign n12 = x2 & ~n11 ;
  assign n13 = ~x1 & ~n12 ;
  assign n14 = ~x0 & x2 ;
  assign n15 = n11 & ~n14 ;
  assign n16 = n15 ^ x5 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = ~x0 & x4 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = n19 & n20 ;
  assign n22 = n21 ^ n15 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n18 & n23 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ n19 ;
  assign n27 = n13 & n26 ;
  assign n28 = n27 ^ n13 ;
  assign n29 = ~n10 & ~n28 ;
  assign y0 = ~n29 ;
endmodule
