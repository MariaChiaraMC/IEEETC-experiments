module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 ;
  assign n13 = ~x5 & ~x9 ;
  assign n14 = ~x11 & ~n13 ;
  assign n15 = ~x3 & ~x10 ;
  assign n16 = ~x0 & ~x1 ;
  assign n17 = n15 & n16 ;
  assign n18 = ~n14 & n17 ;
  assign n19 = n18 ^ x6 ;
  assign n20 = n19 ^ x6 ;
  assign n21 = x7 ^ x6 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n23 ^ x6 ;
  assign n25 = n24 ^ x6 ;
  assign n26 = n20 & n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n24 ^ x8 ;
  assign n29 = n28 ^ n27 ;
  assign n31 = x5 & x9 ;
  assign n30 = n22 ^ x0 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = n24 & ~n32 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = n29 & n35 ;
  assign n37 = n36 ^ n24 ;
  assign n38 = n27 & n37 ;
  assign n39 = n38 ^ n26 ;
  assign n40 = n39 ^ n24 ;
  assign n41 = n40 ^ n18 ;
  assign y0 = n41 ;
endmodule
