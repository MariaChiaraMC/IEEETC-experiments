module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 ;
  assign n9 = ~x6 & ~x7 ;
  assign n10 = ~x2 & ~x7 ;
  assign n11 = x6 & ~n10 ;
  assign n12 = n11 ^ x0 ;
  assign n13 = x1 ^ x0 ;
  assign n14 = n13 ^ x0 ;
  assign n15 = n12 & ~n14 ;
  assign n16 = n15 ^ x0 ;
  assign n17 = n16 ^ n9 ;
  assign n18 = n9 ^ x5 ;
  assign n19 = n18 ^ n9 ;
  assign n20 = n17 & ~n19 ;
  assign n21 = n20 ^ n15 ;
  assign n22 = n21 ^ x0 ;
  assign n23 = n22 ^ n18 ;
  assign n24 = ~n9 & ~n23 ;
  assign n25 = n24 ^ n9 ;
  assign n26 = n25 ^ n18 ;
  assign y0 = n26 ;
endmodule
