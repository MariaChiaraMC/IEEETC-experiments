module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 ;
  assign n11 = ~x4 & ~x9 ;
  assign n22 = ~x5 & ~x6 ;
  assign n23 = x2 & x3 ;
  assign n24 = x2 ^ x0 ;
  assign n25 = n24 ^ x3 ;
  assign n26 = n23 & n25 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = n22 & ~n27 ;
  assign n12 = ~x2 & ~x3 ;
  assign n13 = ~x0 & n12 ;
  assign n14 = ~x5 & n13 ;
  assign n15 = ~x6 & ~x7 ;
  assign n16 = x8 & n15 ;
  assign n17 = n14 & n16 ;
  assign n29 = n28 ^ n17 ;
  assign n30 = n29 ^ n17 ;
  assign n18 = x7 & n13 ;
  assign n19 = x5 & ~n18 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n20 ^ n17 ;
  assign n31 = n30 ^ n21 ;
  assign n32 = x8 ^ x6 ;
  assign n33 = x8 ^ x7 ;
  assign n34 = n33 ^ x7 ;
  assign n35 = n14 ^ x7 ;
  assign n36 = ~n34 & n35 ;
  assign n37 = n36 ^ x7 ;
  assign n38 = n32 & n37 ;
  assign n39 = n38 ^ x6 ;
  assign n40 = n39 ^ n17 ;
  assign n41 = n40 ^ n17 ;
  assign n42 = n41 ^ n30 ;
  assign n43 = ~n30 & n42 ;
  assign n44 = n43 ^ n30 ;
  assign n45 = n31 & ~n44 ;
  assign n46 = n45 ^ n43 ;
  assign n47 = n46 ^ n17 ;
  assign n48 = n47 ^ n30 ;
  assign n49 = ~x1 & ~n48 ;
  assign n50 = n49 ^ n17 ;
  assign n51 = n11 & n50 ;
  assign y0 = n51 ;
endmodule
