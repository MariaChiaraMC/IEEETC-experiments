module top( x0 , y0 );
  input x0 ;
  output y0 ;
  assign y0 = x0 ;
endmodule
