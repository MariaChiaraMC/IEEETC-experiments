module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 ;
  assign n17 = x8 & x9 ;
  assign n18 = ~x7 & n17 ;
  assign n19 = ~x0 & ~x1 ;
  assign n20 = ~x2 & n19 ;
  assign n21 = n18 & n20 ;
  assign n22 = ~x4 & x6 ;
  assign n23 = x5 & x10 ;
  assign n24 = ~x14 & x15 ;
  assign n25 = n23 & n24 ;
  assign n26 = n22 & n25 ;
  assign n27 = n21 & n26 ;
  assign n28 = ~x4 & ~x14 ;
  assign n29 = ~x7 & x15 ;
  assign n30 = n20 & n29 ;
  assign n31 = x10 ^ x6 ;
  assign n32 = n17 ^ x10 ;
  assign n33 = n32 ^ n17 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = ~x8 & ~x9 ;
  assign n36 = n35 ^ x5 ;
  assign n37 = ~x5 & ~n36 ;
  assign n38 = n37 ^ n17 ;
  assign n39 = n38 ^ x5 ;
  assign n40 = n34 & ~n39 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n41 ^ x5 ;
  assign n43 = ~n31 & ~n42 ;
  assign n44 = n30 & n43 ;
  assign n45 = n28 & n44 ;
  assign n46 = ~x10 & n22 ;
  assign n47 = x0 & ~x14 ;
  assign n48 = x9 ^ x7 ;
  assign n56 = n48 ^ x1 ;
  assign n49 = x8 ^ x1 ;
  assign n50 = n49 ^ n48 ;
  assign n51 = n50 ^ x1 ;
  assign n52 = n48 ^ x9 ;
  assign n53 = n52 ^ n49 ;
  assign n54 = n53 ^ n51 ;
  assign n55 = n51 & n54 ;
  assign n57 = n56 ^ n55 ;
  assign n58 = n57 ^ n51 ;
  assign n59 = x2 ^ x1 ;
  assign n60 = n55 ^ n51 ;
  assign n61 = ~n59 & n60 ;
  assign n62 = n61 ^ x1 ;
  assign n63 = ~n58 & n62 ;
  assign n64 = n63 ^ x1 ;
  assign n65 = n64 ^ x1 ;
  assign n66 = n47 & n65 ;
  assign n67 = n46 & n66 ;
  assign n68 = n67 ^ x5 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = n69 ^ x15 ;
  assign n71 = x7 & ~x14 ;
  assign n72 = n20 & n71 ;
  assign n73 = ~x6 & n72 ;
  assign n74 = x8 ^ x4 ;
  assign n75 = x10 ^ x8 ;
  assign n76 = n75 ^ x10 ;
  assign n77 = ~x9 & x10 ;
  assign n78 = n77 ^ x10 ;
  assign n79 = ~n76 & ~n78 ;
  assign n80 = n79 ^ x10 ;
  assign n81 = n74 & ~n80 ;
  assign n82 = n73 & n81 ;
  assign n83 = ~x8 & x9 ;
  assign n84 = x2 & ~x6 ;
  assign n85 = n83 & n84 ;
  assign n86 = x4 & n19 ;
  assign n87 = x10 & x14 ;
  assign n88 = n86 & n87 ;
  assign n89 = n85 & n88 ;
  assign n90 = ~n82 & ~n89 ;
  assign n91 = x2 & x9 ;
  assign n92 = x8 & ~x10 ;
  assign n93 = n22 & n92 ;
  assign n94 = x0 & x1 ;
  assign n95 = n71 & n94 ;
  assign n96 = n93 & n95 ;
  assign n97 = n91 & n96 ;
  assign n98 = n97 ^ n90 ;
  assign n99 = n90 & ~n98 ;
  assign n100 = n99 ^ n67 ;
  assign n101 = n100 ^ n90 ;
  assign n102 = ~n70 & ~n101 ;
  assign n103 = n102 ^ n99 ;
  assign n104 = n103 ^ n90 ;
  assign n105 = ~x15 & n104 ;
  assign n106 = n105 ^ x15 ;
  assign n107 = ~n45 & n106 ;
  assign n108 = n107 ^ x3 ;
  assign n109 = n108 ^ n107 ;
  assign n110 = x6 & ~x14 ;
  assign n111 = x4 & x7 ;
  assign n112 = ~x2 & n111 ;
  assign n113 = x9 & x10 ;
  assign n114 = ~x0 & ~n113 ;
  assign n115 = x9 ^ x8 ;
  assign n116 = n115 ^ x9 ;
  assign n117 = x10 & ~x15 ;
  assign n118 = n117 ^ x9 ;
  assign n119 = n116 & n118 ;
  assign n120 = n119 ^ x9 ;
  assign n121 = x1 & n120 ;
  assign n122 = n114 & n121 ;
  assign n123 = n112 & n122 ;
  assign n124 = n110 & n123 ;
  assign n125 = ~x1 & n110 ;
  assign n126 = ~x4 & n92 ;
  assign n127 = x0 & ~x15 ;
  assign n128 = n48 & n127 ;
  assign n129 = n126 & n128 ;
  assign n130 = ~x0 & ~x8 ;
  assign n131 = n112 & n130 ;
  assign n132 = n77 & n131 ;
  assign n133 = ~n129 & ~n132 ;
  assign n134 = n125 & ~n133 ;
  assign n135 = ~n124 & ~n134 ;
  assign n136 = ~x1 & x7 ;
  assign n137 = x10 & x15 ;
  assign n138 = n136 & n137 ;
  assign n139 = n130 & n138 ;
  assign n140 = n139 ^ x6 ;
  assign n141 = n140 ^ n139 ;
  assign n142 = ~x10 & n128 ;
  assign n143 = ~n83 & n142 ;
  assign n144 = n143 ^ n139 ;
  assign n145 = n141 & n144 ;
  assign n146 = n145 ^ n139 ;
  assign n147 = n28 & n146 ;
  assign n148 = ~x0 & ~n83 ;
  assign n149 = x4 & ~n148 ;
  assign n150 = ~x6 & x14 ;
  assign n151 = ~x0 & ~n87 ;
  assign n152 = x7 & ~n151 ;
  assign n153 = ~n150 & ~n152 ;
  assign n154 = n153 ^ n149 ;
  assign n155 = ~n17 & ~n35 ;
  assign n156 = ~x15 & n125 ;
  assign n157 = ~n155 & n156 ;
  assign n158 = n157 ^ x0 ;
  assign n159 = n158 ^ n157 ;
  assign n160 = n157 ^ x1 ;
  assign n161 = ~n159 & n160 ;
  assign n162 = n161 ^ n157 ;
  assign n163 = n162 ^ n149 ;
  assign n164 = ~n154 & n163 ;
  assign n165 = n164 ^ n161 ;
  assign n166 = n165 ^ n157 ;
  assign n167 = n166 ^ n153 ;
  assign n168 = n149 & ~n167 ;
  assign n169 = n168 ^ n149 ;
  assign n170 = ~n147 & ~n169 ;
  assign n171 = n170 ^ x2 ;
  assign n172 = n171 ^ n170 ;
  assign n173 = n172 ^ n135 ;
  assign n174 = x6 & x15 ;
  assign n175 = n94 & n174 ;
  assign n176 = n175 ^ n111 ;
  assign n177 = n111 & n176 ;
  assign n178 = n177 ^ n170 ;
  assign n179 = n178 ^ n111 ;
  assign n180 = ~n173 & ~n179 ;
  assign n181 = n180 ^ n177 ;
  assign n182 = n181 ^ n111 ;
  assign n183 = n135 & n182 ;
  assign n184 = n183 ^ n135 ;
  assign n185 = ~x5 & ~n184 ;
  assign n186 = ~x7 & x9 ;
  assign n187 = x6 & x10 ;
  assign n188 = x14 & ~n187 ;
  assign n189 = n188 ^ n110 ;
  assign n190 = n189 ^ n188 ;
  assign n191 = x5 & n117 ;
  assign n192 = n191 ^ n188 ;
  assign n193 = n192 ^ n188 ;
  assign n194 = n190 & n193 ;
  assign n195 = n194 ^ n188 ;
  assign n196 = ~x1 & n195 ;
  assign n197 = n196 ^ n188 ;
  assign n198 = x4 & n197 ;
  assign n199 = x2 & ~n198 ;
  assign n200 = n186 & ~n199 ;
  assign n201 = ~x4 & x5 ;
  assign n202 = x14 & ~x15 ;
  assign n203 = x7 & ~x9 ;
  assign n204 = ~x1 & x6 ;
  assign n205 = n203 & n204 ;
  assign n206 = n202 & n205 ;
  assign n207 = n201 & n206 ;
  assign n208 = ~x10 & n207 ;
  assign n209 = ~n200 & ~n208 ;
  assign n210 = ~x6 & ~x10 ;
  assign n211 = ~x14 & ~x15 ;
  assign n212 = n210 & n211 ;
  assign n213 = ~x1 & n186 ;
  assign n214 = n212 & n213 ;
  assign n215 = n201 & n214 ;
  assign n216 = ~x2 & ~n215 ;
  assign n217 = n130 & ~n216 ;
  assign n218 = ~n209 & n217 ;
  assign n219 = ~n185 & ~n218 ;
  assign n220 = n219 ^ n107 ;
  assign n221 = n109 & n220 ;
  assign n222 = n221 ^ n107 ;
  assign n223 = ~n27 & n222 ;
  assign n224 = ~x13 & ~n223 ;
  assign n225 = ~x3 & n23 ;
  assign n226 = x14 ^ x13 ;
  assign n227 = n226 ^ x13 ;
  assign n228 = x13 ^ x11 ;
  assign n229 = n227 & n228 ;
  assign n230 = n229 ^ x13 ;
  assign n231 = ~x15 & n230 ;
  assign n232 = n86 & n231 ;
  assign n233 = n85 & n232 ;
  assign n234 = n225 & n233 ;
  assign n235 = ~n224 & ~n234 ;
  assign n236 = ~x12 & ~n235 ;
  assign y0 = n236 ;
endmodule
