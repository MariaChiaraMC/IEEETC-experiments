module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 ;
  assign n65 = ~x1 & x6 ;
  assign n66 = ~x4 & ~n65 ;
  assign n9 = x1 & ~x6 ;
  assign n10 = x4 & ~n9 ;
  assign n11 = x2 ^ x0 ;
  assign n12 = x3 ^ x2 ;
  assign n13 = n11 & n12 ;
  assign n15 = x1 & ~x5 ;
  assign n14 = x5 & ~x6 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n15 ^ x3 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = ~n16 & n19 ;
  assign n21 = n20 ^ n14 ;
  assign n22 = n13 & n21 ;
  assign n23 = n10 & n22 ;
  assign n24 = ~x0 & x2 ;
  assign n25 = x3 & ~x4 ;
  assign n26 = n24 & n25 ;
  assign n27 = x1 & ~x3 ;
  assign n28 = ~x2 & n27 ;
  assign n29 = ~n26 & ~n28 ;
  assign n30 = x4 ^ x0 ;
  assign n37 = n30 ^ x6 ;
  assign n38 = n37 ^ x0 ;
  assign n31 = n30 ^ x1 ;
  assign n32 = n31 ^ x5 ;
  assign n39 = n38 ^ n32 ;
  assign n40 = n39 ^ x5 ;
  assign n41 = ~x5 & ~n40 ;
  assign n42 = n41 ^ n30 ;
  assign n43 = n42 ^ n32 ;
  assign n44 = n43 ^ x5 ;
  assign n45 = n44 ^ x0 ;
  assign n46 = n32 ^ x5 ;
  assign n47 = n46 ^ x0 ;
  assign n48 = ~n43 & ~n47 ;
  assign n49 = n48 ^ n30 ;
  assign n50 = n49 ^ n32 ;
  assign n51 = n50 ^ x5 ;
  assign n52 = n51 ^ x0 ;
  assign n53 = n45 & n52 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ x5 ;
  assign n35 = n34 ^ x0 ;
  assign n36 = n34 & n35 ;
  assign n54 = n53 ^ n36 ;
  assign n55 = n54 ^ n41 ;
  assign n56 = n55 ^ n30 ;
  assign n57 = n56 ^ n32 ;
  assign n58 = n57 ^ x5 ;
  assign n59 = n58 ^ x0 ;
  assign n60 = ~n29 & n59 ;
  assign n61 = ~n23 & ~n60 ;
  assign n67 = n66 ^ n61 ;
  assign n68 = n67 ^ n61 ;
  assign n62 = ~x0 & ~x5 ;
  assign n63 = n62 ^ n61 ;
  assign n64 = n63 ^ n61 ;
  assign n69 = n68 ^ n64 ;
  assign n70 = x2 & ~n10 ;
  assign n71 = x3 & n70 ;
  assign n72 = n71 ^ n61 ;
  assign n73 = n72 ^ n61 ;
  assign n74 = n73 ^ n68 ;
  assign n75 = ~n68 & ~n74 ;
  assign n76 = n75 ^ n68 ;
  assign n77 = ~n69 & ~n76 ;
  assign n78 = n77 ^ n75 ;
  assign n79 = n78 ^ n61 ;
  assign n80 = n79 ^ n68 ;
  assign n81 = x7 & n80 ;
  assign n82 = n81 ^ n61 ;
  assign y0 = ~n82 ;
endmodule
