module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n11 = x4 & x5 ;
  assign n12 = ~x3 & ~x6 ;
  assign n13 = ~n11 & n12 ;
  assign n17 = ~x4 & ~x5 ;
  assign n14 = ~x0 & ~x2 ;
  assign n15 = ~x8 & n14 ;
  assign n16 = ~x7 & n15 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = n18 ^ x1 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = n20 ^ n13 ;
  assign n22 = x7 & ~x9 ;
  assign n23 = ~x8 & ~n22 ;
  assign n24 = x2 ^ x0 ;
  assign n25 = ~n23 & n24 ;
  assign n26 = n25 ^ x1 ;
  assign n27 = n25 & ~n26 ;
  assign n28 = n27 ^ n16 ;
  assign n29 = n28 ^ n25 ;
  assign n30 = n21 & n29 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n31 ^ n25 ;
  assign n33 = n13 & n32 ;
  assign y0 = n33 ;
endmodule
