module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n15 = x6 & ~x7 ;
  assign n16 = ~x1 & ~x2 ;
  assign n17 = x4 & x5 ;
  assign n18 = n16 & n17 ;
  assign n19 = ~x0 & ~x3 ;
  assign n20 = x9 & n19 ;
  assign n21 = n18 & n20 ;
  assign n22 = n15 & n21 ;
  assign n23 = x10 & x11 ;
  assign n24 = n23 ^ x8 ;
  assign n25 = x12 & x13 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n24 & ~n26 ;
  assign n28 = n27 ^ x8 ;
  assign n29 = n22 & n28 ;
  assign y0 = n29 ;
endmodule
