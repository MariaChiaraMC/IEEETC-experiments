module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n8 = ~x3 & ~x5 ;
  assign n9 = x4 & x6 ;
  assign n10 = ~x3 & ~n9 ;
  assign n11 = x2 & ~n10 ;
  assign n12 = ~n8 & n11 ;
  assign n13 = ~x1 & ~n12 ;
  assign n14 = ~x0 & ~n13 ;
  assign n15 = x4 ^ x2 ;
  assign n16 = x2 ^ x0 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n8 ^ x4 ;
  assign n19 = n18 ^ n8 ;
  assign n20 = x1 & x3 ;
  assign n21 = n20 ^ n8 ;
  assign n22 = n19 & n21 ;
  assign n23 = n22 ^ n8 ;
  assign n24 = n23 ^ n15 ;
  assign n25 = n17 & ~n24 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = n26 ^ n8 ;
  assign n28 = n27 ^ n16 ;
  assign n29 = ~n15 & ~n28 ;
  assign n30 = n29 ^ n15 ;
  assign n31 = n30 ^ x0 ;
  assign n32 = ~n14 & n31 ;
  assign y0 = ~n32 ;
endmodule
