module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n10 = x4 ^ x2 ;
  assign n9 = x7 ^ x4 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = n12 ^ x4 ;
  assign n14 = x5 ^ x4 ;
  assign n15 = x6 ^ x4 ;
  assign n16 = ~n14 & ~n15 ;
  assign n17 = n10 ^ x4 ;
  assign n18 = ~n12 & n17 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = n16 & ~n19 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = ~n13 & n21 ;
  assign n23 = n22 ^ n18 ;
  assign n24 = n23 ^ x4 ;
  assign n25 = ~x3 & ~n24 ;
  assign n26 = x4 & ~x5 ;
  assign n27 = x6 ^ x2 ;
  assign n28 = x6 ^ x3 ;
  assign n29 = n28 ^ x6 ;
  assign n30 = ~n27 & n29 ;
  assign n31 = n30 ^ x6 ;
  assign n32 = n26 & ~n31 ;
  assign n33 = ~x1 & ~n32 ;
  assign n34 = ~n25 & n33 ;
  assign y0 = ~n34 ;
endmodule
