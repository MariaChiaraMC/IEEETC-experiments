module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 ;
  assign n11 = ~x1 & ~x6 ;
  assign n109 = ~x3 & x5 ;
  assign n110 = n11 & ~n109 ;
  assign n111 = x3 & ~x5 ;
  assign n112 = x7 & ~n111 ;
  assign n113 = n110 & n112 ;
  assign n10 = ~x5 & ~x7 ;
  assign n114 = ~x3 & x6 ;
  assign n115 = n10 & n114 ;
  assign n116 = x1 & n115 ;
  assign n117 = ~n113 & ~n116 ;
  assign n118 = ~x2 & x4 ;
  assign n119 = ~n117 & n118 ;
  assign n9 = x1 & x5 ;
  assign n12 = n10 & n11 ;
  assign n13 = ~n9 & ~n12 ;
  assign n14 = x3 & ~n13 ;
  assign n15 = ~x4 & n14 ;
  assign n19 = x5 ^ x4 ;
  assign n20 = n19 ^ x6 ;
  assign n16 = x3 ^ x1 ;
  assign n17 = n16 ^ x6 ;
  assign n18 = n17 ^ n16 ;
  assign n21 = n20 ^ n18 ;
  assign n23 = x5 ^ x3 ;
  assign n28 = n23 ^ x7 ;
  assign n22 = n16 ^ x5 ;
  assign n24 = n23 ^ n22 ;
  assign n29 = n28 ^ n24 ;
  assign n30 = n29 ^ n23 ;
  assign n36 = n30 ^ n16 ;
  assign n37 = n36 ^ n18 ;
  assign n32 = n23 ^ n18 ;
  assign n25 = n24 ^ n20 ;
  assign n26 = n25 ^ n16 ;
  assign n33 = n32 ^ n26 ;
  assign n34 = n33 ^ n16 ;
  assign n38 = n37 ^ n34 ;
  assign n27 = n26 ^ n18 ;
  assign n31 = n30 ^ n27 ;
  assign n35 = n34 ^ n31 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = ~n21 & n39 ;
  assign n41 = n40 ^ n30 ;
  assign n42 = n41 ^ n27 ;
  assign n43 = n42 ^ n21 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = n21 ^ n18 ;
  assign n46 = n27 ^ n18 ;
  assign n47 = n46 ^ n21 ;
  assign n48 = n47 ^ n34 ;
  assign n49 = n45 & ~n48 ;
  assign n50 = n49 ^ n38 ;
  assign n51 = n30 ^ n18 ;
  assign n52 = n51 ^ n27 ;
  assign n53 = n52 ^ n34 ;
  assign n54 = n35 & ~n53 ;
  assign n55 = n54 ^ n30 ;
  assign n56 = n55 ^ n18 ;
  assign n57 = n56 ^ n34 ;
  assign n58 = n57 ^ n38 ;
  assign n59 = n50 & ~n58 ;
  assign n60 = n59 ^ n30 ;
  assign n61 = n60 ^ n21 ;
  assign n62 = n61 ^ n34 ;
  assign n63 = n62 ^ n38 ;
  assign n64 = n44 & ~n63 ;
  assign n65 = n64 ^ n49 ;
  assign n66 = n65 ^ n18 ;
  assign n67 = n66 ^ n27 ;
  assign n68 = n67 ^ n26 ;
  assign n69 = n68 ^ x2 ;
  assign n70 = n69 ^ n68 ;
  assign n76 = x5 ^ x1 ;
  assign n71 = x4 ^ x1 ;
  assign n72 = n71 ^ x5 ;
  assign n77 = n76 ^ n72 ;
  assign n82 = n77 ^ n72 ;
  assign n73 = n72 ^ n16 ;
  assign n74 = n73 ^ x1 ;
  assign n75 = n74 ^ x1 ;
  assign n78 = n77 ^ n74 ;
  assign n79 = n78 ^ x1 ;
  assign n80 = ~n75 & n79 ;
  assign n81 = n80 ^ n77 ;
  assign n83 = n82 ^ n81 ;
  assign n84 = x6 ^ x1 ;
  assign n85 = n84 ^ x1 ;
  assign n86 = n85 ^ n82 ;
  assign n87 = n85 ^ n78 ;
  assign n88 = ~n86 & ~n87 ;
  assign n89 = n88 ^ n74 ;
  assign n90 = n89 ^ n77 ;
  assign n91 = n90 ^ x1 ;
  assign n92 = x4 & ~x7 ;
  assign n93 = n92 ^ n74 ;
  assign n94 = n93 ^ n77 ;
  assign n95 = ~n85 & n94 ;
  assign n96 = n95 ^ n74 ;
  assign n97 = n96 ^ x1 ;
  assign n98 = n91 & ~n97 ;
  assign n99 = n98 ^ n77 ;
  assign n100 = n99 ^ x1 ;
  assign n101 = n100 ^ n82 ;
  assign n102 = ~n83 & ~n101 ;
  assign n103 = n102 ^ n80 ;
  assign n104 = n103 ^ n72 ;
  assign n105 = n104 ^ n68 ;
  assign n106 = n70 & ~n105 ;
  assign n107 = n106 ^ n68 ;
  assign n108 = ~n15 & ~n107 ;
  assign n120 = n119 ^ n108 ;
  assign n121 = x0 & ~n120 ;
  assign n122 = n121 ^ n108 ;
  assign y0 = ~n122 ;
endmodule
