// Benchmark "./mlp4.pla" written by ABC on Thu Apr 23 10:59:56 2020

module \./mlp4.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z7  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z7;
  assign z7 = 1'b1;
endmodule


