// Benchmark "./p82.pla" written by ABC on Thu Apr 23 11:00:00 2020

module \./p82.pla  ( 
    x0, x1, x2, x3, x4,
    z10  );
  input  x0, x1, x2, x3, x4;
  output z10;
  assign z10 = 1'b1;
endmodule


