module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 ;
  assign n9 = ~x2 & ~x5 ;
  assign n10 = ~x3 & ~n9 ;
  assign n11 = x3 & n9 ;
  assign n12 = n11 ^ x2 ;
  assign n13 = n12 ^ x4 ;
  assign n14 = x6 ^ x2 ;
  assign n15 = x7 ^ x5 ;
  assign n16 = x4 ^ x2 ;
  assign n17 = ~n15 & n16 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n14 & n19 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = ~n13 & ~n21 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = ~x4 & n23 ;
  assign n25 = ~n10 & n24 ;
  assign n34 = x3 ^ x2 ;
  assign n28 = x5 ^ x3 ;
  assign n29 = n28 ^ x2 ;
  assign n26 = n15 ^ x5 ;
  assign n27 = n26 ^ x2 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n29 ^ x2 ;
  assign n32 = ~n30 & n31 ;
  assign n33 = n32 ^ n29 ;
  assign n35 = n34 ^ n33 ;
  assign n36 = x4 ^ x3 ;
  assign n37 = n36 ^ x3 ;
  assign n38 = n37 ^ x2 ;
  assign n39 = n38 ^ x2 ;
  assign n40 = n39 ^ n26 ;
  assign n41 = n40 ^ n34 ;
  assign n42 = ~n40 & n41 ;
  assign n43 = n42 ^ x2 ;
  assign n44 = n43 ^ n38 ;
  assign n46 = n36 ^ x6 ;
  assign n47 = n46 ^ n36 ;
  assign n45 = n38 ^ n29 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = n38 & ~n48 ;
  assign n50 = n49 ^ x2 ;
  assign n51 = n50 ^ n29 ;
  assign n52 = n51 ^ n34 ;
  assign n53 = n44 & ~n52 ;
  assign n54 = n53 ^ x2 ;
  assign n55 = ~n35 & n54 ;
  assign n56 = n55 ^ n32 ;
  assign n57 = n56 ^ n29 ;
  assign n58 = n57 ^ x3 ;
  assign n59 = n58 ^ n34 ;
  assign n60 = ~n25 & ~n59 ;
  assign y0 = ~n60 ;
endmodule
