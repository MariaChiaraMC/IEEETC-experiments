module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 ;
  assign n7 = x3 ^ x2 ;
  assign n13 = n7 ^ x4 ;
  assign n10 = x4 ^ x1 ;
  assign n11 = n10 ^ x5 ;
  assign n8 = x5 ^ x2 ;
  assign n9 = n8 ^ n7 ;
  assign n12 = n11 ^ n9 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = n15 ^ n7 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n17 ^ x2 ;
  assign n19 = n18 ^ n11 ;
  assign n20 = n19 ^ n7 ;
  assign n21 = n20 ^ x2 ;
  assign n27 = n21 ^ x2 ;
  assign n28 = n27 ^ n16 ;
  assign n29 = n28 ^ n18 ;
  assign n30 = ~n16 & n29 ;
  assign n22 = n21 ^ n16 ;
  assign n23 = n16 ^ n7 ;
  assign n24 = n23 ^ n16 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = ~n22 & n25 ;
  assign n31 = n30 ^ n26 ;
  assign n32 = n31 ^ n16 ;
  assign n33 = n32 ^ n21 ;
  assign n34 = n27 ^ n21 ;
  assign n35 = n26 ^ n23 ;
  assign n36 = n35 ^ n21 ;
  assign n37 = n34 & ~n36 ;
  assign n38 = n37 ^ n26 ;
  assign n39 = n38 ^ n16 ;
  assign n40 = n39 ^ n27 ;
  assign n41 = n40 ^ n18 ;
  assign n42 = ~n33 & n41 ;
  assign n43 = n42 ^ n37 ;
  assign n44 = ~x0 & n43 ;
  assign n45 = x1 & ~x2 ;
  assign n46 = x5 & n45 ;
  assign n47 = x1 & ~x5 ;
  assign n48 = ~x1 & x5 ;
  assign n49 = ~n47 & ~n48 ;
  assign n50 = x4 & ~n49 ;
  assign n51 = x3 & ~n50 ;
  assign n52 = n7 ^ x2 ;
  assign n53 = n52 ^ x0 ;
  assign n54 = ~x1 & ~x5 ;
  assign n55 = n54 ^ x5 ;
  assign n56 = x2 & ~n55 ;
  assign n57 = n56 ^ x5 ;
  assign n58 = ~n53 & n57 ;
  assign n59 = n58 ^ n56 ;
  assign n60 = n59 ^ x5 ;
  assign n61 = n60 ^ x2 ;
  assign n62 = x0 & n61 ;
  assign n63 = ~n51 & n62 ;
  assign n64 = ~n46 & ~n63 ;
  assign n65 = ~n44 & n64 ;
  assign y0 = n65 ;
endmodule
