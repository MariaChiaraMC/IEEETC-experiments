module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n13 = x2 & x3 ;
  assign n14 = x9 & ~n13 ;
  assign n15 = ~x7 & ~n14 ;
  assign n16 = x0 & x1 ;
  assign n17 = x5 & ~x6 ;
  assign n18 = ~x11 & n17 ;
  assign n19 = n16 & n18 ;
  assign n20 = ~n15 & n19 ;
  assign n21 = x8 & x9 ;
  assign n22 = ~x3 & ~x10 ;
  assign n23 = ~x2 & ~n22 ;
  assign n24 = x7 & ~n23 ;
  assign n25 = n21 & n24 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = x7 & ~n13 ;
  assign n29 = ~x8 & ~n28 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = n27 & n30 ;
  assign n32 = n31 ^ n25 ;
  assign n33 = n20 & n32 ;
  assign y0 = n33 ;
endmodule
