module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 ;
  assign n11 = x2 & ~x4 ;
  assign n12 = x5 & ~x6 ;
  assign n15 = n12 ^ x3 ;
  assign n16 = n15 ^ n12 ;
  assign n13 = n12 ^ x1 ;
  assign n14 = n13 ^ n12 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = x9 ^ x8 ;
  assign n19 = n12 ^ x9 ;
  assign n20 = n19 ^ n12 ;
  assign n21 = ~x5 & x6 ;
  assign n22 = n21 ^ n12 ;
  assign n23 = n22 ^ n12 ;
  assign n24 = ~n20 & n23 ;
  assign n25 = n24 ^ n12 ;
  assign n26 = ~n18 & n25 ;
  assign n27 = n26 ^ n12 ;
  assign n28 = n27 ^ n12 ;
  assign n29 = n28 ^ n12 ;
  assign n30 = n29 ^ n16 ;
  assign n31 = ~n16 & ~n30 ;
  assign n32 = n31 ^ n16 ;
  assign n33 = n17 & ~n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n34 ^ n12 ;
  assign n36 = n35 ^ n16 ;
  assign n37 = ~x7 & ~n36 ;
  assign n38 = n37 ^ n12 ;
  assign n39 = n11 & n38 ;
  assign n40 = ~x3 & x4 ;
  assign n41 = x2 & n40 ;
  assign n42 = ~x3 & x6 ;
  assign n43 = ~x8 & ~x9 ;
  assign n44 = n42 & n43 ;
  assign n45 = ~x2 & n44 ;
  assign n46 = ~x0 & ~x2 ;
  assign n47 = ~x3 & ~x6 ;
  assign n48 = x8 & x9 ;
  assign n49 = n48 ^ x6 ;
  assign n50 = n49 ^ x8 ;
  assign n51 = ~n47 & ~n50 ;
  assign n52 = n51 ^ x8 ;
  assign n53 = n46 & n52 ;
  assign n54 = ~n45 & ~n53 ;
  assign n55 = ~x7 & ~n54 ;
  assign n56 = ~x6 & ~x7 ;
  assign n57 = ~x7 & x8 ;
  assign n58 = ~x3 & n57 ;
  assign n59 = ~n56 & ~n58 ;
  assign n60 = x3 & ~x6 ;
  assign n61 = x9 & ~n60 ;
  assign n62 = x8 & ~x9 ;
  assign n63 = x3 & n62 ;
  assign n64 = n63 ^ x8 ;
  assign n65 = ~n61 & n64 ;
  assign n66 = ~x0 & n65 ;
  assign n67 = ~n59 & ~n66 ;
  assign n68 = x2 & ~n67 ;
  assign n69 = ~x8 & x9 ;
  assign n70 = ~x3 & n56 ;
  assign n71 = n69 & n70 ;
  assign n72 = ~n68 & ~n71 ;
  assign n73 = ~n55 & n72 ;
  assign n74 = ~x5 & n73 ;
  assign n96 = x2 & x5 ;
  assign n75 = ~x9 & n60 ;
  assign n76 = n75 ^ x9 ;
  assign n77 = n76 ^ x2 ;
  assign n85 = n77 ^ n76 ;
  assign n78 = x2 & n47 ;
  assign n79 = n78 ^ n77 ;
  assign n80 = n79 ^ n76 ;
  assign n81 = n77 ^ n75 ;
  assign n82 = n81 ^ n78 ;
  assign n83 = n82 ^ n80 ;
  assign n84 = ~n80 & ~n83 ;
  assign n86 = n85 ^ n84 ;
  assign n87 = n86 ^ n80 ;
  assign n88 = n76 ^ x0 ;
  assign n89 = n84 ^ n80 ;
  assign n90 = n88 & ~n89 ;
  assign n91 = n90 ^ n76 ;
  assign n92 = ~n87 & n91 ;
  assign n93 = n92 ^ n76 ;
  assign n94 = n93 ^ x9 ;
  assign n95 = n94 ^ n76 ;
  assign n97 = n96 ^ n95 ;
  assign n98 = n97 ^ n57 ;
  assign n105 = n98 ^ n97 ;
  assign n99 = n98 ^ n12 ;
  assign n100 = n99 ^ n97 ;
  assign n101 = n98 ^ n95 ;
  assign n102 = n101 ^ n12 ;
  assign n103 = n102 ^ n100 ;
  assign n104 = n100 & n103 ;
  assign n106 = n105 ^ n104 ;
  assign n107 = n106 ^ n100 ;
  assign n108 = x3 & ~x7 ;
  assign n109 = n108 ^ n97 ;
  assign n110 = n104 ^ n100 ;
  assign n111 = ~n109 & n110 ;
  assign n112 = n111 ^ n97 ;
  assign n113 = n107 & ~n112 ;
  assign n114 = n113 ^ n97 ;
  assign n115 = n114 ^ n96 ;
  assign n116 = n115 ^ n97 ;
  assign n117 = ~n74 & ~n116 ;
  assign n118 = ~x4 & ~n117 ;
  assign n119 = x1 & ~n118 ;
  assign n120 = ~n41 & n119 ;
  assign n121 = n120 ^ n39 ;
  assign n122 = ~x2 & ~x5 ;
  assign n123 = ~x7 & ~n43 ;
  assign n124 = x3 & ~n49 ;
  assign n125 = n123 & ~n124 ;
  assign n126 = n122 & ~n125 ;
  assign n127 = ~x5 & ~x6 ;
  assign n128 = ~x5 & x7 ;
  assign n129 = x2 & ~n128 ;
  assign n130 = ~n127 & n129 ;
  assign n131 = ~n126 & ~n130 ;
  assign n132 = ~x4 & ~n131 ;
  assign n133 = ~n62 & ~n69 ;
  assign n134 = n78 & ~n133 ;
  assign n135 = ~x7 & n40 ;
  assign n136 = n127 & n135 ;
  assign n137 = ~x1 & ~n136 ;
  assign n138 = ~n134 & n137 ;
  assign n139 = ~n132 & n138 ;
  assign n140 = x5 & x6 ;
  assign n141 = n140 ^ x2 ;
  assign n142 = n141 ^ n140 ;
  assign n143 = n142 ^ x4 ;
  assign n144 = x7 ^ x5 ;
  assign n145 = x7 & ~n144 ;
  assign n146 = n145 ^ n140 ;
  assign n147 = n146 ^ x7 ;
  assign n148 = n143 & n147 ;
  assign n149 = n148 ^ n145 ;
  assign n150 = n149 ^ x7 ;
  assign n151 = ~x4 & n150 ;
  assign n152 = ~n139 & ~n151 ;
  assign n153 = ~n41 & n152 ;
  assign n154 = n153 ^ x0 ;
  assign n155 = n154 ^ n153 ;
  assign n156 = n42 & n96 ;
  assign n157 = x3 & n140 ;
  assign n158 = n133 ^ x5 ;
  assign n159 = n158 ^ n133 ;
  assign n160 = n133 ^ n43 ;
  assign n161 = ~n159 & ~n160 ;
  assign n162 = n161 ^ n133 ;
  assign n163 = ~x7 & n162 ;
  assign n164 = n60 & ~n163 ;
  assign n167 = ~n57 & ~n108 ;
  assign n168 = ~x9 & ~n167 ;
  assign n165 = n62 & n128 ;
  assign n166 = ~x3 & ~n165 ;
  assign n169 = n168 ^ n166 ;
  assign n170 = ~n21 & ~n169 ;
  assign n171 = n170 ^ n168 ;
  assign n172 = ~n164 & n171 ;
  assign n173 = n172 ^ x5 ;
  assign n174 = n173 ^ x2 ;
  assign n182 = n174 ^ n173 ;
  assign n175 = n57 & n60 ;
  assign n176 = n175 ^ n174 ;
  assign n177 = n176 ^ n173 ;
  assign n178 = n174 ^ n172 ;
  assign n179 = n178 ^ n175 ;
  assign n180 = n179 ^ n177 ;
  assign n181 = n177 & n180 ;
  assign n183 = n182 ^ n181 ;
  assign n184 = n183 ^ n177 ;
  assign n185 = x8 & n47 ;
  assign n186 = ~x7 & ~n185 ;
  assign n187 = n60 ^ x9 ;
  assign n188 = ~n42 & ~n187 ;
  assign n189 = ~x8 & n188 ;
  assign n190 = n186 & ~n189 ;
  assign n191 = n190 ^ n173 ;
  assign n192 = n181 ^ n177 ;
  assign n193 = n191 & n192 ;
  assign n194 = n193 ^ n173 ;
  assign n195 = ~n184 & n194 ;
  assign n196 = n195 ^ n173 ;
  assign n197 = n196 ^ x5 ;
  assign n198 = n197 ^ n173 ;
  assign n199 = ~n157 & n198 ;
  assign n200 = n199 ^ x1 ;
  assign n201 = n200 ^ n199 ;
  assign n202 = x8 ^ x3 ;
  assign n203 = n202 ^ x3 ;
  assign n204 = x7 ^ x3 ;
  assign n205 = n204 ^ x3 ;
  assign n206 = ~n203 & ~n205 ;
  assign n207 = n206 ^ x3 ;
  assign n208 = ~x3 & x9 ;
  assign n209 = n208 ^ x6 ;
  assign n210 = ~n207 & ~n209 ;
  assign n211 = n210 ^ n208 ;
  assign n212 = ~x6 & n211 ;
  assign n213 = n212 ^ x3 ;
  assign n214 = n213 ^ x6 ;
  assign n215 = n96 & ~n214 ;
  assign n216 = ~x6 & n48 ;
  assign n217 = n108 & n216 ;
  assign n218 = ~x5 & n60 ;
  assign n219 = ~n128 & ~n218 ;
  assign n220 = ~n217 & n219 ;
  assign n221 = ~x2 & ~n220 ;
  assign n222 = x6 ^ x5 ;
  assign n223 = x5 ^ x2 ;
  assign n224 = n222 & n223 ;
  assign n225 = n58 & n224 ;
  assign n226 = ~x9 & n225 ;
  assign n227 = ~n221 & ~n226 ;
  assign n228 = ~n215 & n227 ;
  assign n229 = n228 ^ n199 ;
  assign n230 = n201 & n229 ;
  assign n231 = n230 ^ n199 ;
  assign n232 = ~x4 & n231 ;
  assign n233 = ~n156 & n232 ;
  assign n234 = n233 ^ n153 ;
  assign n235 = n155 & n234 ;
  assign n236 = n235 ^ n153 ;
  assign n237 = n236 ^ n39 ;
  assign n238 = n121 & ~n237 ;
  assign n239 = n238 ^ n235 ;
  assign n240 = n239 ^ n153 ;
  assign n241 = n240 ^ n120 ;
  assign n242 = ~n39 & ~n241 ;
  assign n243 = n242 ^ n39 ;
  assign y0 = n243 ;
endmodule
