module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 ;
  assign n129 = ~x7 & x8 ;
  assign n130 = ~x5 & n129 ;
  assign n131 = x4 & n130 ;
  assign n99 = ~x7 & ~x8 ;
  assign n181 = x5 & n99 ;
  assign n182 = ~n131 & ~n181 ;
  assign n183 = x1 & x2 ;
  assign n184 = ~n182 & n183 ;
  assign n159 = x5 & ~x8 ;
  assign n10 = ~x1 & ~x2 ;
  assign n185 = ~x7 & n10 ;
  assign n36 = x2 ^ x1 ;
  assign n186 = x7 & n36 ;
  assign n187 = ~n185 & ~n186 ;
  assign n188 = n159 & ~n187 ;
  assign n189 = x4 & n188 ;
  assign n190 = ~n184 & ~n189 ;
  assign n191 = ~x3 & ~n190 ;
  assign n27 = x2 & ~x3 ;
  assign n28 = ~x1 & n27 ;
  assign n132 = n28 & n131 ;
  assign n133 = x3 ^ x2 ;
  assign n138 = x4 ^ x3 ;
  assign n15 = x8 ^ x3 ;
  assign n134 = n15 ^ x5 ;
  assign n135 = n134 ^ x4 ;
  assign n136 = n135 ^ x3 ;
  assign n145 = n136 ^ x3 ;
  assign n137 = n136 ^ x5 ;
  assign n146 = n145 ^ n137 ;
  assign n147 = ~n138 & ~n146 ;
  assign n139 = x7 ^ x5 ;
  assign n140 = n139 ^ n138 ;
  assign n141 = n137 & n140 ;
  assign n153 = n147 ^ n141 ;
  assign n142 = n141 ^ n136 ;
  assign n143 = n142 ^ n138 ;
  assign n144 = n143 ^ n137 ;
  assign n148 = n147 ^ n136 ;
  assign n149 = n148 ^ n138 ;
  assign n150 = n149 ^ n137 ;
  assign n151 = n150 ^ n133 ;
  assign n152 = n144 & n151 ;
  assign n154 = n153 ^ n152 ;
  assign n155 = n133 & n154 ;
  assign n156 = x1 & n155 ;
  assign n157 = ~x2 & ~x3 ;
  assign n158 = ~x4 & x7 ;
  assign n160 = n158 & n159 ;
  assign n161 = n157 & n160 ;
  assign n162 = ~n156 & ~n161 ;
  assign n53 = x2 & x4 ;
  assign n100 = x7 & x8 ;
  assign n103 = x1 & n100 ;
  assign n163 = n53 & n103 ;
  assign n164 = x4 ^ x1 ;
  assign n165 = n164 ^ x8 ;
  assign n166 = x8 ^ x2 ;
  assign n167 = n166 ^ x2 ;
  assign n168 = x4 ^ x2 ;
  assign n169 = n168 ^ x2 ;
  assign n170 = ~n167 & n169 ;
  assign n171 = n170 ^ x2 ;
  assign n172 = n165 & ~n171 ;
  assign n173 = ~x7 & n172 ;
  assign n174 = ~n163 & ~n173 ;
  assign n175 = x3 & x5 ;
  assign n176 = ~n174 & n175 ;
  assign n177 = n162 & ~n176 ;
  assign n178 = ~n132 & n177 ;
  assign n11 = x0 & x2 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = ~x7 & n12 ;
  assign n14 = n13 ^ n11 ;
  assign n16 = x0 & ~x1 ;
  assign n17 = x4 & x8 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = n17 ^ x4 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = n21 ^ n17 ;
  assign n23 = ~n16 & n22 ;
  assign n24 = n15 & n23 ;
  assign n25 = n14 & n24 ;
  assign n54 = n15 & n53 ;
  assign n55 = ~x2 & x3 ;
  assign n56 = x1 & x4 ;
  assign n57 = n55 & ~n56 ;
  assign n58 = ~n54 & ~n57 ;
  assign n26 = ~x4 & x8 ;
  assign n29 = n26 & n28 ;
  assign n30 = x4 & ~x8 ;
  assign n31 = x1 & ~x2 ;
  assign n32 = n30 & n31 ;
  assign n33 = ~n29 & ~n32 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ n33 ;
  assign n34 = n33 ^ x3 ;
  assign n35 = n34 ^ n33 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n33 ^ n17 ;
  assign n41 = n40 ^ n33 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = n38 & n42 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = n39 & n44 ;
  assign n46 = n45 ^ n43 ;
  assign n47 = n46 ^ n33 ;
  assign n48 = n47 ^ n38 ;
  assign n49 = ~x0 & ~n48 ;
  assign n50 = n49 ^ n33 ;
  assign n59 = n58 ^ n50 ;
  assign n60 = n59 ^ n50 ;
  assign n51 = n50 ^ x0 ;
  assign n52 = n51 ^ n50 ;
  assign n61 = n60 ^ n52 ;
  assign n62 = n30 & n55 ;
  assign n63 = ~x1 & ~n62 ;
  assign n64 = n63 ^ n50 ;
  assign n65 = n64 ^ n50 ;
  assign n66 = n65 ^ n60 ;
  assign n67 = ~n60 & n66 ;
  assign n68 = n67 ^ n60 ;
  assign n69 = n61 & ~n68 ;
  assign n70 = n69 ^ n67 ;
  assign n71 = n70 ^ n50 ;
  assign n72 = n71 ^ n60 ;
  assign n73 = x7 & n72 ;
  assign n74 = n73 ^ n50 ;
  assign n75 = n74 ^ x5 ;
  assign n76 = n75 ^ n74 ;
  assign n77 = x4 ^ x0 ;
  assign n78 = n77 ^ x7 ;
  assign n79 = x8 ^ x1 ;
  assign n87 = n79 ^ x8 ;
  assign n88 = n87 ^ x8 ;
  assign n89 = n87 & n88 ;
  assign n81 = n79 ^ x7 ;
  assign n80 = n79 ^ x4 ;
  assign n82 = n81 ^ n80 ;
  assign n83 = n81 ^ n79 ;
  assign n84 = n83 ^ x8 ;
  assign n85 = n82 & ~n84 ;
  assign n92 = n89 ^ n85 ;
  assign n86 = n85 ^ n78 ;
  assign n90 = n89 ^ n87 ;
  assign n91 = n86 & n90 ;
  assign n93 = n92 ^ n91 ;
  assign n94 = n78 & n93 ;
  assign n95 = n94 ^ n85 ;
  assign n96 = n95 ^ n89 ;
  assign n97 = n96 ^ n91 ;
  assign n98 = n55 & n97 ;
  assign n109 = x0 & ~n17 ;
  assign n101 = ~x1 & ~n100 ;
  assign n102 = ~n99 & n101 ;
  assign n104 = ~n102 & ~n103 ;
  assign n105 = n11 & ~n104 ;
  assign n106 = ~x4 & n105 ;
  assign n110 = n109 ^ n106 ;
  assign n111 = n110 ^ n106 ;
  assign n107 = n106 ^ n102 ;
  assign n108 = n107 ^ n106 ;
  assign n112 = n111 ^ n108 ;
  assign n113 = n106 ^ x2 ;
  assign n114 = n113 ^ n106 ;
  assign n115 = n114 ^ n111 ;
  assign n116 = n111 & ~n115 ;
  assign n117 = n116 ^ n111 ;
  assign n118 = n112 & n117 ;
  assign n119 = n118 ^ n116 ;
  assign n120 = n119 ^ n106 ;
  assign n121 = n120 ^ n111 ;
  assign n122 = ~x3 & n121 ;
  assign n123 = n122 ^ n106 ;
  assign n124 = ~n98 & ~n123 ;
  assign n125 = n124 ^ n74 ;
  assign n126 = n76 & n125 ;
  assign n127 = n126 ^ n74 ;
  assign n128 = ~n25 & n127 ;
  assign n179 = n178 ^ n128 ;
  assign n180 = n179 ^ n178 ;
  assign n192 = n191 ^ n180 ;
  assign n193 = n192 ^ n179 ;
  assign n194 = n179 ^ x0 ;
  assign n195 = n194 ^ n179 ;
  assign n196 = ~n193 & ~n195 ;
  assign n197 = n196 ^ n179 ;
  assign n198 = ~x6 & n197 ;
  assign n199 = n198 ^ n128 ;
  assign y0 = ~n199 ;
endmodule
