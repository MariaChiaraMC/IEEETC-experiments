module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 ;
  assign n15 = ~x3 & x4 ;
  assign n16 = n15 ^ x2 ;
  assign n17 = n15 ^ x6 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = ~x1 & ~x7 ;
  assign n21 = x0 & ~n20 ;
  assign n22 = n21 ^ x3 ;
  assign n23 = ~n15 & ~n22 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n19 & ~n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n26 ^ n21 ;
  assign n28 = n27 ^ n15 ;
  assign n29 = ~n16 & n28 ;
  assign n30 = n29 ^ x2 ;
  assign n31 = x5 & ~n30 ;
  assign n32 = x13 & n31 ;
  assign n33 = x8 ^ x0 ;
  assign n34 = n33 ^ x8 ;
  assign n35 = x10 ^ x8 ;
  assign n36 = ~n34 & ~n35 ;
  assign n37 = n36 ^ x8 ;
  assign n38 = ~n20 & ~n37 ;
  assign n39 = n38 ^ x0 ;
  assign n40 = x5 & x6 ;
  assign n41 = ~x2 & ~x12 ;
  assign n42 = n40 & n41 ;
  assign n43 = n15 & n42 ;
  assign n44 = ~x11 & ~n43 ;
  assign n45 = n44 ^ n21 ;
  assign n46 = n45 ^ n39 ;
  assign n47 = ~x6 & n15 ;
  assign n48 = x5 & n47 ;
  assign n49 = x2 & n48 ;
  assign n50 = n49 ^ x9 ;
  assign n51 = n21 & ~n50 ;
  assign n52 = n51 ^ x9 ;
  assign n53 = ~n46 & n52 ;
  assign n54 = n53 ^ n51 ;
  assign n55 = n54 ^ x9 ;
  assign n56 = n55 ^ n21 ;
  assign n57 = n39 & n56 ;
  assign n58 = ~n32 & ~n57 ;
  assign y0 = ~n58 ;
endmodule
