// Benchmark "./newtpla1.pla" written by ABC on Thu Apr 23 10:59:58 2020

module \./newtpla1.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9,
    z0  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
  output z0;
  assign z0 = x0 | x2;
endmodule


