module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 ;
  assign n11 = x3 & ~x9 ;
  assign n12 = x2 & ~x5 ;
  assign n13 = ~x6 & n12 ;
  assign n14 = ~x7 & n13 ;
  assign n15 = ~x5 & x7 ;
  assign n16 = x5 & ~x7 ;
  assign n17 = ~n15 & ~n16 ;
  assign n18 = ~x1 & ~x2 ;
  assign n19 = x6 & n18 ;
  assign n20 = ~n17 & n19 ;
  assign n21 = ~n14 & ~n20 ;
  assign n22 = n11 & ~n21 ;
  assign n23 = ~x4 & n22 ;
  assign n24 = ~x3 & ~x6 ;
  assign n25 = ~x4 & x9 ;
  assign n26 = n24 & ~n25 ;
  assign n27 = ~x7 & ~x9 ;
  assign n28 = n18 & ~n27 ;
  assign n29 = n26 & n28 ;
  assign n30 = n17 & n29 ;
  assign n31 = ~x5 & ~x6 ;
  assign n32 = x2 & ~x4 ;
  assign n33 = ~x9 & n32 ;
  assign n34 = ~x7 & x9 ;
  assign n35 = ~x2 & x4 ;
  assign n36 = n34 & n35 ;
  assign n37 = ~n33 & ~n36 ;
  assign n38 = x1 & ~n37 ;
  assign n39 = n18 & n34 ;
  assign n40 = ~x4 & n39 ;
  assign n41 = ~n38 & ~n40 ;
  assign n42 = n31 & ~n41 ;
  assign n43 = x7 & x9 ;
  assign n44 = x1 & ~x5 ;
  assign n45 = n43 & n44 ;
  assign n46 = x7 & ~x9 ;
  assign n47 = n46 ^ x9 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = n46 ^ n16 ;
  assign n50 = n49 ^ n46 ;
  assign n51 = n48 & n50 ;
  assign n52 = n51 ^ n46 ;
  assign n53 = ~x4 & n52 ;
  assign n54 = n53 ^ n46 ;
  assign n55 = ~x1 & n54 ;
  assign n56 = ~n45 & ~n55 ;
  assign n57 = x2 & x6 ;
  assign n58 = ~n56 & n57 ;
  assign n59 = x1 & x6 ;
  assign n60 = x7 ^ x4 ;
  assign n61 = n60 ^ x9 ;
  assign n62 = n61 ^ x2 ;
  assign n63 = x9 ^ x7 ;
  assign n64 = x7 ^ x5 ;
  assign n65 = n64 ^ x7 ;
  assign n66 = n63 & n65 ;
  assign n67 = n66 ^ x7 ;
  assign n68 = n67 ^ n61 ;
  assign n69 = ~n62 & ~n68 ;
  assign n70 = n69 ^ n66 ;
  assign n71 = n70 ^ x7 ;
  assign n72 = n71 ^ x2 ;
  assign n73 = n61 & n72 ;
  assign n74 = n73 ^ n61 ;
  assign n75 = n59 & n74 ;
  assign n76 = ~n58 & ~n75 ;
  assign n77 = ~n42 & n76 ;
  assign n78 = x3 & ~n77 ;
  assign n79 = ~x6 & n43 ;
  assign n80 = ~x3 & ~x5 ;
  assign n81 = n79 & n80 ;
  assign n82 = n81 ^ x5 ;
  assign n83 = n82 ^ n81 ;
  assign n84 = x6 & n27 ;
  assign n85 = n84 ^ n81 ;
  assign n86 = n85 ^ n81 ;
  assign n87 = n83 & n86 ;
  assign n88 = n87 ^ n81 ;
  assign n89 = x1 & n88 ;
  assign n90 = n89 ^ n81 ;
  assign n91 = n32 & n90 ;
  assign n92 = n80 & n84 ;
  assign n93 = x5 & x6 ;
  assign n94 = n34 & n93 ;
  assign n95 = x5 & x7 ;
  assign n96 = ~x6 & ~x9 ;
  assign n97 = ~x3 & n96 ;
  assign n98 = ~n95 & n97 ;
  assign n99 = ~n94 & ~n98 ;
  assign n100 = x2 & ~n99 ;
  assign n101 = ~n92 & ~n100 ;
  assign n102 = x1 & x4 ;
  assign n103 = ~n101 & n102 ;
  assign n104 = ~n91 & ~n103 ;
  assign n105 = ~n78 & n104 ;
  assign n106 = ~n30 & n105 ;
  assign n107 = n106 ^ x8 ;
  assign n108 = n107 ^ n106 ;
  assign n109 = ~x2 & n59 ;
  assign n111 = x5 & x9 ;
  assign n110 = ~x4 & ~x5 ;
  assign n112 = n111 ^ n110 ;
  assign n113 = ~x3 & n112 ;
  assign n114 = n113 ^ n111 ;
  assign n115 = n109 & n114 ;
  assign n116 = ~x2 & ~x9 ;
  assign n117 = x5 & ~x6 ;
  assign n118 = ~x4 & n117 ;
  assign n119 = ~x1 & ~x3 ;
  assign n120 = n118 & n119 ;
  assign n121 = n116 & n120 ;
  assign n122 = ~x4 & ~x6 ;
  assign n123 = ~n11 & ~n122 ;
  assign n124 = n123 ^ n12 ;
  assign n125 = ~x6 & n11 ;
  assign n126 = n125 ^ x1 ;
  assign n127 = n126 ^ n125 ;
  assign n128 = n125 ^ n96 ;
  assign n129 = ~n127 & ~n128 ;
  assign n130 = n129 ^ n125 ;
  assign n131 = n130 ^ n123 ;
  assign n132 = ~n124 & ~n131 ;
  assign n133 = n132 ^ n129 ;
  assign n134 = n133 ^ n125 ;
  assign n135 = n134 ^ n12 ;
  assign n136 = ~n123 & n135 ;
  assign n137 = n136 ^ n123 ;
  assign n138 = ~n121 & n137 ;
  assign n139 = ~n115 & n138 ;
  assign n140 = ~x7 & ~n139 ;
  assign n141 = x3 & ~n43 ;
  assign n142 = ~x1 & ~n31 ;
  assign n143 = ~n111 & ~n142 ;
  assign n144 = ~n141 & ~n143 ;
  assign n145 = ~x2 & x7 ;
  assign n146 = x3 & x7 ;
  assign n147 = ~n145 & ~n146 ;
  assign n148 = ~n93 & ~n147 ;
  assign n149 = ~x1 & ~n46 ;
  assign n150 = ~n148 & n149 ;
  assign n151 = n144 & ~n150 ;
  assign n152 = x2 ^ x1 ;
  assign n153 = n152 ^ x3 ;
  assign n154 = x6 ^ x1 ;
  assign n155 = n154 ^ x6 ;
  assign n156 = n111 ^ x6 ;
  assign n157 = ~n155 & n156 ;
  assign n158 = n157 ^ x6 ;
  assign n159 = n158 ^ n152 ;
  assign n160 = n153 & ~n159 ;
  assign n161 = n160 ^ n157 ;
  assign n162 = n161 ^ x6 ;
  assign n163 = n162 ^ x3 ;
  assign n164 = ~n152 & ~n163 ;
  assign n165 = n164 ^ n152 ;
  assign n166 = n165 ^ x2 ;
  assign n167 = n151 & ~n166 ;
  assign n168 = n167 ^ x4 ;
  assign n169 = n168 ^ n167 ;
  assign n170 = n169 ^ n140 ;
  assign n171 = x7 ^ x2 ;
  assign n172 = n171 ^ n43 ;
  assign n173 = x7 ^ x3 ;
  assign n174 = n43 ^ x3 ;
  assign n175 = n174 ^ x3 ;
  assign n176 = n173 & n175 ;
  assign n177 = n176 ^ x3 ;
  assign n178 = ~n172 & n177 ;
  assign n179 = n178 ^ n43 ;
  assign n180 = n31 & n179 ;
  assign n186 = x3 & ~n116 ;
  assign n181 = ~x2 & x5 ;
  assign n182 = n34 & n181 ;
  assign n187 = n186 ^ n182 ;
  assign n188 = n187 ^ n182 ;
  assign n183 = ~n43 & ~n146 ;
  assign n184 = n183 ^ n182 ;
  assign n185 = n184 ^ n182 ;
  assign n189 = n188 ^ n185 ;
  assign n190 = n182 ^ x5 ;
  assign n191 = n190 ^ n182 ;
  assign n192 = n191 ^ n188 ;
  assign n193 = ~n188 & ~n192 ;
  assign n194 = n193 ^ n188 ;
  assign n195 = n189 & ~n194 ;
  assign n196 = n195 ^ n193 ;
  assign n197 = n196 ^ n182 ;
  assign n198 = n197 ^ n188 ;
  assign n199 = x6 & ~n198 ;
  assign n200 = n199 ^ n182 ;
  assign n201 = ~n180 & ~n200 ;
  assign n202 = ~x1 & n201 ;
  assign n203 = x5 & n79 ;
  assign n204 = ~x7 & n116 ;
  assign n205 = ~n93 & n204 ;
  assign n206 = ~n203 & ~n205 ;
  assign n207 = x5 ^ x3 ;
  assign n208 = ~n206 & ~n207 ;
  assign n209 = x1 & ~n208 ;
  assign n210 = n80 ^ x9 ;
  assign n211 = n210 ^ n80 ;
  assign n212 = x3 & x5 ;
  assign n213 = n212 ^ n80 ;
  assign n214 = ~n211 & n213 ;
  assign n215 = n214 ^ n80 ;
  assign n216 = n63 & n215 ;
  assign n217 = n216 ^ x2 ;
  assign n218 = n217 ^ n216 ;
  assign n219 = ~n95 & ~n141 ;
  assign n220 = ~x9 & ~n15 ;
  assign n221 = ~n219 & ~n220 ;
  assign n222 = n221 ^ n216 ;
  assign n223 = ~n218 & n222 ;
  assign n224 = n223 ^ n216 ;
  assign n225 = x6 & n224 ;
  assign n226 = n209 & ~n225 ;
  assign n227 = n226 ^ n202 ;
  assign n228 = ~n202 & n227 ;
  assign n229 = n228 ^ n167 ;
  assign n230 = n229 ^ n202 ;
  assign n231 = ~n170 & ~n230 ;
  assign n232 = n231 ^ n228 ;
  assign n233 = n232 ^ n202 ;
  assign n234 = ~n140 & ~n233 ;
  assign n235 = n234 ^ n140 ;
  assign n236 = n235 ^ n106 ;
  assign n237 = n108 & ~n236 ;
  assign n238 = n237 ^ n106 ;
  assign n239 = ~n23 & n238 ;
  assign n242 = n239 ^ x7 ;
  assign n243 = n242 ^ n239 ;
  assign n240 = n239 ^ n32 ;
  assign n241 = n240 ^ n239 ;
  assign n244 = n243 ^ n241 ;
  assign n245 = x1 & x5 ;
  assign n246 = x8 & n96 ;
  assign n247 = n245 & n246 ;
  assign n248 = n247 ^ n239 ;
  assign n249 = n248 ^ n239 ;
  assign n250 = n249 ^ n243 ;
  assign n251 = n243 & n250 ;
  assign n252 = n251 ^ n243 ;
  assign n253 = n244 & n252 ;
  assign n254 = n253 ^ n251 ;
  assign n255 = n254 ^ n239 ;
  assign n256 = n255 ^ n243 ;
  assign n257 = ~x0 & ~n256 ;
  assign n258 = n257 ^ n239 ;
  assign n366 = ~x6 & x8 ;
  assign n367 = x6 & ~x8 ;
  assign n368 = ~n366 & ~n367 ;
  assign n369 = ~x1 & x4 ;
  assign n370 = n34 & n369 ;
  assign n371 = ~n368 & n370 ;
  assign n372 = ~n13 & ~n181 ;
  assign n373 = n371 & ~n372 ;
  assign n303 = ~x5 & x6 ;
  assign n374 = ~n95 & ~n303 ;
  assign n375 = ~x1 & n374 ;
  assign n289 = x5 & ~x8 ;
  assign n376 = ~n289 & ~n366 ;
  assign n377 = x9 & n376 ;
  assign n378 = n375 & n377 ;
  assign n290 = x2 & x4 ;
  assign n264 = x6 & x8 ;
  assign n379 = n45 & n264 ;
  assign n380 = n46 & n117 ;
  assign n381 = x1 & n380 ;
  assign n382 = ~n247 & ~n381 ;
  assign n383 = ~n379 & n382 ;
  assign n384 = n290 & n383 ;
  assign n385 = ~n378 & n384 ;
  assign n386 = n43 & n366 ;
  assign n387 = ~x5 & n386 ;
  assign n388 = ~x2 & ~n387 ;
  assign n389 = n43 & n367 ;
  assign n390 = n27 & n31 ;
  assign n391 = ~n389 & ~n390 ;
  assign n392 = n391 ^ x1 ;
  assign n393 = n392 ^ n391 ;
  assign n394 = n393 ^ n388 ;
  assign n395 = n27 & n289 ;
  assign n396 = n395 ^ x6 ;
  assign n397 = ~x6 & ~n396 ;
  assign n398 = n397 ^ n391 ;
  assign n399 = n398 ^ x6 ;
  assign n400 = ~n394 & n399 ;
  assign n401 = n400 ^ n397 ;
  assign n402 = n401 ^ x6 ;
  assign n403 = n388 & ~n402 ;
  assign n404 = n403 ^ n388 ;
  assign n405 = ~n385 & ~n404 ;
  assign n406 = n44 & n46 ;
  assign n407 = ~n368 & n406 ;
  assign n408 = ~n405 & ~n407 ;
  assign n266 = ~x2 & ~x4 ;
  assign n409 = n27 & n264 ;
  assign n410 = ~n389 & ~n409 ;
  assign n411 = n245 & ~n410 ;
  assign n412 = n34 & n117 ;
  assign n413 = ~n390 & ~n412 ;
  assign n414 = x1 & ~x8 ;
  assign n415 = ~n413 & n414 ;
  assign n416 = x5 & n386 ;
  assign n417 = ~x4 & ~n416 ;
  assign n418 = ~n415 & n417 ;
  assign n419 = ~n411 & n418 ;
  assign n420 = ~n266 & ~n419 ;
  assign n421 = ~n408 & n420 ;
  assign n422 = x8 ^ x6 ;
  assign n423 = x9 ^ x8 ;
  assign n424 = ~n422 & ~n423 ;
  assign n425 = n266 & n424 ;
  assign n360 = x9 & n264 ;
  assign n426 = x7 & ~n360 ;
  assign n427 = n426 ^ n95 ;
  assign n428 = n427 ^ n95 ;
  assign n429 = n95 ^ x5 ;
  assign n430 = n429 ^ n95 ;
  assign n431 = ~n428 & ~n430 ;
  assign n432 = n431 ^ n95 ;
  assign n433 = ~x1 & n432 ;
  assign n434 = n433 ^ n95 ;
  assign n435 = n425 & n434 ;
  assign n436 = n39 & n303 ;
  assign n437 = x8 & n436 ;
  assign n438 = ~n435 & ~n437 ;
  assign n439 = ~n421 & n438 ;
  assign n440 = ~x0 & ~n439 ;
  assign n441 = ~n373 & ~n440 ;
  assign n259 = ~x1 & ~x5 ;
  assign n260 = x7 & ~x8 ;
  assign n261 = n259 & n260 ;
  assign n262 = n35 & n261 ;
  assign n263 = x5 & n46 ;
  assign n265 = n264 ^ n263 ;
  assign n267 = n266 ^ x1 ;
  assign n268 = n267 ^ n266 ;
  assign n269 = n266 ^ x2 ;
  assign n270 = ~n268 & n269 ;
  assign n271 = n270 ^ n266 ;
  assign n272 = n271 ^ n263 ;
  assign n273 = n265 & n272 ;
  assign n274 = n273 ^ n270 ;
  assign n275 = n274 ^ n266 ;
  assign n276 = n275 ^ n264 ;
  assign n277 = n263 & n276 ;
  assign n278 = n277 ^ n263 ;
  assign n279 = ~n262 & ~n278 ;
  assign n283 = ~x2 & ~x6 ;
  assign n280 = x6 ^ x5 ;
  assign n281 = x5 ^ x4 ;
  assign n282 = n280 & n281 ;
  assign n284 = n283 ^ n282 ;
  assign n285 = ~x8 & n284 ;
  assign n286 = n285 ^ x1 ;
  assign n287 = n286 ^ n285 ;
  assign n288 = n287 ^ n27 ;
  assign n291 = n289 & n290 ;
  assign n292 = n264 & n266 ;
  assign n293 = n292 ^ n291 ;
  assign n294 = ~n291 & n293 ;
  assign n295 = n294 ^ n285 ;
  assign n296 = n295 ^ n291 ;
  assign n297 = ~n288 & n296 ;
  assign n298 = n297 ^ n294 ;
  assign n299 = n298 ^ n291 ;
  assign n300 = n27 & ~n299 ;
  assign n301 = n300 ^ n27 ;
  assign n302 = n279 & ~n301 ;
  assign n304 = x4 & n303 ;
  assign n305 = n260 & n304 ;
  assign n309 = x4 & x7 ;
  assign n310 = n181 & ~n309 ;
  assign n306 = x7 ^ x6 ;
  assign n307 = ~x4 & n306 ;
  assign n308 = n307 ^ x6 ;
  assign n311 = n310 ^ n308 ;
  assign n312 = n311 ^ n310 ;
  assign n313 = ~x6 & ~x7 ;
  assign n314 = x2 & ~n313 ;
  assign n315 = ~n16 & n314 ;
  assign n316 = n315 ^ n310 ;
  assign n317 = ~n312 & n316 ;
  assign n318 = n317 ^ n310 ;
  assign n319 = x8 & n318 ;
  assign n320 = ~n305 & ~n319 ;
  assign n321 = n320 ^ x1 ;
  assign n322 = n321 ^ n320 ;
  assign n323 = n117 ^ x4 ;
  assign n324 = ~n303 & ~n323 ;
  assign n325 = x7 & n324 ;
  assign n326 = ~x2 & ~n325 ;
  assign n332 = n93 & n309 ;
  assign n327 = x4 & x6 ;
  assign n328 = ~n118 & ~n327 ;
  assign n329 = ~x7 & ~n328 ;
  assign n333 = n332 ^ n329 ;
  assign n334 = n333 ^ n329 ;
  assign n330 = n329 ^ x2 ;
  assign n331 = n330 ^ n329 ;
  assign n335 = n334 ^ n331 ;
  assign n336 = n110 & n313 ;
  assign n337 = n336 ^ n329 ;
  assign n338 = n337 ^ n329 ;
  assign n339 = n338 ^ n334 ;
  assign n340 = ~n334 & n339 ;
  assign n341 = n340 ^ n334 ;
  assign n342 = ~n335 & ~n341 ;
  assign n343 = n342 ^ n340 ;
  assign n344 = n343 ^ n329 ;
  assign n345 = n344 ^ n334 ;
  assign n346 = ~x8 & n345 ;
  assign n347 = n346 ^ n329 ;
  assign n348 = ~n326 & n347 ;
  assign n349 = n348 ^ n320 ;
  assign n350 = n322 & ~n349 ;
  assign n351 = n350 ^ n320 ;
  assign n352 = x9 & ~n351 ;
  assign n353 = n302 & ~n352 ;
  assign n354 = ~x0 & ~n353 ;
  assign n355 = x6 & n261 ;
  assign n356 = n35 ^ n32 ;
  assign n357 = x9 & n356 ;
  assign n358 = n357 ^ n32 ;
  assign n359 = n355 & n358 ;
  assign n361 = ~x7 & n245 ;
  assign n362 = n360 & n361 ;
  assign n363 = n290 & n362 ;
  assign n364 = ~n359 & ~n363 ;
  assign n365 = ~n354 & n364 ;
  assign n442 = n441 ^ n365 ;
  assign n443 = x3 & n442 ;
  assign n444 = n443 ^ n441 ;
  assign n445 = n258 & n444 ;
  assign y0 = ~n445 ;
endmodule
