// Benchmark "./exp.pla" written by ABC on Thu Apr 23 10:59:51 2020

module \./exp.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z17  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z17;
  wire new_n10_, new_n11_, new_n12_, new_n13_, new_n14_, new_n15_, new_n16_,
    new_n17_, new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_,
    new_n24_, new_n25_, new_n26_, new_n27_, new_n28_;
  assign new_n10_ = x1 & ~x5;
  assign new_n11_ = x2 & x6;
  assign new_n12_ = x0 & new_n11_;
  assign new_n13_ = ~x2 & ~x6;
  assign new_n14_ = ~new_n12_ & ~new_n13_;
  assign new_n15_ = new_n10_ & ~new_n14_;
  assign new_n16_ = ~x1 & x5;
  assign new_n17_ = x6 & ~new_n16_;
  assign new_n18_ = ~x0 & ~new_n17_;
  assign new_n19_ = ~new_n15_ & ~new_n18_;
  assign new_n20_ = ~x6 & ~new_n10_;
  assign new_n21_ = ~x3 & ~new_n20_;
  assign new_n22_ = ~new_n19_ & new_n21_;
  assign new_n23_ = x0 & x3;
  assign new_n24_ = x5 & ~new_n13_;
  assign new_n25_ = ~x5 & ~new_n11_;
  assign new_n26_ = ~new_n24_ & ~new_n25_;
  assign new_n27_ = new_n23_ & new_n26_;
  assign new_n28_ = ~x1 & new_n27_;
  assign z17 = new_n22_ | new_n28_;
endmodule


