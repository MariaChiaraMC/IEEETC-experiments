module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 ;
  assign n12 = x2 & ~x8 ;
  assign n27 = ~x4 & ~x5 ;
  assign n65 = ~x3 & ~x6 ;
  assign n66 = n27 & n65 ;
  assign n67 = n12 & ~n66 ;
  assign n68 = x7 & n67 ;
  assign n69 = ~x7 & x8 ;
  assign n10 = x5 & x6 ;
  assign n70 = x4 & n10 ;
  assign n71 = ~x2 & x8 ;
  assign n72 = ~x3 & n71 ;
  assign n73 = ~n70 & n72 ;
  assign n74 = ~n69 & ~n73 ;
  assign n75 = ~n68 & n74 ;
  assign n49 = x7 & ~x8 ;
  assign n50 = ~x0 & ~n49 ;
  assign n15 = x2 ^ x0 ;
  assign n16 = n15 ^ x7 ;
  assign n17 = n16 ^ x7 ;
  assign n18 = n17 ^ x0 ;
  assign n19 = n18 ^ x0 ;
  assign n20 = x8 ^ x0 ;
  assign n21 = n20 ^ x7 ;
  assign n22 = n21 ^ x0 ;
  assign n23 = n19 & ~n22 ;
  assign n24 = n23 ^ x7 ;
  assign n25 = n24 ^ x0 ;
  assign n26 = n25 ^ n18 ;
  assign n28 = n27 ^ x7 ;
  assign n29 = n28 ^ x0 ;
  assign n30 = n27 & n29 ;
  assign n31 = n27 ^ n21 ;
  assign n32 = n31 ^ x0 ;
  assign n33 = n32 ^ n18 ;
  assign n34 = x6 & ~n33 ;
  assign n35 = n34 ^ x6 ;
  assign n36 = n35 ^ n27 ;
  assign n37 = n36 ^ x0 ;
  assign n38 = n37 ^ n18 ;
  assign n39 = n30 & n38 ;
  assign n40 = n39 ^ x0 ;
  assign n41 = n26 & n40 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = n42 ^ x7 ;
  assign n44 = n43 ^ x0 ;
  assign n45 = n44 ^ x7 ;
  assign n46 = n45 ^ x7 ;
  assign n47 = n46 ^ x3 ;
  assign n11 = ~x4 & ~n10 ;
  assign n13 = ~n11 & n12 ;
  assign n14 = n13 ^ x3 ;
  assign n48 = n47 ^ n14 ;
  assign n51 = n50 ^ n48 ;
  assign n52 = n51 ^ n48 ;
  assign n53 = n48 ^ n47 ;
  assign n54 = n53 ^ x3 ;
  assign n55 = n52 & ~n54 ;
  assign n56 = n55 ^ n47 ;
  assign n57 = x7 & n47 ;
  assign n58 = n57 ^ x3 ;
  assign n59 = n56 & ~n58 ;
  assign n60 = n59 ^ n57 ;
  assign n61 = ~x3 & n60 ;
  assign n62 = n61 ^ n55 ;
  assign n63 = n62 ^ n46 ;
  assign n64 = n63 ^ n47 ;
  assign n76 = n75 ^ n64 ;
  assign n77 = n76 ^ n64 ;
  assign n78 = n64 ^ x0 ;
  assign n79 = n78 ^ n64 ;
  assign n80 = ~n77 & ~n79 ;
  assign n81 = n80 ^ n64 ;
  assign n82 = x1 & ~n81 ;
  assign n83 = n82 ^ n64 ;
  assign y0 = ~n83 ;
endmodule
