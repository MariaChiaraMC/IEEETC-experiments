// Benchmark "./pla/x2dn.pla_dbb_orig_11NonExact" written by ABC on Fri Nov 20 10:30:31 2020

module \./pla/x2dn.pla_dbb_orig_11NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = 1'b1;
endmodule


