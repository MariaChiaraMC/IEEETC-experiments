module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 ;
  output y0 ;
  wire n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 ;
  assign n19 = x6 & x16 ;
  assign n20 = ~x6 & ~x16 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = x4 & ~x8 ;
  assign n23 = ~x7 & x15 ;
  assign n24 = x5 & n23 ;
  assign n25 = n22 & n24 ;
  assign n26 = ~n21 & n25 ;
  assign n27 = x15 ^ x6 ;
  assign n28 = x15 ^ x13 ;
  assign n29 = n28 ^ x13 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = ~x7 & x16 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = n22 & ~n32 ;
  assign n34 = n33 ^ x13 ;
  assign n35 = ~n30 & n34 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = ~n27 & n36 ;
  assign n38 = n37 ^ n33 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = ~x5 & n39 ;
  assign n41 = ~x15 & ~x16 ;
  assign n42 = x5 & ~x15 ;
  assign n43 = x5 & ~x16 ;
  assign n44 = ~n42 & ~n43 ;
  assign n45 = ~n41 & ~n44 ;
  assign n46 = ~x7 & ~n41 ;
  assign n47 = ~n19 & ~n46 ;
  assign n48 = ~n45 & n47 ;
  assign n49 = x13 & ~n48 ;
  assign n50 = ~n40 & ~n49 ;
  assign n51 = ~n26 & n50 ;
  assign n52 = ~x14 & ~n51 ;
  assign n69 = ~n23 & n45 ;
  assign n70 = x5 & ~x6 ;
  assign n71 = x6 & x7 ;
  assign n72 = x5 & x16 ;
  assign n73 = x15 & ~n72 ;
  assign n74 = ~n71 & n73 ;
  assign n75 = ~n70 & n74 ;
  assign n76 = ~n69 & ~n75 ;
  assign n77 = ~x2 & ~x9 ;
  assign n78 = n77 ^ x16 ;
  assign n79 = n77 ^ x15 ;
  assign n80 = n79 ^ x15 ;
  assign n81 = ~x6 & ~x7 ;
  assign n82 = ~n71 & ~n81 ;
  assign n83 = n82 ^ x15 ;
  assign n84 = n80 & n83 ;
  assign n85 = n84 ^ x15 ;
  assign n86 = ~n78 & n85 ;
  assign n87 = n86 ^ x16 ;
  assign n88 = n76 & ~n87 ;
  assign n53 = ~x10 & ~x11 ;
  assign n54 = x1 & ~x12 ;
  assign n55 = ~n53 & n54 ;
  assign n56 = n41 & ~n55 ;
  assign n57 = x4 & x7 ;
  assign n58 = ~n41 & ~n57 ;
  assign n59 = x16 ^ x6 ;
  assign n60 = x15 ^ x5 ;
  assign n61 = n60 ^ x16 ;
  assign n62 = n59 & n61 ;
  assign n63 = n62 ^ n58 ;
  assign n64 = n41 & ~n63 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = ~n58 & n65 ;
  assign n67 = ~x3 & ~n66 ;
  assign n68 = ~n56 & ~n67 ;
  assign n89 = n88 ^ n68 ;
  assign n90 = ~x14 & ~n89 ;
  assign n91 = n90 ^ n88 ;
  assign n92 = ~x13 & ~n91 ;
  assign n93 = ~n52 & ~n92 ;
  assign n94 = ~x17 & ~n93 ;
  assign n95 = ~x8 & ~x13 ;
  assign n96 = ~x5 & n21 ;
  assign n97 = ~x7 & ~n96 ;
  assign n98 = ~n95 & ~n97 ;
  assign n101 = ~n21 & ~n42 ;
  assign n99 = ~x17 & ~n19 ;
  assign n100 = ~x15 & ~n99 ;
  assign n102 = n101 ^ n100 ;
  assign n103 = ~x5 & n102 ;
  assign n104 = n102 ^ n100 ;
  assign n105 = ~n20 & n95 ;
  assign n106 = ~x7 & ~n105 ;
  assign n107 = n106 ^ n103 ;
  assign n108 = n104 & n107 ;
  assign n109 = n108 ^ n106 ;
  assign n110 = n103 & n109 ;
  assign n111 = n110 ^ n101 ;
  assign n112 = ~n98 & n111 ;
  assign n113 = x14 ^ x13 ;
  assign n114 = n113 ^ x14 ;
  assign n115 = ~x8 & ~x17 ;
  assign n116 = x14 & n77 ;
  assign n117 = ~n115 & n116 ;
  assign n118 = n117 ^ x14 ;
  assign n119 = ~n114 & ~n118 ;
  assign n120 = n119 ^ x14 ;
  assign n121 = n112 & ~n120 ;
  assign n122 = ~n94 & ~n121 ;
  assign n123 = ~x0 & ~n122 ;
  assign y0 = n123 ;
endmodule
