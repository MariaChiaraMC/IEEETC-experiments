module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 ;
  assign n20 = x16 & x17 ;
  assign n21 = ~x10 & x18 ;
  assign n22 = n20 & n21 ;
  assign n23 = x2 & x10 ;
  assign n29 = x11 & x13 ;
  assign n30 = x14 & ~n29 ;
  assign n31 = ~x15 & ~n30 ;
  assign n32 = ~x3 & x13 ;
  assign n33 = x12 & ~n32 ;
  assign n34 = ~n31 & n33 ;
  assign n35 = ~x14 & x15 ;
  assign n36 = ~x12 & n35 ;
  assign n37 = x11 & n32 ;
  assign n38 = ~n36 & ~n37 ;
  assign n39 = x4 & n38 ;
  assign n40 = ~n34 & n39 ;
  assign n41 = x6 ^ x3 ;
  assign n42 = n41 ^ x6 ;
  assign n43 = x7 ^ x6 ;
  assign n44 = n42 & n43 ;
  assign n45 = n44 ^ x6 ;
  assign n46 = ~n35 & n45 ;
  assign n47 = ~n40 & ~n46 ;
  assign n24 = x0 & x3 ;
  assign n25 = x9 & n24 ;
  assign n26 = x8 & n25 ;
  assign n48 = n47 ^ n26 ;
  assign n49 = n48 ^ n26 ;
  assign n27 = n26 ^ x5 ;
  assign n28 = n27 ^ n26 ;
  assign n50 = n49 ^ n28 ;
  assign n51 = n26 ^ x0 ;
  assign n52 = n51 ^ n26 ;
  assign n53 = n52 ^ n49 ;
  assign n54 = ~n49 & n53 ;
  assign n55 = n54 ^ n49 ;
  assign n56 = ~n50 & ~n55 ;
  assign n57 = n56 ^ n54 ;
  assign n58 = n57 ^ n26 ;
  assign n59 = n58 ^ n49 ;
  assign n60 = x1 & ~n59 ;
  assign n61 = n60 ^ n26 ;
  assign n62 = n23 & n61 ;
  assign n63 = ~n22 & ~n62 ;
  assign y0 = ~n63 ;
endmodule
