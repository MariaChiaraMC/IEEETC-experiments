module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n13 = x5 & x9 ;
  assign n14 = ~x7 & ~n13 ;
  assign n15 = ~x8 & ~n14 ;
  assign n16 = x6 & ~n15 ;
  assign n17 = ~x5 & ~x9 ;
  assign n18 = ~x11 & ~n17 ;
  assign n19 = x10 & ~n18 ;
  assign n20 = ~n16 & n19 ;
  assign n21 = x4 & ~n20 ;
  assign n22 = ~x1 & ~x3 ;
  assign n23 = ~x0 & n22 ;
  assign n24 = ~n21 & n23 ;
  assign n25 = x4 & ~x7 ;
  assign n26 = x0 & n25 ;
  assign n27 = ~x8 & n26 ;
  assign n28 = ~n24 & ~n27 ;
  assign y0 = ~n28 ;
endmodule
