module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 ;
  assign n16 = ~x1 & ~x8 ;
  assign n17 = ~x3 & ~n16 ;
  assign n18 = x5 & ~n17 ;
  assign n19 = ~x2 & n18 ;
  assign n21 = ~x9 & ~x14 ;
  assign n20 = x8 ^ x4 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n21 ^ x3 ;
  assign n24 = x8 ^ x3 ;
  assign n25 = n23 & n24 ;
  assign n26 = n25 ^ x3 ;
  assign n27 = ~n22 & n26 ;
  assign n28 = n27 ^ x4 ;
  assign n29 = n19 & n28 ;
  assign n30 = ~x8 & ~n21 ;
  assign n31 = x4 ^ x1 ;
  assign n32 = n31 ^ x3 ;
  assign n33 = n32 ^ x5 ;
  assign n34 = x2 ^ x1 ;
  assign n35 = ~x2 & ~n34 ;
  assign n36 = n35 ^ x3 ;
  assign n37 = n36 ^ x2 ;
  assign n38 = n33 & n37 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n39 ^ x2 ;
  assign n41 = ~x5 & ~n40 ;
  assign n42 = n41 ^ x4 ;
  assign n43 = ~n30 & ~n42 ;
  assign n44 = ~n29 & ~n43 ;
  assign y0 = ~n44 ;
endmodule
