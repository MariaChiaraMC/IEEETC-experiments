module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 ;
  assign n17 = x9 & x15 ;
  assign n18 = ~x2 & ~x15 ;
  assign n19 = ~x0 & x7 ;
  assign n20 = x8 & n19 ;
  assign n21 = n18 & n20 ;
  assign n22 = x1 & ~n21 ;
  assign n23 = x3 & ~x6 ;
  assign n24 = ~x1 & ~n23 ;
  assign n25 = n18 & ~n24 ;
  assign n26 = ~x11 & ~x15 ;
  assign n27 = x13 & ~n26 ;
  assign n28 = x13 & x14 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = x0 & ~x3 ;
  assign n31 = n30 ^ x2 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = n30 ^ n19 ;
  assign n34 = n32 & n33 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n35 ^ n27 ;
  assign n37 = n29 & ~n36 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = n38 ^ n30 ;
  assign n40 = n39 ^ n28 ;
  assign n41 = ~n27 & ~n40 ;
  assign n42 = n41 ^ n27 ;
  assign n43 = ~n25 & n42 ;
  assign n44 = x11 & n28 ;
  assign n45 = x4 & x12 ;
  assign n46 = ~x5 & x10 ;
  assign n47 = n45 & n46 ;
  assign n48 = ~n44 & n47 ;
  assign n49 = ~n43 & n48 ;
  assign n50 = ~n22 & n49 ;
  assign n51 = ~n17 & ~n50 ;
  assign y0 = ~n51 ;
endmodule
