module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 ;
  assign n24 = ~x12 & ~x13 ;
  assign n34 = x11 & n24 ;
  assign n63 = ~x6 & n34 ;
  assign n15 = x0 & x4 ;
  assign n16 = x6 & x13 ;
  assign n17 = ~n15 & n16 ;
  assign n18 = n17 ^ x11 ;
  assign n19 = n17 ^ x12 ;
  assign n20 = n19 ^ x12 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = ~x4 & ~x8 ;
  assign n23 = x3 & n22 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n23 & n25 ;
  assign n27 = n26 ^ x12 ;
  assign n28 = n27 ^ n23 ;
  assign n29 = n21 & n28 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n30 ^ n23 ;
  assign n32 = ~n18 & n31 ;
  assign n33 = n32 ^ n17 ;
  assign n35 = n34 ^ n33 ;
  assign n36 = n35 ^ x9 ;
  assign n46 = n36 ^ n35 ;
  assign n37 = x9 & ~x13 ;
  assign n38 = ~x11 & ~n37 ;
  assign n39 = ~x6 & ~n38 ;
  assign n40 = n39 ^ n36 ;
  assign n41 = n40 ^ n35 ;
  assign n42 = n36 ^ n33 ;
  assign n43 = n42 ^ n39 ;
  assign n44 = n43 ^ n41 ;
  assign n45 = n41 & n44 ;
  assign n47 = n46 ^ n45 ;
  assign n48 = n47 ^ n41 ;
  assign n49 = x11 & x12 ;
  assign n50 = x4 & x6 ;
  assign n51 = ~n49 & ~n50 ;
  assign n52 = x0 & n24 ;
  assign n53 = n52 ^ x12 ;
  assign n54 = n51 & n53 ;
  assign n55 = n54 ^ n35 ;
  assign n56 = n45 ^ n41 ;
  assign n57 = n55 & n56 ;
  assign n58 = n57 ^ n35 ;
  assign n59 = ~n48 & n58 ;
  assign n60 = n59 ^ n35 ;
  assign n61 = n60 ^ n34 ;
  assign n62 = n61 ^ n35 ;
  assign n64 = n63 ^ n62 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = ~x9 & n22 ;
  assign n67 = n66 ^ n62 ;
  assign n68 = n67 ^ n62 ;
  assign n69 = n65 & n68 ;
  assign n70 = n69 ^ n62 ;
  assign n71 = x10 & n70 ;
  assign n72 = n71 ^ n62 ;
  assign y0 = n72 ;
endmodule
