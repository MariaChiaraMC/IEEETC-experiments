module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 ;
  assign n87 = x6 & x7 ;
  assign n88 = ~x2 & ~x4 ;
  assign n89 = x3 & n88 ;
  assign n31 = ~x3 & x4 ;
  assign n90 = ~x2 & n31 ;
  assign n91 = ~n89 & ~n90 ;
  assign n92 = n87 & ~n91 ;
  assign n93 = ~x5 & n92 ;
  assign n63 = x5 & ~x6 ;
  assign n94 = n63 & n89 ;
  assign n95 = x0 & ~n94 ;
  assign n99 = x2 & ~x7 ;
  assign n100 = x4 & n99 ;
  assign n96 = x4 & x6 ;
  assign n97 = ~x3 & x5 ;
  assign n98 = ~n96 & n97 ;
  assign n101 = n100 ^ n98 ;
  assign n102 = n101 ^ n95 ;
  assign n103 = ~x3 & ~x6 ;
  assign n104 = ~x5 & ~n103 ;
  assign n105 = n104 ^ n87 ;
  assign n106 = ~n100 & ~n105 ;
  assign n107 = n106 ^ n104 ;
  assign n108 = n102 & ~n107 ;
  assign n109 = n108 ^ n106 ;
  assign n110 = n109 ^ n104 ;
  assign n111 = n110 ^ n100 ;
  assign n112 = n95 & n111 ;
  assign n113 = ~n93 & n112 ;
  assign n114 = x3 & ~x5 ;
  assign n115 = n96 & n114 ;
  assign n116 = ~n94 & ~n115 ;
  assign n117 = x7 & ~n116 ;
  assign n118 = ~x0 & ~n117 ;
  assign n119 = x5 ^ x3 ;
  assign n120 = ~x7 & n96 ;
  assign n121 = n120 ^ x4 ;
  assign n122 = n121 ^ x2 ;
  assign n129 = n122 ^ n121 ;
  assign n123 = n122 ^ n103 ;
  assign n124 = n123 ^ n121 ;
  assign n125 = n122 ^ n120 ;
  assign n126 = n125 ^ n103 ;
  assign n127 = n126 ^ n124 ;
  assign n128 = n124 & n127 ;
  assign n130 = n129 ^ n128 ;
  assign n131 = n130 ^ n124 ;
  assign n132 = n121 ^ n87 ;
  assign n133 = n128 ^ n124 ;
  assign n134 = n132 & n133 ;
  assign n135 = n134 ^ n121 ;
  assign n136 = ~n131 & ~n135 ;
  assign n137 = n136 ^ n121 ;
  assign n138 = n137 ^ x4 ;
  assign n139 = n138 ^ n121 ;
  assign n140 = ~n119 & ~n139 ;
  assign n141 = n118 & ~n140 ;
  assign n142 = ~n113 & ~n141 ;
  assign n9 = ~x0 & x2 ;
  assign n10 = n9 ^ x4 ;
  assign n11 = n10 ^ x3 ;
  assign n12 = n9 ^ x6 ;
  assign n13 = n12 ^ x6 ;
  assign n14 = x5 & x6 ;
  assign n15 = ~x5 & ~x6 ;
  assign n16 = x2 & n15 ;
  assign n17 = ~n14 & ~n16 ;
  assign n18 = x0 & n17 ;
  assign n19 = n18 ^ x6 ;
  assign n20 = ~n13 & ~n19 ;
  assign n21 = n20 ^ x6 ;
  assign n22 = n21 ^ n10 ;
  assign n23 = ~n11 & ~n22 ;
  assign n24 = n23 ^ n20 ;
  assign n25 = n24 ^ x6 ;
  assign n26 = n25 ^ x3 ;
  assign n27 = ~n10 & n26 ;
  assign n28 = n27 ^ n10 ;
  assign n32 = n14 & n31 ;
  assign n33 = n32 ^ x0 ;
  assign n34 = n33 ^ n32 ;
  assign n29 = x7 ^ x2 ;
  assign n30 = ~x2 & n29 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = x6 ^ x5 ;
  assign n37 = n31 ^ x6 ;
  assign n38 = n36 & ~n37 ;
  assign n39 = n38 ^ x5 ;
  assign n40 = n39 ^ x2 ;
  assign n41 = n34 ^ x2 ;
  assign n42 = ~n40 & n41 ;
  assign n43 = n42 ^ n32 ;
  assign n44 = n43 ^ x2 ;
  assign n45 = n44 ^ n39 ;
  assign n46 = n32 ^ x2 ;
  assign n47 = n46 ^ n34 ;
  assign n48 = ~x4 & ~n47 ;
  assign n49 = n48 ^ x7 ;
  assign n50 = n45 & ~n49 ;
  assign n51 = n50 ^ n39 ;
  assign n52 = n51 ^ n34 ;
  assign n53 = n52 ^ x7 ;
  assign n54 = ~n35 & n53 ;
  assign n55 = n54 ^ n42 ;
  assign n56 = n55 ^ x2 ;
  assign n57 = n56 ^ n34 ;
  assign n58 = n57 ^ x7 ;
  assign n59 = n28 & ~n58 ;
  assign n60 = x3 ^ x0 ;
  assign n61 = x5 ^ x4 ;
  assign n62 = n61 ^ x5 ;
  assign n64 = n63 ^ x5 ;
  assign n65 = ~n62 & ~n64 ;
  assign n66 = n65 ^ x5 ;
  assign n67 = n66 ^ x3 ;
  assign n68 = n60 & ~n67 ;
  assign n69 = n68 ^ n65 ;
  assign n70 = n69 ^ x5 ;
  assign n71 = n70 ^ x0 ;
  assign n72 = x3 & ~n71 ;
  assign n73 = n72 ^ x3 ;
  assign n74 = n73 ^ x2 ;
  assign n75 = n74 ^ n73 ;
  assign n76 = n75 ^ x7 ;
  assign n77 = n15 ^ x4 ;
  assign n78 = n15 & ~n77 ;
  assign n79 = n78 ^ n73 ;
  assign n80 = n79 ^ n15 ;
  assign n81 = ~n76 & n80 ;
  assign n82 = n81 ^ n78 ;
  assign n83 = n82 ^ n15 ;
  assign n84 = x7 & n83 ;
  assign n85 = n84 ^ x7 ;
  assign n86 = ~n59 & ~n85 ;
  assign n143 = n142 ^ n86 ;
  assign n144 = n143 ^ n142 ;
  assign n145 = ~x2 & n32 ;
  assign n146 = n145 ^ n142 ;
  assign n147 = n146 ^ n142 ;
  assign n148 = ~n144 & ~n147 ;
  assign n149 = n148 ^ n142 ;
  assign n150 = x1 & ~n149 ;
  assign n151 = n150 ^ n142 ;
  assign y0 = n151 ;
endmodule
