// Benchmark "./pla/b11.pla_res_28NonExact" written by ABC on Fri Nov 20 10:19:55 2020

module \./pla/b11.pla_res_28NonExact  ( 
    x0, x1,
    z0  );
  input  x0, x1;
  output z0;
  assign z0 = ~x0 & x1;
endmodule


