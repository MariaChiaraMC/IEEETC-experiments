module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 ;
  assign n12 = ~x0 & ~x3 ;
  assign n13 = ~x4 & n12 ;
  assign n7 = x0 & x3 ;
  assign n8 = x1 & x4 ;
  assign n9 = n7 & n8 ;
  assign n14 = n13 ^ n9 ;
  assign n15 = n14 ^ n9 ;
  assign n10 = n9 ^ x5 ;
  assign n11 = n10 ^ n9 ;
  assign n16 = n15 ^ n11 ;
  assign n17 = n9 ^ x1 ;
  assign n18 = n17 ^ n9 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n15 & ~n19 ;
  assign n21 = n20 ^ n15 ;
  assign n22 = ~n16 & n21 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n23 ^ n9 ;
  assign n25 = n24 ^ n15 ;
  assign n26 = ~x2 & n25 ;
  assign n27 = n26 ^ n9 ;
  assign y0 = ~n27 ;
endmodule
