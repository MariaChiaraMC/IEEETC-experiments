module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 ;
  assign n11 = ~x0 & ~x6 ;
  assign n12 = ~x1 & ~x2 ;
  assign n13 = n11 & n12 ;
  assign n18 = ~x4 & ~x6 ;
  assign n26 = x2 & ~n18 ;
  assign n27 = ~x1 & ~n26 ;
  assign n28 = x0 & x6 ;
  assign n29 = x4 ^ x3 ;
  assign n30 = n29 ^ x3 ;
  assign n31 = x3 ^ x2 ;
  assign n32 = ~n30 & n31 ;
  assign n33 = n32 ^ x3 ;
  assign n34 = ~x6 & n33 ;
  assign n35 = n34 ^ x4 ;
  assign n36 = ~n28 & ~n35 ;
  assign n37 = ~n27 & ~n36 ;
  assign n14 = ~x1 & ~x3 ;
  assign n15 = x0 & ~n12 ;
  assign n16 = ~n14 & n15 ;
  assign n17 = x2 ^ x1 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = x4 ^ x2 ;
  assign n21 = n20 ^ x4 ;
  assign n22 = ~n19 & n21 ;
  assign n23 = n22 ^ x4 ;
  assign n24 = n17 & n23 ;
  assign n25 = ~n16 & ~n24 ;
  assign n38 = n37 ^ n25 ;
  assign n39 = x7 & n38 ;
  assign n40 = n39 ^ n37 ;
  assign n41 = ~x8 & ~n40 ;
  assign n42 = ~x5 & x7 ;
  assign n43 = x1 & n42 ;
  assign n44 = x3 & ~n43 ;
  assign n45 = n11 & ~n44 ;
  assign n46 = ~n28 & ~n45 ;
  assign n47 = x3 ^ x1 ;
  assign n48 = n47 ^ x3 ;
  assign n49 = x5 ^ x3 ;
  assign n50 = ~n48 & ~n49 ;
  assign n51 = n50 ^ x3 ;
  assign n52 = x6 & n51 ;
  assign n53 = n46 & ~n52 ;
  assign n56 = n53 ^ x7 ;
  assign n57 = n56 ^ n53 ;
  assign n54 = n53 ^ x3 ;
  assign n55 = n54 ^ n53 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = x1 & x4 ;
  assign n60 = n59 ^ n53 ;
  assign n61 = n60 ^ n53 ;
  assign n62 = n61 ^ n57 ;
  assign n63 = n57 & n62 ;
  assign n64 = n63 ^ n57 ;
  assign n65 = ~n58 & n64 ;
  assign n66 = n65 ^ n63 ;
  assign n67 = n66 ^ n53 ;
  assign n68 = n67 ^ n57 ;
  assign n69 = ~x8 & ~n68 ;
  assign n70 = n69 ^ n53 ;
  assign n71 = ~n41 & n70 ;
  assign n72 = ~n13 & n71 ;
  assign y0 = ~n72 ;
endmodule
