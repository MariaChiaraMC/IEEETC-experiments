module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
  assign n16 = ~x8 & ~x11 ;
  assign n17 = ~x0 & n16 ;
  assign n18 = x2 & ~x12 ;
  assign n19 = x7 & ~x13 ;
  assign n20 = n18 & n19 ;
  assign n21 = ~x1 & ~x14 ;
  assign n22 = ~x4 & n21 ;
  assign n23 = n20 & n22 ;
  assign n24 = n17 & n23 ;
  assign n25 = ~x5 & x10 ;
  assign n26 = x9 & n25 ;
  assign n27 = ~x6 & n26 ;
  assign n28 = n27 ^ x3 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = x5 & x6 ;
  assign n31 = ~x9 & n30 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = n29 & n32 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = n24 & n34 ;
  assign y0 = n35 ;
endmodule
