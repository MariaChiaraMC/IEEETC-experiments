// Benchmark "./pla/bcd.div3.pla_res_0NonExact" written by ABC on Fri Nov 20 10:20:12 2020

module \./pla/bcd.div3.pla_res_0NonExact  ( 
    x0, x1,
    z0  );
  input  x0, x1;
  output z0;
  assign z0 = x0 & x1;
endmodule


