module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 ;
  assign n24 = ~x6 & x7 ;
  assign n25 = x5 & n24 ;
  assign n26 = x0 & x4 ;
  assign n27 = ~x3 & ~n26 ;
  assign n28 = x6 & ~x7 ;
  assign n29 = x5 & n28 ;
  assign n30 = n27 & ~n29 ;
  assign n31 = ~n25 & n30 ;
  assign n9 = x7 ^ x6 ;
  assign n10 = x6 ^ x5 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = x7 ^ x3 ;
  assign n13 = n12 ^ x3 ;
  assign n14 = x4 ^ x3 ;
  assign n15 = n13 & ~n14 ;
  assign n16 = n15 ^ x3 ;
  assign n17 = n16 ^ n9 ;
  assign n18 = n11 & n17 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = n20 ^ n10 ;
  assign n22 = n9 & n21 ;
  assign n23 = n22 ^ n9 ;
  assign n32 = n31 ^ n23 ;
  assign n33 = n32 ^ x0 ;
  assign n40 = n33 ^ n32 ;
  assign n34 = n33 ^ x6 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = n31 ^ x6 ;
  assign n37 = n36 ^ x6 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = ~n35 & ~n38 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = n41 ^ n35 ;
  assign n43 = ~x5 & x7 ;
  assign n44 = n43 ^ n32 ;
  assign n45 = n39 ^ n35 ;
  assign n46 = n44 & ~n45 ;
  assign n47 = n46 ^ n32 ;
  assign n48 = n42 & n47 ;
  assign n49 = n48 ^ n32 ;
  assign n50 = n49 ^ n31 ;
  assign n51 = n50 ^ n32 ;
  assign n52 = x1 & n51 ;
  assign n53 = x4 & x5 ;
  assign n54 = ~x0 & x3 ;
  assign n55 = n28 & n54 ;
  assign n56 = n53 & n55 ;
  assign n57 = ~x4 & x7 ;
  assign n58 = ~n24 & ~n57 ;
  assign n59 = ~x1 & ~x3 ;
  assign n60 = x0 & n59 ;
  assign n61 = ~x4 & ~x6 ;
  assign n62 = ~x5 & ~n61 ;
  assign n63 = n60 & n62 ;
  assign n64 = n63 ^ x1 ;
  assign n65 = n64 ^ n63 ;
  assign n66 = ~x5 & x6 ;
  assign n67 = n54 & ~n66 ;
  assign n68 = ~x4 & ~x5 ;
  assign n69 = n67 & ~n68 ;
  assign n70 = n69 ^ n63 ;
  assign n71 = n70 ^ n63 ;
  assign n72 = ~n65 & n71 ;
  assign n73 = n72 ^ n63 ;
  assign n74 = n58 & n73 ;
  assign n75 = n74 ^ n63 ;
  assign n76 = ~n56 & ~n75 ;
  assign n77 = ~n52 & n76 ;
  assign n78 = ~x2 & ~n77 ;
  assign n79 = x5 ^ x4 ;
  assign n80 = x2 & n28 ;
  assign n81 = n80 ^ x5 ;
  assign n82 = n81 ^ n80 ;
  assign n83 = n80 ^ n24 ;
  assign n84 = n83 ^ n80 ;
  assign n85 = ~n82 & n84 ;
  assign n86 = n85 ^ n80 ;
  assign n87 = ~n79 & n86 ;
  assign n88 = n87 ^ n80 ;
  assign n89 = n88 ^ x2 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = n88 ^ n61 ;
  assign n92 = n91 ^ n88 ;
  assign n93 = n90 & n92 ;
  assign n94 = n93 ^ n88 ;
  assign n95 = x3 & n94 ;
  assign n96 = n95 ^ n88 ;
  assign n99 = n96 ^ n80 ;
  assign n100 = n99 ^ n96 ;
  assign n97 = n96 ^ n68 ;
  assign n98 = n97 ^ n96 ;
  assign n101 = n100 ^ n98 ;
  assign n102 = n96 ^ x3 ;
  assign n103 = n102 ^ n96 ;
  assign n104 = n103 ^ n100 ;
  assign n105 = n100 & ~n104 ;
  assign n106 = n105 ^ n100 ;
  assign n107 = n101 & n106 ;
  assign n108 = n107 ^ n105 ;
  assign n109 = n108 ^ n96 ;
  assign n110 = n109 ^ n100 ;
  assign n111 = ~x1 & n110 ;
  assign n112 = n111 ^ n96 ;
  assign n113 = ~x0 & n112 ;
  assign n114 = ~n78 & ~n113 ;
  assign y0 = ~n114 ;
endmodule
