module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n10 = ~x2 & ~x6 ;
  assign n11 = ~x4 & n10 ;
  assign n13 = x5 & n11 ;
  assign n14 = ~x6 & ~x7 ;
  assign n15 = x3 & ~n14 ;
  assign n16 = ~x4 & n15 ;
  assign n17 = ~n13 & ~n16 ;
  assign n18 = x4 ^ x2 ;
  assign n19 = ~x3 & n18 ;
  assign n20 = n18 ^ x5 ;
  assign n21 = ~x4 & ~x6 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n20 & n22 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n19 & n24 ;
  assign n26 = n25 ^ x2 ;
  assign n27 = n17 & ~n26 ;
  assign n9 = ~x3 & ~x5 ;
  assign n12 = n9 & n11 ;
  assign n28 = n27 ^ n12 ;
  assign n29 = n12 ^ x7 ;
  assign n30 = n12 ^ x1 ;
  assign n31 = n12 & ~n30 ;
  assign n32 = n31 ^ n12 ;
  assign n33 = ~n29 & n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n34 ^ n12 ;
  assign n36 = n35 ^ x1 ;
  assign n37 = ~n28 & ~n36 ;
  assign n38 = n37 ^ n12 ;
  assign y0 = n38 ;
endmodule
