module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 ;
  assign n9 = x2 ^ x1 ;
  assign n7 = x4 ^ x3 ;
  assign n8 = n7 ^ x0 ;
  assign n10 = n9 ^ n8 ;
  assign n11 = n10 ^ n7 ;
  assign n15 = n8 ^ x4 ;
  assign n12 = n7 ^ x2 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = n13 ^ n7 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n16 ^ n8 ;
  assign n18 = n9 & ~n17 ;
  assign n19 = n18 ^ n7 ;
  assign n20 = n19 ^ n11 ;
  assign n21 = n14 ^ n9 ;
  assign n22 = n21 ^ n11 ;
  assign n23 = ~n7 & n22 ;
  assign n24 = n23 ^ n9 ;
  assign n25 = ~n20 & n24 ;
  assign n26 = n11 & n25 ;
  assign n27 = n26 ^ n18 ;
  assign n28 = n27 ^ n23 ;
  assign n29 = n28 ^ n25 ;
  assign n30 = n29 ^ n7 ;
  assign n36 = n30 ^ x0 ;
  assign n37 = n36 ^ n30 ;
  assign n31 = ~x3 & ~x4 ;
  assign n32 = x3 & x4 ;
  assign n33 = ~n31 & ~n32 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ n30 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = ~x1 & x2 ;
  assign n40 = x1 & ~x2 ;
  assign n41 = ~n39 & ~n40 ;
  assign n42 = n41 ^ n30 ;
  assign n43 = n42 ^ n30 ;
  assign n44 = n43 ^ n37 ;
  assign n45 = n37 & ~n44 ;
  assign n46 = n45 ^ n37 ;
  assign n47 = n38 & n46 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = n48 ^ n30 ;
  assign n50 = n49 ^ n37 ;
  assign n51 = ~x5 & ~n50 ;
  assign n52 = n51 ^ n30 ;
  assign y0 = ~n52 ;
endmodule
