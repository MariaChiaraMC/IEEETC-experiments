module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n13 = ~x2 & ~x8 ;
  assign n14 = ~x2 & x3 ;
  assign n15 = x8 & ~n14 ;
  assign n16 = ~x4 & ~n15 ;
  assign n17 = ~n13 & ~n16 ;
  assign n18 = x7 & ~n17 ;
  assign n19 = x2 & ~x3 ;
  assign n20 = x8 ^ x7 ;
  assign n22 = x8 ^ x4 ;
  assign n21 = x8 ^ x2 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n23 ^ n20 ;
  assign n25 = n22 ^ x8 ;
  assign n26 = x10 ^ x3 ;
  assign n27 = n22 ^ n20 ;
  assign n28 = ~n26 & n27 ;
  assign n29 = n28 ^ x3 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n25 & n30 ;
  assign n32 = n31 ^ n22 ;
  assign n33 = ~n24 & ~n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = ~n20 & n34 ;
  assign n36 = n35 ^ x7 ;
  assign n37 = ~n19 & n36 ;
  assign n38 = ~n18 & n37 ;
  assign y0 = n38 ;
endmodule
