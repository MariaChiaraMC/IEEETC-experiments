module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 ;
  output y0 ;
  wire n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 ;
  assign n26 = ~x15 & ~x16 ;
  assign n27 = x5 & ~x17 ;
  assign n28 = ~x2 & ~x3 ;
  assign n29 = ~x4 & n28 ;
  assign n30 = ~n27 & n29 ;
  assign n31 = x17 ^ x14 ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = n26 & ~n32 ;
  assign n34 = x1 & ~n33 ;
  assign n35 = x15 & x17 ;
  assign n36 = x16 & n35 ;
  assign n37 = ~x5 & x24 ;
  assign n38 = ~x2 & ~x14 ;
  assign n39 = ~x3 & ~x4 ;
  assign n40 = n38 & n39 ;
  assign n41 = n37 & n40 ;
  assign n42 = n36 & n41 ;
  assign n43 = x13 & n42 ;
  assign n44 = ~x1 & n29 ;
  assign n45 = ~x5 & n44 ;
  assign n46 = x13 & n26 ;
  assign n47 = ~n45 & n46 ;
  assign n48 = ~n43 & ~n47 ;
  assign n49 = ~n34 & ~n48 ;
  assign n50 = ~x13 & x14 ;
  assign n51 = n36 & ~n44 ;
  assign n52 = x24 & n45 ;
  assign n53 = n26 & n52 ;
  assign n54 = ~n51 & ~n53 ;
  assign n55 = n50 & ~n54 ;
  assign n56 = ~n49 & ~n55 ;
  assign n57 = ~x0 & ~n56 ;
  assign n58 = x4 ^ x0 ;
  assign n59 = x5 & ~n58 ;
  assign n60 = n59 ^ x0 ;
  assign n61 = x14 & n60 ;
  assign n62 = n36 ^ n26 ;
  assign n63 = n62 ^ n36 ;
  assign n64 = n36 ^ x17 ;
  assign n65 = n64 ^ n36 ;
  assign n66 = n63 & ~n65 ;
  assign n67 = n66 ^ n36 ;
  assign n68 = x13 & n67 ;
  assign n69 = n68 ^ n36 ;
  assign n70 = n61 & n69 ;
  assign n71 = ~x14 & x17 ;
  assign n72 = x0 & ~x5 ;
  assign n73 = n71 & n72 ;
  assign n74 = ~x4 & n73 ;
  assign n75 = n46 & n74 ;
  assign n76 = ~n70 & ~n75 ;
  assign n77 = ~x1 & n28 ;
  assign n78 = ~n76 & n77 ;
  assign n79 = ~n57 & ~n78 ;
  assign n80 = ~x10 & ~n79 ;
  assign n81 = ~x13 & x19 ;
  assign n82 = x18 & x21 ;
  assign n83 = n81 & n82 ;
  assign n84 = ~x20 & n83 ;
  assign n85 = x13 & ~x22 ;
  assign n86 = x10 & ~n85 ;
  assign n87 = ~x0 & n86 ;
  assign n88 = n52 & n87 ;
  assign n89 = ~n84 & n88 ;
  assign n90 = ~n80 & ~n89 ;
  assign n91 = x11 & ~n90 ;
  assign n92 = ~x4 & ~x17 ;
  assign n93 = x10 & ~x11 ;
  assign n94 = n92 & n93 ;
  assign n95 = ~x0 & ~x1 ;
  assign n96 = x15 & n95 ;
  assign n97 = n28 & n96 ;
  assign n98 = n94 & n97 ;
  assign n99 = x14 ^ x13 ;
  assign n100 = n37 & n99 ;
  assign n101 = n100 ^ x16 ;
  assign n102 = n101 ^ n100 ;
  assign n103 = x5 & ~x13 ;
  assign n104 = ~x14 & n103 ;
  assign n105 = n104 ^ n100 ;
  assign n106 = ~n102 & n105 ;
  assign n107 = n106 ^ n100 ;
  assign n108 = n98 & n107 ;
  assign n109 = ~n91 & ~n108 ;
  assign n110 = ~x12 & ~n109 ;
  assign n111 = x10 & x13 ;
  assign n112 = x12 & n111 ;
  assign n113 = n95 & n112 ;
  assign n114 = x11 & n41 ;
  assign n115 = n113 & n114 ;
  assign n116 = ~x15 & n115 ;
  assign n117 = ~n110 & ~n116 ;
  assign n118 = ~x6 & ~x23 ;
  assign n119 = ~x8 & n118 ;
  assign n120 = ~x7 & n119 ;
  assign n121 = ~x9 & n120 ;
  assign n122 = ~n117 & n121 ;
  assign y0 = n122 ;
endmodule
