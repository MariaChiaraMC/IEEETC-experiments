module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 ;
  assign n7 = x1 & ~x5 ;
  assign n8 = x2 & ~x5 ;
  assign n9 = x2 & ~x3 ;
  assign n10 = ~n8 & ~n9 ;
  assign n11 = ~n7 & ~n10 ;
  assign n12 = ~x4 & x5 ;
  assign n13 = ~x3 & n12 ;
  assign n14 = ~n11 & ~n13 ;
  assign n15 = ~x0 & ~n14 ;
  assign n16 = x2 ^ x0 ;
  assign n17 = n16 ^ x5 ;
  assign n24 = n17 ^ x3 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = n18 ^ x3 ;
  assign n20 = x4 ^ x3 ;
  assign n21 = n20 ^ x5 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = ~n19 & ~n22 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ n19 ;
  assign n27 = x3 ^ x0 ;
  assign n28 = n27 ^ x3 ;
  assign n29 = n23 ^ n19 ;
  assign n30 = n28 & ~n29 ;
  assign n31 = n30 ^ x3 ;
  assign n32 = ~n26 & n31 ;
  assign n33 = n32 ^ x3 ;
  assign n34 = n33 ^ x3 ;
  assign n35 = n34 ^ x1 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = n36 ^ n15 ;
  assign n38 = ~x2 & ~x5 ;
  assign n39 = n38 ^ x2 ;
  assign n40 = n39 ^ x2 ;
  assign n41 = n16 ^ x2 ;
  assign n42 = n40 & n41 ;
  assign n43 = n42 ^ x2 ;
  assign n44 = x3 & n43 ;
  assign n45 = n44 ^ x2 ;
  assign n46 = n45 ^ x4 ;
  assign n47 = n45 & ~n46 ;
  assign n48 = n47 ^ n34 ;
  assign n49 = n48 ^ n45 ;
  assign n50 = n37 & n49 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = n51 ^ n45 ;
  assign n53 = ~n15 & n52 ;
  assign n54 = n53 ^ n15 ;
  assign y0 = n54 ;
endmodule
