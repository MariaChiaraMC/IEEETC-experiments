// Benchmark "./pla/Z5xp1.pla_res_8NonExact" written by ABC on Fri Nov 20 10:31:40 2020

module \./pla/Z5xp1.pla_res_8NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = x0;
endmodule


