module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 ;
  assign n20 = ~x0 & x2 ;
  assign n21 = ~x13 & ~x14 ;
  assign n22 = x15 & ~n21 ;
  assign n23 = x4 & ~x5 ;
  assign n24 = ~n22 & n23 ;
  assign n25 = ~x1 & n24 ;
  assign n26 = x10 & n25 ;
  assign n27 = x1 & x5 ;
  assign n28 = x4 & ~x16 ;
  assign n29 = ~x18 & ~n28 ;
  assign n30 = ~n22 & ~n29 ;
  assign n31 = n27 & n30 ;
  assign n32 = ~x17 & n31 ;
  assign n33 = ~n26 & ~n32 ;
  assign n34 = n20 & ~n33 ;
  assign n35 = x1 & x11 ;
  assign n36 = n23 & n35 ;
  assign n37 = x13 & x14 ;
  assign n38 = x15 & n37 ;
  assign n39 = ~x2 & x10 ;
  assign n40 = ~x17 & n39 ;
  assign n41 = ~n38 & n40 ;
  assign n42 = n36 & n41 ;
  assign n43 = ~x0 & n42 ;
  assign n44 = n43 ^ n34 ;
  assign n45 = ~x17 & n20 ;
  assign n46 = n27 & n45 ;
  assign n47 = ~n29 & ~n37 ;
  assign n48 = n46 & n47 ;
  assign n49 = ~x2 & ~x9 ;
  assign n50 = ~x1 & n49 ;
  assign n51 = n50 ^ x7 ;
  assign n52 = n51 ^ n48 ;
  assign n55 = ~x16 & n46 ;
  assign n53 = ~x17 & n23 ;
  assign n54 = ~n38 & n53 ;
  assign n56 = n55 ^ n54 ;
  assign n57 = ~n50 & ~n56 ;
  assign n58 = n57 ^ n54 ;
  assign n59 = ~n52 & ~n58 ;
  assign n60 = n59 ^ n57 ;
  assign n61 = n60 ^ n54 ;
  assign n62 = n61 ^ n50 ;
  assign n63 = ~n48 & n62 ;
  assign n64 = n63 ^ x3 ;
  assign n65 = n64 ^ n63 ;
  assign n66 = x6 & n55 ;
  assign n67 = ~x1 & x6 ;
  assign n68 = ~x8 & ~n67 ;
  assign n69 = ~n25 & n68 ;
  assign n70 = x0 & ~n69 ;
  assign n71 = ~x2 & n70 ;
  assign n72 = ~n66 & ~n71 ;
  assign n73 = n72 ^ n63 ;
  assign n74 = ~n65 & n73 ;
  assign n75 = n74 ^ n63 ;
  assign n76 = n75 ^ n34 ;
  assign n77 = n44 & ~n76 ;
  assign n78 = n77 ^ n74 ;
  assign n79 = n78 ^ n63 ;
  assign n80 = n79 ^ n43 ;
  assign n81 = ~n34 & ~n80 ;
  assign n82 = n81 ^ n34 ;
  assign n83 = x12 & n82 ;
  assign y0 = n83 ;
endmodule
