module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 ;
  assign n13 = x7 & ~x11 ;
  assign n14 = ~x9 & x10 ;
  assign n15 = x8 & n14 ;
  assign n16 = n13 & ~n15 ;
  assign n17 = x5 & ~n16 ;
  assign n18 = x11 ^ x4 ;
  assign n19 = n18 ^ x0 ;
  assign n20 = x4 ^ x0 ;
  assign n21 = x8 ^ x5 ;
  assign n22 = n20 & n21 ;
  assign n23 = n22 ^ x5 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = x7 & ~n24 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = ~n19 & ~n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = ~x0 & n28 ;
  assign n30 = n29 ^ x0 ;
  assign n31 = n30 ^ n17 ;
  assign n32 = ~x5 & n14 ;
  assign n33 = x7 & ~x8 ;
  assign n34 = x4 & ~n33 ;
  assign n35 = n32 & ~n34 ;
  assign n36 = n35 ^ x6 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = x4 & ~n32 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = ~n37 & n39 ;
  assign n41 = n40 ^ n35 ;
  assign n42 = n41 ^ n17 ;
  assign n43 = n31 & ~n42 ;
  assign n44 = n43 ^ n40 ;
  assign n45 = n44 ^ n35 ;
  assign n46 = n45 ^ n30 ;
  assign n47 = ~n17 & ~n46 ;
  assign n48 = n47 ^ n17 ;
  assign y0 = ~n48 ;
endmodule
