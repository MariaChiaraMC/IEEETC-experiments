module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 ;
  assign n15 = x4 ^ x2 ;
  assign n22 = n15 ^ x2 ;
  assign n16 = n15 ^ x6 ;
  assign n17 = n16 ^ x2 ;
  assign n18 = x6 ^ x1 ;
  assign n19 = n18 ^ x6 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = ~n17 & ~n20 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n23 ^ n17 ;
  assign n25 = x3 ^ x2 ;
  assign n26 = n21 ^ n17 ;
  assign n27 = n25 & ~n26 ;
  assign n28 = n27 ^ x2 ;
  assign n29 = n24 & ~n28 ;
  assign n30 = n29 ^ x2 ;
  assign n31 = n30 ^ x4 ;
  assign n32 = n31 ^ x2 ;
  assign n33 = x5 & ~n32 ;
  assign n34 = x2 & ~x12 ;
  assign n35 = ~x11 & n34 ;
  assign n36 = x8 & ~x10 ;
  assign n37 = x5 & x6 ;
  assign n38 = n36 & n37 ;
  assign n39 = ~x7 & ~x13 ;
  assign n40 = n38 & n39 ;
  assign n41 = n35 & n40 ;
  assign n42 = x2 & ~x4 ;
  assign n43 = x3 & ~n42 ;
  assign n44 = ~n41 & n43 ;
  assign n45 = x9 & ~n44 ;
  assign n46 = ~n33 & n45 ;
  assign n47 = ~x4 & ~x6 ;
  assign n48 = ~x2 & ~x5 ;
  assign n49 = n47 & n48 ;
  assign n50 = ~x3 & ~n49 ;
  assign n51 = ~x1 & ~n50 ;
  assign n52 = ~x0 & ~n51 ;
  assign n53 = n46 & n52 ;
  assign y0 = n53 ;
endmodule
