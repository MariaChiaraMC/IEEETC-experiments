module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n11 = x4 & ~x8 ;
  assign n12 = x0 & x2 ;
  assign n13 = ~x6 & ~x7 ;
  assign n14 = ~n12 & n13 ;
  assign n15 = ~x1 & ~n14 ;
  assign n16 = ~n11 & ~n15 ;
  assign n17 = ~x4 & x8 ;
  assign n18 = ~x2 & x6 ;
  assign n19 = ~x5 & x9 ;
  assign n20 = ~n18 & ~n19 ;
  assign n21 = ~n17 & n20 ;
  assign n22 = n11 ^ x3 ;
  assign n23 = n22 ^ x3 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n15 ^ x7 ;
  assign n26 = x3 & ~n25 ;
  assign n27 = n26 ^ x7 ;
  assign n28 = n24 & ~n27 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = n29 ^ x7 ;
  assign n31 = n30 ^ x3 ;
  assign n32 = n21 & ~n31 ;
  assign n33 = ~n16 & n32 ;
  assign y0 = n33 ;
endmodule
