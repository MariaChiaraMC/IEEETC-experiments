module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 ;
  output y0 ;
  wire n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 ;
  assign n32 = x0 & ~x24 ;
  assign n34 = ~x11 & ~x13 ;
  assign n35 = x2 & x10 ;
  assign n36 = n34 & n35 ;
  assign n37 = ~x12 & n36 ;
  assign n38 = ~x8 & ~n37 ;
  assign n40 = n38 ^ x26 ;
  assign n49 = n40 ^ n38 ;
  assign n33 = ~x2 & ~x4 ;
  assign n39 = n38 ^ n33 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = n42 ^ n38 ;
  assign n44 = ~x4 & ~x9 ;
  assign n45 = n44 ^ n41 ;
  assign n46 = n45 ^ n41 ;
  assign n47 = n46 ^ n43 ;
  assign n48 = ~n43 & n47 ;
  assign n50 = n49 ^ n48 ;
  assign n51 = n50 ^ n43 ;
  assign n52 = n38 ^ x5 ;
  assign n53 = n48 ^ n43 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = n54 ^ n38 ;
  assign n56 = ~n51 & n55 ;
  assign n57 = n56 ^ n38 ;
  assign n58 = n57 ^ x26 ;
  assign n59 = n58 ^ n38 ;
  assign n60 = n32 & n59 ;
  assign n61 = ~x3 & x5 ;
  assign n62 = ~x7 & ~n61 ;
  assign n63 = ~n33 & ~n62 ;
  assign n64 = n63 ^ x5 ;
  assign n65 = n63 ^ x0 ;
  assign n66 = n65 ^ n63 ;
  assign n67 = ~n64 & n66 ;
  assign n68 = n67 ^ x5 ;
  assign n78 = x4 ^ x2 ;
  assign n79 = n78 ^ x22 ;
  assign n80 = n79 ^ x4 ;
  assign n85 = n80 ^ n78 ;
  assign n86 = n85 ^ x4 ;
  assign n87 = n86 ^ x4 ;
  assign n88 = n78 ^ x29 ;
  assign n89 = n88 ^ n78 ;
  assign n90 = n89 ^ x4 ;
  assign n91 = ~n87 & ~n90 ;
  assign n81 = n78 ^ x28 ;
  assign n82 = n81 ^ n80 ;
  assign n83 = n82 ^ x4 ;
  assign n84 = ~n80 & n83 ;
  assign n92 = n91 ^ n84 ;
  assign n93 = n92 ^ n80 ;
  assign n94 = n84 ^ x4 ;
  assign n95 = n94 ^ n86 ;
  assign n96 = ~x4 & ~n95 ;
  assign n97 = n96 ^ n84 ;
  assign n98 = ~n93 & n97 ;
  assign n99 = n98 ^ n91 ;
  assign n100 = n99 ^ n96 ;
  assign n101 = n100 ^ n80 ;
  assign n102 = n101 ^ x4 ;
  assign n103 = n102 ^ n86 ;
  assign n104 = n103 ^ x2 ;
  assign n69 = ~x7 & x30 ;
  assign n70 = n69 ^ n63 ;
  assign n71 = n70 ^ n65 ;
  assign n72 = n71 ^ x3 ;
  assign n73 = n72 ^ n71 ;
  assign n74 = n71 ^ n65 ;
  assign n75 = n74 ^ n63 ;
  assign n76 = n75 ^ n67 ;
  assign n77 = n73 & ~n76 ;
  assign n105 = n104 ^ n77 ;
  assign n106 = ~x5 & n105 ;
  assign n107 = n106 ^ n77 ;
  assign n108 = n107 ^ n66 ;
  assign n109 = ~n68 & n108 ;
  assign n110 = n109 ^ n77 ;
  assign n111 = n110 ^ n106 ;
  assign n112 = n111 ^ n66 ;
  assign n113 = n112 ^ x0 ;
  assign n114 = ~x27 & n113 ;
  assign n115 = x23 ^ x0 ;
  assign n116 = x24 & n115 ;
  assign n117 = ~n114 & ~n116 ;
  assign n118 = ~x25 & ~n117 ;
  assign n119 = x22 & x28 ;
  assign n120 = x2 & ~n119 ;
  assign n121 = ~x5 & n120 ;
  assign n122 = n62 & ~n121 ;
  assign n123 = n32 & ~n122 ;
  assign n124 = ~n118 & ~n123 ;
  assign n125 = x3 & x5 ;
  assign n126 = ~n33 & ~n125 ;
  assign n127 = ~x5 & ~x6 ;
  assign n128 = n69 & ~n127 ;
  assign n129 = n128 ^ x24 ;
  assign n130 = n129 ^ n126 ;
  assign n160 = x3 & ~x25 ;
  assign n161 = n33 & n160 ;
  assign n162 = ~x27 & n161 ;
  assign n131 = ~x19 & ~x20 ;
  assign n132 = x14 & x18 ;
  assign n133 = ~n131 & ~n132 ;
  assign n134 = x0 & x21 ;
  assign n135 = ~x15 & ~n134 ;
  assign n136 = ~n133 & n135 ;
  assign n137 = ~x17 & ~n136 ;
  assign n138 = x16 ^ x15 ;
  assign n139 = n138 ^ x16 ;
  assign n140 = n139 ^ x18 ;
  assign n147 = n140 ^ n138 ;
  assign n141 = n140 ^ x18 ;
  assign n142 = n141 ^ n138 ;
  assign n143 = x18 ^ x0 ;
  assign n144 = n143 ^ x18 ;
  assign n145 = n144 ^ n142 ;
  assign n146 = ~n142 & ~n145 ;
  assign n148 = n147 ^ n146 ;
  assign n149 = n148 ^ n142 ;
  assign n150 = n138 ^ x17 ;
  assign n151 = n146 ^ n142 ;
  assign n152 = ~n150 & ~n151 ;
  assign n153 = n152 ^ n138 ;
  assign n154 = ~n149 & ~n153 ;
  assign n155 = n154 ^ n138 ;
  assign n156 = n155 ^ x18 ;
  assign n157 = n156 ^ n138 ;
  assign n158 = ~n137 & ~n157 ;
  assign n159 = x3 & ~n158 ;
  assign n163 = n162 ^ n159 ;
  assign n164 = ~x24 & n163 ;
  assign n165 = n164 ^ n162 ;
  assign n166 = ~n130 & n165 ;
  assign n167 = n166 ^ n164 ;
  assign n168 = n167 ^ n162 ;
  assign n169 = n168 ^ x24 ;
  assign n170 = ~n126 & ~n169 ;
  assign n171 = n124 & ~n170 ;
  assign n172 = ~x26 & ~n171 ;
  assign n173 = ~x1 & ~n172 ;
  assign n174 = ~n60 & n173 ;
  assign y0 = ~n174 ;
endmodule
