module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n13 = x4 & ~x11 ;
  assign n14 = ~x5 & ~x10 ;
  assign n15 = ~n13 & ~n14 ;
  assign n16 = x5 & ~x7 ;
  assign n17 = ~x0 & ~n16 ;
  assign n18 = ~x6 & n17 ;
  assign n19 = ~n15 & n18 ;
  assign n20 = x7 & ~x11 ;
  assign n21 = ~x5 & n20 ;
  assign n22 = x11 ^ x4 ;
  assign n23 = n22 ^ x4 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = ~x8 & ~x9 ;
  assign n26 = n25 ^ x10 ;
  assign n27 = x4 & ~n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n24 & n28 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n30 ^ n25 ;
  assign n32 = n31 ^ x4 ;
  assign n33 = ~n21 & n32 ;
  assign n34 = n19 & n33 ;
  assign y0 = n34 ;
endmodule
