module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 ;
  assign n9 = x2 ^ x1 ;
  assign n10 = x4 & x5 ;
  assign n11 = ~x3 & n10 ;
  assign n12 = n11 ^ x2 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = ~x4 & ~x5 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = n13 & n15 ;
  assign n17 = n16 ^ n11 ;
  assign n18 = n9 & n17 ;
  assign n19 = ~x6 & n18 ;
  assign n20 = x1 & ~x2 ;
  assign n21 = ~x3 & x4 ;
  assign n22 = x5 & x7 ;
  assign n23 = n21 & ~n22 ;
  assign n24 = x6 & ~n23 ;
  assign n25 = ~x5 & x7 ;
  assign n26 = ~n10 & ~n25 ;
  assign n27 = ~x2 & ~n26 ;
  assign n28 = n24 & n27 ;
  assign n29 = x4 ^ x3 ;
  assign n31 = n29 ^ x4 ;
  assign n32 = n31 ^ x5 ;
  assign n39 = n32 ^ n29 ;
  assign n30 = n29 ^ x5 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ n29 ;
  assign n35 = n29 ^ x6 ;
  assign n36 = n35 ^ n30 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = ~n34 & n37 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = n40 ^ n34 ;
  assign n42 = n29 ^ x7 ;
  assign n43 = n38 ^ n34 ;
  assign n44 = ~n42 & ~n43 ;
  assign n45 = n44 ^ n29 ;
  assign n46 = n41 & n45 ;
  assign n47 = n46 ^ n29 ;
  assign n48 = n47 ^ n29 ;
  assign n49 = n48 ^ n29 ;
  assign n50 = x1 & n49 ;
  assign n51 = ~x2 & x3 ;
  assign n52 = n14 & n51 ;
  assign n53 = ~x7 & n52 ;
  assign n54 = ~n50 & ~n53 ;
  assign n55 = ~n28 & n54 ;
  assign n56 = ~n20 & ~n55 ;
  assign n57 = ~n19 & ~n56 ;
  assign n60 = n57 ^ n22 ;
  assign n61 = n60 ^ n57 ;
  assign n58 = n57 ^ n51 ;
  assign n59 = n58 ^ n57 ;
  assign n62 = n61 ^ n59 ;
  assign n63 = x4 & ~x6 ;
  assign n64 = ~x1 & n63 ;
  assign n65 = n64 ^ n57 ;
  assign n66 = n65 ^ n57 ;
  assign n67 = n66 ^ n61 ;
  assign n68 = n61 & n67 ;
  assign n69 = n68 ^ n61 ;
  assign n70 = n62 & n69 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = n71 ^ n57 ;
  assign n73 = n72 ^ n61 ;
  assign n74 = x0 & ~n73 ;
  assign n75 = n74 ^ n57 ;
  assign y0 = ~n75 ;
endmodule
