module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n8 = x3 ^ x0 ;
  assign n10 = n8 ^ x1 ;
  assign n11 = n10 ^ x5 ;
  assign n7 = x5 ^ x3 ;
  assign n12 = n11 ^ n7 ;
  assign n16 = n12 ^ n8 ;
  assign n9 = n8 ^ n7 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = n9 & n13 ;
  assign n15 = n14 ^ n9 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n7 ^ x5 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n18 ^ x4 ;
  assign n21 = n19 & ~n20 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = n22 ^ x2 ;
  assign n24 = n19 ^ x2 ;
  assign n25 = ~n18 & ~n24 ;
  assign n26 = n25 ^ n18 ;
  assign n27 = n26 ^ n16 ;
  assign n28 = ~n23 & n27 ;
  assign n29 = n28 ^ x2 ;
  assign n30 = ~n17 & ~n29 ;
  assign y0 = n30 ;
endmodule
