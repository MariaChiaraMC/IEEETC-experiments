module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 ;
  assign n16 = x13 ^ x7 ;
  assign n17 = x6 & ~x14 ;
  assign n18 = ~x1 & x3 ;
  assign n19 = ~x7 & x9 ;
  assign n20 = n18 & n19 ;
  assign n24 = ~x0 & x2 ;
  assign n25 = ~x8 & x10 ;
  assign n26 = x4 & n25 ;
  assign n27 = n24 & n26 ;
  assign n21 = x8 & ~x10 ;
  assign n22 = ~x4 & n21 ;
  assign n23 = x0 & n22 ;
  assign n28 = n27 ^ n23 ;
  assign n29 = ~x5 & n28 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n20 & n30 ;
  assign n32 = n17 & n31 ;
  assign n33 = n32 ^ n16 ;
  assign n34 = n33 ^ x13 ;
  assign n35 = n34 ^ n33 ;
  assign n36 = ~x9 & ~x10 ;
  assign n37 = n17 & n36 ;
  assign n38 = ~x8 & n37 ;
  assign n39 = ~x1 & n24 ;
  assign n40 = ~x4 & x5 ;
  assign n41 = n39 & n40 ;
  assign n42 = x3 & x13 ;
  assign n43 = n41 & n42 ;
  assign n44 = n38 & n43 ;
  assign n45 = n44 ^ n33 ;
  assign n46 = n45 ^ n16 ;
  assign n47 = ~n35 & ~n46 ;
  assign n48 = n47 ^ n44 ;
  assign n49 = x6 ^ x4 ;
  assign n50 = n49 ^ x14 ;
  assign n51 = n24 ^ x4 ;
  assign n52 = n51 ^ n24 ;
  assign n53 = ~x0 & ~x2 ;
  assign n54 = ~x9 & n53 ;
  assign n55 = n54 ^ n24 ;
  assign n56 = n52 & n55 ;
  assign n57 = n56 ^ n24 ;
  assign n58 = n57 ^ n49 ;
  assign n59 = ~n50 & ~n58 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = n60 ^ n24 ;
  assign n62 = n61 ^ x14 ;
  assign n63 = ~n49 & n62 ;
  assign n64 = n63 ^ n49 ;
  assign n65 = n25 & ~n64 ;
  assign n66 = ~x2 & ~x8 ;
  assign n67 = x0 & ~x4 ;
  assign n68 = ~n66 & n67 ;
  assign n69 = n37 & n68 ;
  assign n70 = ~n65 & ~n69 ;
  assign n71 = n18 & ~n70 ;
  assign n72 = x4 & x14 ;
  assign n73 = x6 & n72 ;
  assign n74 = x1 & n73 ;
  assign n75 = x3 & n74 ;
  assign n76 = ~x1 & ~x3 ;
  assign n77 = n38 & n76 ;
  assign n78 = n67 & n77 ;
  assign n79 = n75 & ~n78 ;
  assign n80 = n78 ^ x0 ;
  assign n81 = ~x8 & x9 ;
  assign n82 = ~x10 & n81 ;
  assign n83 = n82 ^ n79 ;
  assign n84 = n80 & n83 ;
  assign n85 = n84 ^ n82 ;
  assign n86 = n79 & n85 ;
  assign n87 = n86 ^ n78 ;
  assign n88 = ~x2 & n87 ;
  assign n89 = ~n71 & ~n88 ;
  assign n90 = ~x5 & ~n89 ;
  assign n91 = ~x9 & n26 ;
  assign n92 = ~n22 & ~n91 ;
  assign n93 = x5 & ~x6 ;
  assign n94 = n53 & n76 ;
  assign n95 = n93 & n94 ;
  assign n96 = ~n92 & n95 ;
  assign n97 = ~x14 & n96 ;
  assign n98 = ~n90 & ~n97 ;
  assign n99 = ~n44 & n98 ;
  assign n100 = n99 ^ n16 ;
  assign n101 = ~n48 & n100 ;
  assign n102 = n101 ^ n99 ;
  assign n103 = n16 & n102 ;
  assign n104 = n103 ^ n47 ;
  assign n105 = n104 ^ x7 ;
  assign n106 = n105 ^ n44 ;
  assign n109 = n106 ^ n93 ;
  assign n110 = n109 ^ n106 ;
  assign n107 = n106 ^ n39 ;
  assign n108 = n107 ^ n106 ;
  assign n111 = n110 ^ n108 ;
  assign n112 = ~x3 & x4 ;
  assign n113 = n81 & n112 ;
  assign n114 = ~x13 & ~x14 ;
  assign n115 = x10 & n114 ;
  assign n116 = n113 & n115 ;
  assign n117 = n116 ^ n106 ;
  assign n118 = n117 ^ n106 ;
  assign n119 = n118 ^ n110 ;
  assign n120 = n110 & n119 ;
  assign n121 = n120 ^ n110 ;
  assign n122 = n111 & n121 ;
  assign n123 = n122 ^ n120 ;
  assign n124 = n123 ^ n106 ;
  assign n125 = n124 ^ n110 ;
  assign n126 = x12 & ~n125 ;
  assign n127 = n126 ^ n106 ;
  assign n128 = ~x11 & ~n127 ;
  assign y0 = n128 ;
endmodule
