module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 ;
  assign n9 = x3 ^ x2 ;
  assign n10 = x4 & ~x5 ;
  assign n11 = n10 ^ x3 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = x6 ^ x5 ;
  assign n14 = x7 ^ x4 ;
  assign n15 = x6 ^ x4 ;
  assign n16 = ~n14 & ~n15 ;
  assign n17 = n16 ^ x4 ;
  assign n18 = ~n13 & n17 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = n19 ^ n10 ;
  assign n21 = ~n12 & n20 ;
  assign n22 = n21 ^ n10 ;
  assign n23 = ~n9 & ~n22 ;
  assign n24 = n23 ^ x2 ;
  assign n25 = ~x1 & ~n24 ;
  assign n26 = ~x0 & ~n25 ;
  assign y0 = n26 ;
endmodule
