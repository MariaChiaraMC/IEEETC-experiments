module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 ;
  assign n11 = ~x2 & ~x6 ;
  assign n12 = ~x0 & n11 ;
  assign n13 = ~x3 & ~x7 ;
  assign n14 = n12 & n13 ;
  assign n15 = x8 & ~n14 ;
  assign n16 = ~x1 & x4 ;
  assign n17 = ~n15 & n16 ;
  assign n18 = x2 & x3 ;
  assign n19 = x6 ^ x0 ;
  assign n20 = n18 & n19 ;
  assign n21 = n20 ^ n12 ;
  assign n22 = n21 ^ x7 ;
  assign n29 = n22 ^ n21 ;
  assign n23 = n22 ^ x8 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n22 ^ n20 ;
  assign n26 = n25 ^ x8 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n24 & ~n27 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = n30 ^ n24 ;
  assign n32 = n21 ^ x3 ;
  assign n33 = n28 ^ n24 ;
  assign n34 = ~n32 & n33 ;
  assign n35 = n34 ^ n21 ;
  assign n36 = ~n31 & n35 ;
  assign n37 = n36 ^ n21 ;
  assign n38 = n37 ^ n12 ;
  assign n39 = n38 ^ n21 ;
  assign n40 = n17 & n39 ;
  assign n41 = n40 ^ x9 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = x4 & ~x8 ;
  assign n44 = ~x4 & x8 ;
  assign n45 = x6 ^ x2 ;
  assign n46 = x1 & ~n45 ;
  assign n47 = n46 ^ n13 ;
  assign n48 = x3 & x7 ;
  assign n49 = n48 ^ n46 ;
  assign n50 = n49 ^ n48 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = n12 ^ x8 ;
  assign n53 = ~x8 & ~n52 ;
  assign n54 = n53 ^ n48 ;
  assign n55 = n54 ^ x8 ;
  assign n56 = ~n51 & n55 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n57 ^ x8 ;
  assign n59 = n47 & ~n58 ;
  assign n60 = n59 ^ n46 ;
  assign n61 = ~n44 & n60 ;
  assign n62 = ~n43 & n61 ;
  assign n63 = n62 ^ n40 ;
  assign n64 = n42 & n63 ;
  assign n65 = n64 ^ n40 ;
  assign n66 = x5 & n65 ;
  assign n67 = ~x5 & ~x9 ;
  assign n68 = n60 & n67 ;
  assign n69 = x8 ^ x4 ;
  assign n70 = n68 & ~n69 ;
  assign n71 = ~n66 & ~n70 ;
  assign y0 = ~n71 ;
endmodule
