module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 ;
  assign n7 = x0 & x1 ;
  assign n8 = ~x3 & ~x5 ;
  assign n9 = n7 & n8 ;
  assign n14 = x4 & ~x5 ;
  assign n27 = x3 & ~x5 ;
  assign n28 = x1 & ~n27 ;
  assign n29 = ~n14 & n28 ;
  assign n30 = ~x4 & ~x5 ;
  assign n31 = ~n7 & n30 ;
  assign n32 = ~x1 & ~x5 ;
  assign n33 = ~x0 & ~n32 ;
  assign n34 = ~x3 & n33 ;
  assign n35 = ~n31 & ~n34 ;
  assign n36 = ~n29 & ~n35 ;
  assign n11 = x5 ^ x0 ;
  assign n10 = x5 ^ x3 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = n12 ^ n11 ;
  assign n16 = x5 ^ x1 ;
  assign n17 = n16 ^ n11 ;
  assign n18 = ~n11 & n17 ;
  assign n21 = n18 ^ n14 ;
  assign n15 = n14 ^ n13 ;
  assign n19 = n18 ^ n11 ;
  assign n20 = ~n15 & ~n19 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = ~n13 & n22 ;
  assign n24 = n23 ^ n18 ;
  assign n25 = n24 ^ n20 ;
  assign n26 = n25 ^ x1 ;
  assign n37 = n36 ^ n26 ;
  assign n38 = ~x2 & n37 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = ~n9 & n39 ;
  assign y0 = ~n40 ;
endmodule
