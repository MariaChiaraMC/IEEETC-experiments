module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 ;
  assign n73 = x3 ^ x2 ;
  assign n15 = x1 & ~x8 ;
  assign n19 = ~x0 & x2 ;
  assign n20 = x3 & n19 ;
  assign n16 = x2 & ~x3 ;
  assign n17 = ~x6 & ~n16 ;
  assign n18 = ~x5 & ~n17 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = x0 & ~x3 ;
  assign n23 = n22 ^ n18 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = x6 ^ x5 ;
  assign n26 = x7 & ~n25 ;
  assign n27 = n26 ^ x5 ;
  assign n28 = ~x4 & ~n27 ;
  assign n29 = n28 ^ n22 ;
  assign n30 = ~n24 & n29 ;
  assign n31 = n30 ^ n22 ;
  assign n32 = n21 & n31 ;
  assign n33 = n32 ^ n20 ;
  assign n34 = n15 & n33 ;
  assign n35 = x1 & ~n22 ;
  assign n36 = ~x5 & ~x7 ;
  assign n37 = n36 ^ x1 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = n36 ^ x6 ;
  assign n40 = n39 ^ n36 ;
  assign n41 = ~n38 & n40 ;
  assign n42 = n41 ^ n36 ;
  assign n43 = ~x3 & ~n42 ;
  assign n44 = n43 ^ n36 ;
  assign n45 = ~n35 & n44 ;
  assign n46 = n45 ^ x2 ;
  assign n47 = x5 & ~x7 ;
  assign n48 = x1 & n47 ;
  assign n49 = ~x6 & ~n48 ;
  assign n50 = x4 & ~x8 ;
  assign n51 = ~n49 & n50 ;
  assign n52 = n51 ^ x0 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = x5 & x8 ;
  assign n55 = ~x4 & n54 ;
  assign n56 = n55 ^ n51 ;
  assign n57 = ~n53 & n56 ;
  assign n58 = n57 ^ n51 ;
  assign n59 = n58 ^ n45 ;
  assign n60 = ~n46 & n59 ;
  assign n61 = n60 ^ n57 ;
  assign n62 = n61 ^ n51 ;
  assign n63 = n62 ^ x2 ;
  assign n64 = n45 & ~n63 ;
  assign n65 = n64 ^ n45 ;
  assign n66 = ~n34 & ~n65 ;
  assign n67 = ~x10 & ~x11 ;
  assign n68 = ~n66 & n67 ;
  assign n74 = n73 ^ n68 ;
  assign n75 = n74 ^ n68 ;
  assign n69 = x10 & x11 ;
  assign n70 = x13 & n69 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = n71 ^ n68 ;
  assign n76 = n75 ^ n72 ;
  assign n77 = n68 ^ x8 ;
  assign n78 = n77 ^ n68 ;
  assign n79 = n78 ^ n75 ;
  assign n80 = n75 & ~n79 ;
  assign n81 = n80 ^ n75 ;
  assign n82 = n76 & n81 ;
  assign n83 = n82 ^ n80 ;
  assign n84 = n83 ^ n68 ;
  assign n85 = n84 ^ n75 ;
  assign n86 = x9 & n85 ;
  assign n87 = n86 ^ n68 ;
  assign n88 = ~x12 & n87 ;
  assign y0 = n88 ;
endmodule
