module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 ;
  assign n17 = ~x12 & ~x13 ;
  assign n18 = ~x0 & n17 ;
  assign n71 = ~x3 & ~x5 ;
  assign n19 = ~x7 & ~x8 ;
  assign n20 = x4 & ~x9 ;
  assign n21 = ~x6 & n20 ;
  assign n22 = n19 & n21 ;
  assign n23 = x10 & ~x15 ;
  assign n24 = x3 & x5 ;
  assign n25 = ~x1 & x2 ;
  assign n26 = n24 & n25 ;
  assign n27 = n23 & n26 ;
  assign n28 = n22 & n27 ;
  assign n29 = ~x1 & ~x4 ;
  assign n30 = x5 ^ x3 ;
  assign n31 = ~x2 & n23 ;
  assign n32 = ~x6 & n31 ;
  assign n33 = n32 ^ x5 ;
  assign n34 = n33 ^ n32 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = ~x15 & n19 ;
  assign n37 = x2 & ~n36 ;
  assign n38 = x6 & ~x10 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = ~n37 & ~n39 ;
  assign n41 = n40 ^ n32 ;
  assign n42 = n41 ^ n37 ;
  assign n43 = n35 & ~n42 ;
  assign n44 = n43 ^ n40 ;
  assign n45 = n44 ^ n37 ;
  assign n46 = ~n30 & ~n45 ;
  assign n47 = n29 & n46 ;
  assign n48 = x4 & x15 ;
  assign n49 = x3 & ~x8 ;
  assign n50 = n48 & n49 ;
  assign n51 = x1 & n50 ;
  assign n53 = ~x5 & ~n38 ;
  assign n52 = x6 & x10 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = n53 ^ x7 ;
  assign n56 = n55 ^ n53 ;
  assign n57 = n56 ^ n51 ;
  assign n58 = n57 ^ n50 ;
  assign n59 = ~n54 & ~n58 ;
  assign n60 = n59 ^ n53 ;
  assign n61 = n51 & ~n60 ;
  assign n62 = n61 ^ n51 ;
  assign n63 = ~n47 & ~n62 ;
  assign n64 = x7 & x8 ;
  assign n65 = ~x2 & ~n64 ;
  assign n66 = x9 & ~n65 ;
  assign n67 = ~n63 & n66 ;
  assign n68 = ~n28 & ~n67 ;
  assign n72 = n71 ^ n68 ;
  assign n73 = n72 ^ n68 ;
  assign n69 = n68 ^ n31 ;
  assign n70 = n69 ^ n68 ;
  assign n74 = n73 ^ n70 ;
  assign n75 = x8 & x9 ;
  assign n76 = n29 & n75 ;
  assign n77 = x6 & ~x7 ;
  assign n78 = x11 & n77 ;
  assign n79 = n76 & n78 ;
  assign n80 = n79 ^ n68 ;
  assign n81 = n80 ^ n68 ;
  assign n82 = n81 ^ n73 ;
  assign n83 = n73 & n82 ;
  assign n84 = n83 ^ n73 ;
  assign n85 = n74 & n84 ;
  assign n86 = n85 ^ n83 ;
  assign n87 = n86 ^ n68 ;
  assign n88 = n87 ^ n73 ;
  assign n89 = x14 & ~n88 ;
  assign n90 = n89 ^ n68 ;
  assign n91 = n18 & ~n90 ;
  assign y0 = n91 ;
endmodule
