module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 ;
  assign n8 = x0 & x1 ;
  assign n9 = x3 & x6 ;
  assign n10 = x5 & ~n9 ;
  assign n11 = ~x5 & n9 ;
  assign n12 = ~n10 & ~n11 ;
  assign n13 = ~n8 & ~n12 ;
  assign n14 = ~x2 & n13 ;
  assign n15 = n14 ^ x4 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = ~x0 & x2 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = n18 ^ n15 ;
  assign n25 = n19 ^ n15 ;
  assign n26 = n25 ^ n14 ;
  assign n20 = n19 ^ x5 ;
  assign n21 = n20 ^ x6 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n22 ^ n14 ;
  assign n24 = n23 ^ n16 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = ~n16 & ~n27 ;
  assign n29 = n28 ^ n22 ;
  assign n30 = n29 ^ n26 ;
  assign n36 = n20 ^ n19 ;
  assign n31 = n20 ^ x3 ;
  assign n32 = n31 ^ n20 ;
  assign n33 = n26 ^ n22 ;
  assign n34 = n32 & n33 ;
  assign n35 = n34 ^ n28 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = n37 ^ n32 ;
  assign n39 = n38 ^ n22 ;
  assign n40 = n26 & ~n39 ;
  assign n41 = n40 ^ n16 ;
  assign n42 = n30 & ~n41 ;
  assign n43 = n42 ^ n16 ;
  assign n44 = n43 ^ x4 ;
  assign n45 = n44 ^ n16 ;
  assign y0 = ~n45 ;
endmodule
