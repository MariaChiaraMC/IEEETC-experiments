module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 ;
  assign n11 = x4 ^ x3 ;
  assign n17 = x7 ^ x5 ;
  assign n9 = x5 ^ x3 ;
  assign n18 = n17 ^ n9 ;
  assign n19 = n18 ^ x5 ;
  assign n10 = n9 ^ x6 ;
  assign n12 = n11 ^ n10 ;
  assign n20 = n19 ^ n12 ;
  assign n21 = n20 ^ n11 ;
  assign n22 = ~n11 & n21 ;
  assign n23 = n22 ^ n9 ;
  assign n24 = n23 ^ n12 ;
  assign n25 = n24 ^ n11 ;
  assign n26 = n25 ^ x5 ;
  assign n27 = n12 ^ n11 ;
  assign n28 = n27 ^ x5 ;
  assign n29 = ~n24 & ~n28 ;
  assign n30 = n29 ^ n9 ;
  assign n31 = n30 ^ n12 ;
  assign n32 = n31 ^ n11 ;
  assign n33 = n32 ^ x5 ;
  assign n34 = ~n26 & ~n33 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = n13 ^ n11 ;
  assign n15 = n14 ^ x5 ;
  assign n16 = n14 & ~n15 ;
  assign n35 = n34 ^ n16 ;
  assign n36 = n35 ^ n22 ;
  assign n37 = n36 ^ n9 ;
  assign n38 = n37 ^ n12 ;
  assign n39 = n38 ^ n11 ;
  assign n40 = n39 ^ x5 ;
  assign n41 = n40 ^ x3 ;
  assign y0 = ~n41 ;
endmodule
