module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n7 = x1 ^ x0 ;
  assign n8 = n7 ^ x1 ;
  assign n9 = n8 ^ x2 ;
  assign n10 = n9 ^ x3 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = n9 ^ n8 ;
  assign n13 = n12 ^ n7 ;
  assign n14 = ~n11 & n13 ;
  assign n15 = n14 ^ n8 ;
  assign n16 = x4 & x5 ;
  assign n17 = n8 & ~n16 ;
  assign n18 = n17 ^ n7 ;
  assign n19 = n15 & ~n18 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = ~n7 & n20 ;
  assign n22 = n21 ^ n14 ;
  assign n23 = n22 ^ x0 ;
  assign n24 = n23 ^ n8 ;
  assign y0 = n24 ;
endmodule
