module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 ;
  output y0 ;
  wire n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 ;
  assign n35 = ~x3 & ~x4 ;
  assign n36 = x0 & ~x13 ;
  assign n37 = ~n35 & n36 ;
  assign n58 = x4 ^ x0 ;
  assign n80 = n58 ^ x4 ;
  assign n81 = n80 ^ x4 ;
  assign n82 = n80 & ~n81 ;
  assign n61 = ~x4 & x13 ;
  assign n62 = x15 ^ x14 ;
  assign n63 = x17 ^ x15 ;
  assign n64 = ~n62 & ~n63 ;
  assign n65 = x23 & n64 ;
  assign n66 = n61 & ~n65 ;
  assign n67 = x20 & x21 ;
  assign n45 = x16 & ~x18 ;
  assign n68 = x17 & n45 ;
  assign n69 = x19 & ~n68 ;
  assign n44 = ~x13 & ~x15 ;
  assign n70 = x4 & n44 ;
  assign n71 = ~n69 & n70 ;
  assign n72 = ~n67 & n71 ;
  assign n73 = ~n66 & ~n72 ;
  assign n59 = x4 ^ x3 ;
  assign n60 = n59 ^ n58 ;
  assign n74 = n73 ^ n60 ;
  assign n75 = n74 ^ n60 ;
  assign n76 = n60 ^ n58 ;
  assign n77 = n76 ^ x4 ;
  assign n78 = ~n75 & ~n77 ;
  assign n85 = n82 ^ n78 ;
  assign n79 = n78 ^ x2 ;
  assign n83 = n82 ^ n80 ;
  assign n84 = ~n79 & n83 ;
  assign n86 = n85 ^ n84 ;
  assign n87 = ~x2 & n86 ;
  assign n88 = n87 ^ n78 ;
  assign n89 = n88 ^ n82 ;
  assign n90 = n89 ^ n84 ;
  assign n91 = n90 ^ x0 ;
  assign n92 = ~x5 & ~n91 ;
  assign n38 = x4 & ~x13 ;
  assign n39 = x21 & ~x22 ;
  assign n40 = n38 & n39 ;
  assign n41 = n40 ^ x3 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = n42 ^ x2 ;
  assign n46 = ~x4 & n45 ;
  assign n47 = n44 & n46 ;
  assign n48 = n47 ^ x0 ;
  assign n49 = ~n47 & n48 ;
  assign n50 = n49 ^ n40 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = n43 & n51 ;
  assign n53 = n52 ^ n49 ;
  assign n54 = n53 ^ n47 ;
  assign n55 = x2 & ~n54 ;
  assign n56 = n55 ^ x2 ;
  assign n57 = x5 & ~n56 ;
  assign n93 = n92 ^ n57 ;
  assign n94 = n93 ^ x2 ;
  assign n95 = n94 ^ n57 ;
  assign n163 = n95 ^ n93 ;
  assign n164 = n163 ^ n57 ;
  assign n165 = n164 ^ n57 ;
  assign n166 = ~x3 & x13 ;
  assign n167 = x4 & x14 ;
  assign n168 = n166 & n167 ;
  assign n169 = n168 ^ n93 ;
  assign n170 = n169 ^ n93 ;
  assign n171 = n170 ^ n57 ;
  assign n172 = n165 & ~n171 ;
  assign n96 = x10 ^ x9 ;
  assign n97 = n96 ^ x9 ;
  assign n98 = n97 ^ x7 ;
  assign n99 = x12 ^ x9 ;
  assign n100 = x9 ^ x8 ;
  assign n101 = n100 ^ x9 ;
  assign n102 = n99 & n101 ;
  assign n103 = n102 ^ x9 ;
  assign n104 = n103 ^ n97 ;
  assign n105 = n104 ^ x7 ;
  assign n106 = ~x11 & ~n105 ;
  assign n107 = n106 ^ x9 ;
  assign n108 = n107 ^ n97 ;
  assign n109 = n98 & ~n108 ;
  assign n110 = n109 ^ n106 ;
  assign n111 = x7 & n110 ;
  assign n112 = x6 & ~n111 ;
  assign n113 = x27 & x29 ;
  assign n114 = x28 & x31 ;
  assign n115 = n113 & n114 ;
  assign n116 = ~x30 & n115 ;
  assign n117 = ~x13 & n116 ;
  assign n118 = ~n112 & ~n117 ;
  assign n119 = n35 & ~n118 ;
  assign n120 = x25 & x26 ;
  assign n121 = x3 & x17 ;
  assign n122 = n120 & n121 ;
  assign n123 = x13 & n122 ;
  assign n125 = x24 ^ x17 ;
  assign n133 = n125 ^ x24 ;
  assign n134 = n133 ^ x24 ;
  assign n135 = n133 & n134 ;
  assign n124 = n120 ^ x24 ;
  assign n126 = n125 ^ n124 ;
  assign n127 = n126 ^ n67 ;
  assign n128 = n127 ^ n126 ;
  assign n129 = n126 ^ n125 ;
  assign n130 = n129 ^ x24 ;
  assign n131 = n128 & ~n130 ;
  assign n138 = n135 ^ n131 ;
  assign n132 = n131 ^ x13 ;
  assign n136 = n135 ^ n133 ;
  assign n137 = ~n132 & n136 ;
  assign n139 = n138 ^ n137 ;
  assign n140 = ~x13 & n139 ;
  assign n141 = n140 ^ n131 ;
  assign n142 = n141 ^ n135 ;
  assign n143 = n142 ^ n137 ;
  assign n144 = n143 ^ x17 ;
  assign n145 = x4 & n144 ;
  assign n146 = x15 & ~x18 ;
  assign n147 = x19 & x32 ;
  assign n148 = ~n146 & n147 ;
  assign n149 = n38 & ~n148 ;
  assign n150 = ~n145 & ~n149 ;
  assign n151 = n150 ^ x3 ;
  assign n152 = n151 ^ n150 ;
  assign n153 = x14 & n38 ;
  assign n154 = n153 ^ n150 ;
  assign n155 = ~n152 & ~n154 ;
  assign n156 = n155 ^ n150 ;
  assign n157 = ~n123 & n156 ;
  assign n158 = ~n119 & n157 ;
  assign n159 = n158 ^ n93 ;
  assign n160 = n159 ^ n95 ;
  assign n161 = n160 ^ n57 ;
  assign n162 = n95 & n161 ;
  assign n173 = n172 ^ n162 ;
  assign n174 = n173 ^ n95 ;
  assign n175 = n162 ^ n57 ;
  assign n176 = n175 ^ n164 ;
  assign n177 = ~n57 & n176 ;
  assign n178 = n177 ^ n162 ;
  assign n179 = n174 & n178 ;
  assign n180 = n179 ^ n172 ;
  assign n181 = n180 ^ n177 ;
  assign n182 = n181 ^ n95 ;
  assign n183 = n182 ^ n57 ;
  assign n184 = n183 ^ n164 ;
  assign n185 = n184 ^ n92 ;
  assign n186 = x0 & ~x3 ;
  assign n187 = n186 ^ x2 ;
  assign n188 = n186 ^ n61 ;
  assign n189 = n188 ^ n61 ;
  assign n190 = n38 & n121 ;
  assign n191 = x33 & n190 ;
  assign n192 = n191 ^ n61 ;
  assign n193 = ~n189 & ~n192 ;
  assign n194 = n193 ^ n61 ;
  assign n195 = ~n187 & n194 ;
  assign n196 = n195 ^ x2 ;
  assign n197 = n185 & n196 ;
  assign n198 = ~n37 & n197 ;
  assign n199 = x1 & ~n198 ;
  assign y0 = n199 ;
endmodule
