module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 ;
  assign n47 = x7 ^ x0 ;
  assign n22 = ~x8 & x10 ;
  assign n23 = ~x9 & ~x11 ;
  assign n24 = ~x12 & n23 ;
  assign n25 = n22 & n24 ;
  assign n26 = x14 & x15 ;
  assign n27 = x14 ^ x13 ;
  assign n28 = n27 ^ x15 ;
  assign n29 = n26 & n28 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = n25 & n30 ;
  assign n17 = ~x6 & ~x7 ;
  assign n18 = x3 & ~n17 ;
  assign n19 = x4 & n18 ;
  assign n32 = n31 ^ n19 ;
  assign n33 = n32 ^ n19 ;
  assign n20 = n19 ^ x6 ;
  assign n21 = n20 ^ n19 ;
  assign n34 = n33 ^ n21 ;
  assign n35 = n19 ^ x3 ;
  assign n36 = n35 ^ n19 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n33 & ~n37 ;
  assign n39 = n38 ^ n33 ;
  assign n40 = n34 & n39 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n41 ^ n19 ;
  assign n43 = n42 ^ n33 ;
  assign n44 = x5 & n43 ;
  assign n45 = n44 ^ n19 ;
  assign n46 = n45 ^ x0 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = n48 ^ x3 ;
  assign n50 = n49 ^ n48 ;
  assign n51 = n48 ^ n46 ;
  assign n52 = n51 ^ x0 ;
  assign n53 = ~n50 & ~n52 ;
  assign n54 = n53 ^ n46 ;
  assign n55 = ~x4 & x5 ;
  assign n56 = n31 & ~n55 ;
  assign n57 = ~n46 & n56 ;
  assign n58 = n57 ^ x0 ;
  assign n59 = ~n54 & ~n58 ;
  assign n60 = n59 ^ n57 ;
  assign n61 = ~x0 & n60 ;
  assign n62 = n61 ^ n53 ;
  assign n63 = n62 ^ n45 ;
  assign n64 = n63 ^ n46 ;
  assign y0 = ~n64 ;
endmodule
