module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 ;
  assign n28 = ~x5 & ~x6 ;
  assign n11 = x0 & ~x9 ;
  assign n12 = ~x2 & ~n11 ;
  assign n13 = x6 ^ x5 ;
  assign n14 = n13 ^ x6 ;
  assign n15 = x6 ^ x2 ;
  assign n16 = n15 ^ x8 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = x9 ^ x2 ;
  assign n19 = x2 & n18 ;
  assign n20 = n19 ^ x8 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = ~n17 & n21 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n23 ^ x2 ;
  assign n25 = ~n14 & n24 ;
  assign n26 = n25 ^ n13 ;
  assign n27 = ~n12 & n26 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ x7 ;
  assign n39 = n30 ^ n29 ;
  assign n31 = ~x8 & ~x9 ;
  assign n32 = x0 & ~n31 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ n29 ;
  assign n35 = n30 ^ n27 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = n34 & ~n37 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = n40 ^ n34 ;
  assign n42 = n29 ^ x2 ;
  assign n43 = n38 ^ n34 ;
  assign n44 = ~n42 & n43 ;
  assign n45 = n44 ^ n29 ;
  assign n46 = ~n41 & n45 ;
  assign n47 = n46 ^ n29 ;
  assign n48 = n47 ^ n28 ;
  assign n49 = n48 ^ n29 ;
  assign n50 = x3 & n49 ;
  assign n53 = ~x6 & x9 ;
  assign n54 = x5 & n53 ;
  assign n55 = ~x3 & n54 ;
  assign n51 = n31 ^ x7 ;
  assign n52 = n51 ^ n31 ;
  assign n56 = n55 ^ n52 ;
  assign n57 = n56 ^ n55 ;
  assign n58 = x5 & ~x6 ;
  assign n59 = ~x5 & x6 ;
  assign n60 = ~x3 & x4 ;
  assign n61 = n59 & n60 ;
  assign n62 = ~n58 & ~n61 ;
  assign n63 = n57 ^ n51 ;
  assign n64 = n63 ^ n57 ;
  assign n65 = ~n62 & ~n64 ;
  assign n66 = n65 ^ n55 ;
  assign n67 = x4 & n28 ;
  assign n68 = x1 & n67 ;
  assign n69 = n68 ^ n55 ;
  assign n70 = n63 & ~n69 ;
  assign n71 = n70 ^ n57 ;
  assign n72 = n71 ^ n63 ;
  assign n73 = ~n66 & ~n72 ;
  assign n74 = ~n57 & n73 ;
  assign n75 = n74 ^ n65 ;
  assign n76 = n75 ^ x7 ;
  assign n77 = ~x2 & ~n76 ;
  assign n78 = ~n50 & ~n77 ;
  assign y0 = ~n78 ;
endmodule
