module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 ;
  assign n17 = x6 & x7 ;
  assign n18 = x4 & ~n17 ;
  assign n19 = x12 & ~x13 ;
  assign n20 = ~x14 & n19 ;
  assign n21 = ~x12 & ~x15 ;
  assign n22 = x13 & n21 ;
  assign n23 = ~n20 & ~n22 ;
  assign n24 = n23 ^ x5 ;
  assign n26 = ~x12 & x13 ;
  assign n27 = x14 & ~n26 ;
  assign n25 = x15 & ~n19 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n28 ^ x7 ;
  assign n30 = n23 ^ x7 ;
  assign n31 = n30 ^ x7 ;
  assign n32 = ~n29 & n31 ;
  assign n33 = n32 ^ x7 ;
  assign n34 = n24 & n33 ;
  assign n35 = n34 ^ x5 ;
  assign n36 = n18 & ~n35 ;
  assign n37 = x5 ^ x4 ;
  assign n38 = n37 ^ x10 ;
  assign n39 = x7 ^ x4 ;
  assign n40 = n39 ^ x7 ;
  assign n43 = x14 & x15 ;
  assign n44 = n26 & n43 ;
  assign n45 = x12 & x13 ;
  assign n46 = x15 ^ x14 ;
  assign n47 = n45 & n46 ;
  assign n48 = ~n44 & ~n47 ;
  assign n52 = n48 ^ n19 ;
  assign n49 = n48 ^ x7 ;
  assign n41 = x14 & ~x15 ;
  assign n42 = n41 ^ n19 ;
  assign n50 = n49 ^ n42 ;
  assign n51 = n50 ^ n19 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n48 ^ n42 ;
  assign n55 = n54 ^ n19 ;
  assign n56 = n55 ^ n19 ;
  assign n57 = ~n50 & ~n56 ;
  assign n58 = n57 ^ n50 ;
  assign n59 = ~n55 & ~n58 ;
  assign n60 = n59 ^ n19 ;
  assign n61 = ~n53 & n60 ;
  assign n62 = n61 ^ n57 ;
  assign n63 = n62 ^ n19 ;
  assign n64 = n63 ^ n52 ;
  assign n65 = n64 ^ x7 ;
  assign n66 = n40 & n65 ;
  assign n67 = n66 ^ x7 ;
  assign n68 = n67 ^ n37 ;
  assign n69 = ~n38 & n68 ;
  assign n70 = n69 ^ n66 ;
  assign n71 = n70 ^ x7 ;
  assign n72 = n71 ^ x10 ;
  assign n73 = ~n37 & ~n72 ;
  assign n74 = n73 ^ n37 ;
  assign n75 = n74 ^ x10 ;
  assign n76 = x6 & n75 ;
  assign n77 = n76 ^ x7 ;
  assign n78 = ~n19 & ~n26 ;
  assign n79 = n43 & ~n78 ;
  assign n80 = ~n47 & ~n79 ;
  assign n81 = ~x4 & x5 ;
  assign n82 = ~n80 & n81 ;
  assign n83 = ~x10 & ~n82 ;
  assign n84 = n83 ^ n77 ;
  assign n85 = n84 ^ n76 ;
  assign n86 = n85 ^ n84 ;
  assign n87 = ~x6 & x10 ;
  assign n88 = n87 ^ x5 ;
  assign n89 = ~x4 & ~x5 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = n90 ^ n87 ;
  assign n92 = n91 ^ n90 ;
  assign n93 = n46 ^ x15 ;
  assign n94 = n93 ^ n45 ;
  assign n95 = n21 ^ x13 ;
  assign n96 = n21 & ~n95 ;
  assign n97 = n96 ^ x15 ;
  assign n98 = n97 ^ n21 ;
  assign n99 = n94 & n98 ;
  assign n100 = n99 ^ n96 ;
  assign n101 = n100 ^ n21 ;
  assign n102 = ~n45 & n101 ;
  assign n103 = n102 ^ n45 ;
  assign n104 = ~x4 & ~n103 ;
  assign n105 = x9 ^ x8 ;
  assign n106 = n104 & n105 ;
  assign n107 = n80 & ~n106 ;
  assign n108 = x8 & ~x9 ;
  assign n109 = ~x6 & ~n108 ;
  assign n110 = ~x4 & x9 ;
  assign n111 = n109 & ~n110 ;
  assign n112 = ~n80 & n111 ;
  assign n113 = n112 ^ x10 ;
  assign n114 = n113 ^ n112 ;
  assign n115 = ~x8 & x9 ;
  assign n116 = ~n108 & ~n115 ;
  assign n117 = x6 ^ x4 ;
  assign n118 = ~n116 & ~n117 ;
  assign n119 = n118 ^ x4 ;
  assign n120 = n119 ^ n112 ;
  assign n121 = ~n114 & n120 ;
  assign n122 = n121 ^ n112 ;
  assign n123 = ~n107 & n122 ;
  assign n124 = n123 ^ n90 ;
  assign n125 = n124 ^ n88 ;
  assign n126 = n92 & ~n125 ;
  assign n127 = n126 ^ n123 ;
  assign n128 = ~x9 & n104 ;
  assign n129 = ~x8 & n128 ;
  assign n130 = ~n123 & ~n129 ;
  assign n131 = n130 ^ n88 ;
  assign n132 = ~n127 & ~n131 ;
  assign n133 = n132 ^ n130 ;
  assign n134 = ~n88 & n133 ;
  assign n135 = n134 ^ n126 ;
  assign n136 = n135 ^ x5 ;
  assign n137 = n136 ^ n123 ;
  assign n138 = n137 ^ n84 ;
  assign n139 = n138 ^ n77 ;
  assign n140 = n86 & ~n139 ;
  assign n141 = n140 ^ n137 ;
  assign n142 = ~x14 & x15 ;
  assign n143 = ~x12 & n142 ;
  assign n144 = ~x13 & n41 ;
  assign n145 = ~n143 & ~n144 ;
  assign n146 = ~x4 & ~n145 ;
  assign n147 = n23 & ~n146 ;
  assign n148 = x5 & ~n147 ;
  assign n149 = ~x5 & ~n103 ;
  assign n150 = n80 & ~n149 ;
  assign n151 = x4 & ~n150 ;
  assign n152 = n105 & n151 ;
  assign n153 = ~n148 & ~n152 ;
  assign n154 = n137 & n153 ;
  assign n155 = n154 ^ n77 ;
  assign n156 = n141 & ~n155 ;
  assign n157 = n156 ^ n154 ;
  assign n158 = ~n77 & n157 ;
  assign n159 = n158 ^ n140 ;
  assign n160 = n159 ^ x7 ;
  assign n161 = n160 ^ n137 ;
  assign n162 = ~x11 & n161 ;
  assign n163 = n17 & n108 ;
  assign n164 = n89 & n163 ;
  assign n165 = x6 & ~x10 ;
  assign n166 = x11 ^ x4 ;
  assign n167 = n165 & ~n166 ;
  assign n168 = n167 ^ x4 ;
  assign n169 = ~n80 & ~n168 ;
  assign n170 = ~n104 & ~n169 ;
  assign n171 = n170 ^ x7 ;
  assign n172 = n171 ^ n170 ;
  assign n173 = n172 ^ x5 ;
  assign n174 = x6 & n21 ;
  assign n175 = ~x6 & n108 ;
  assign n176 = n142 & n175 ;
  assign n177 = x12 & n176 ;
  assign n178 = ~n174 & ~n177 ;
  assign n179 = x10 & x13 ;
  assign n180 = ~n178 & n179 ;
  assign n181 = n145 & ~n180 ;
  assign n182 = x10 & x14 ;
  assign n183 = n182 ^ n175 ;
  assign n184 = n78 ^ x15 ;
  assign n185 = n184 ^ n78 ;
  assign n186 = n78 ^ x12 ;
  assign n187 = ~n185 & ~n186 ;
  assign n188 = n187 ^ n78 ;
  assign n189 = n188 ^ n182 ;
  assign n190 = n183 & ~n189 ;
  assign n191 = n190 ^ n187 ;
  assign n192 = n191 ^ n78 ;
  assign n193 = n192 ^ n175 ;
  assign n194 = n182 & ~n193 ;
  assign n195 = n194 ^ n182 ;
  assign n196 = n181 & ~n195 ;
  assign n197 = x4 & ~n196 ;
  assign n198 = n111 & n129 ;
  assign n199 = x4 & ~n109 ;
  assign n200 = n199 ^ n80 ;
  assign n201 = n199 ^ n111 ;
  assign n202 = n201 ^ n111 ;
  assign n203 = x6 & n22 ;
  assign n204 = n203 ^ n111 ;
  assign n205 = n202 & ~n204 ;
  assign n206 = n205 ^ n111 ;
  assign n207 = ~n200 & ~n206 ;
  assign n208 = n207 ^ n80 ;
  assign n209 = ~n198 & n208 ;
  assign n210 = ~x10 & ~n209 ;
  assign n211 = x10 & ~n80 ;
  assign n212 = n211 ^ x6 ;
  assign n213 = n211 ^ n20 ;
  assign n214 = n213 ^ n20 ;
  assign n215 = n108 ^ n20 ;
  assign n216 = n214 & n215 ;
  assign n217 = n216 ^ n20 ;
  assign n218 = n212 & ~n217 ;
  assign n219 = n218 ^ x6 ;
  assign n220 = x4 & n219 ;
  assign n221 = ~n210 & ~n220 ;
  assign n222 = x11 & ~n221 ;
  assign n223 = n222 ^ n197 ;
  assign n224 = ~n197 & n223 ;
  assign n225 = n224 ^ n170 ;
  assign n226 = n225 ^ n197 ;
  assign n227 = n173 & ~n226 ;
  assign n228 = n227 ^ n224 ;
  assign n229 = n228 ^ n197 ;
  assign n230 = x5 & ~n229 ;
  assign n231 = n230 ^ x5 ;
  assign n232 = ~n164 & ~n231 ;
  assign n233 = ~n162 & n232 ;
  assign n234 = ~n36 & n233 ;
  assign n235 = ~x0 & ~x3 ;
  assign n236 = ~x1 & n235 ;
  assign n237 = ~x2 & n236 ;
  assign n238 = ~n234 & n237 ;
  assign y0 = n238 ;
endmodule
