module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n8 = x1 ^ x0 ;
  assign n9 = n8 ^ x2 ;
  assign n10 = n9 ^ x1 ;
  assign n11 = x5 & x6 ;
  assign n12 = n11 ^ x2 ;
  assign n13 = x4 ^ x2 ;
  assign n14 = n12 & n13 ;
  assign n15 = n14 ^ x2 ;
  assign n16 = n15 ^ n9 ;
  assign n17 = n16 ^ x1 ;
  assign n18 = ~x3 & n17 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = n19 ^ n9 ;
  assign n21 = ~n10 & n20 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = x1 & n22 ;
  assign n24 = n23 ^ n8 ;
  assign y0 = n24 ;
endmodule
