module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n18 = ~x0 & ~x11 ;
  assign n19 = x13 ^ x12 ;
  assign n20 = n19 ^ n18 ;
  assign n23 = ~x5 & ~x14 ;
  assign n24 = x1 & x4 ;
  assign n25 = ~x3 & ~x16 ;
  assign n26 = ~x2 & ~x15 ;
  assign n27 = n25 & n26 ;
  assign n28 = n24 & n27 ;
  assign n29 = n23 & n28 ;
  assign n21 = x15 & x16 ;
  assign n22 = x14 & n21 ;
  assign n30 = n29 ^ n22 ;
  assign n31 = ~x13 & n30 ;
  assign n32 = n31 ^ n22 ;
  assign n33 = ~n20 & ~n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n34 ^ n22 ;
  assign n36 = n35 ^ x13 ;
  assign n37 = n18 & n36 ;
  assign y0 = n37 ;
endmodule
