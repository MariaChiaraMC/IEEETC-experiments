module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 ;
  assign n13 = x5 & x11 ;
  assign n14 = ~x0 & ~n13 ;
  assign n15 = x1 & x6 ;
  assign n16 = ~n14 & n15 ;
  assign n17 = ~x0 & ~x4 ;
  assign n18 = ~x1 & ~x5 ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = ~x2 & ~x6 ;
  assign n21 = ~x4 & ~x5 ;
  assign n22 = ~n20 & ~n21 ;
  assign n23 = n19 & n22 ;
  assign n24 = ~n16 & ~n23 ;
  assign n25 = x3 & ~n24 ;
  assign n32 = ~x5 & x10 ;
  assign n33 = ~n13 & ~n32 ;
  assign n34 = x1 & ~n33 ;
  assign n35 = ~n19 & ~n34 ;
  assign n37 = n35 ^ x2 ;
  assign n26 = x11 ^ x10 ;
  assign n27 = x6 & n26 ;
  assign n28 = n27 ^ x10 ;
  assign n29 = n28 ^ x6 ;
  assign n30 = x7 ^ x2 ;
  assign n31 = ~n29 & n30 ;
  assign n38 = n31 ^ x6 ;
  assign n39 = n38 ^ n29 ;
  assign n40 = n39 ^ x7 ;
  assign n41 = n37 & ~n40 ;
  assign n36 = n35 ^ n31 ;
  assign n42 = n41 ^ n36 ;
  assign n43 = n42 ^ x6 ;
  assign n44 = n43 ^ n29 ;
  assign n45 = n44 ^ x7 ;
  assign n46 = x7 & ~n45 ;
  assign n47 = n46 ^ x7 ;
  assign n48 = n47 ^ x7 ;
  assign n49 = n48 ^ x7 ;
  assign n50 = ~n25 & ~n49 ;
  assign n51 = x8 & ~n50 ;
  assign n52 = x2 & ~x7 ;
  assign n53 = x3 & ~x6 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = n54 ^ x4 ;
  assign n56 = x2 & x3 ;
  assign n57 = ~x6 & ~x7 ;
  assign n58 = ~n56 & ~n57 ;
  assign n59 = n58 ^ n54 ;
  assign n60 = n59 ^ n58 ;
  assign n61 = n60 ^ n55 ;
  assign n62 = n32 ^ x0 ;
  assign n63 = ~n32 & n62 ;
  assign n64 = n63 ^ n58 ;
  assign n65 = n64 ^ n32 ;
  assign n66 = ~n61 & n65 ;
  assign n67 = n66 ^ n63 ;
  assign n68 = n67 ^ n32 ;
  assign n69 = n55 & ~n68 ;
  assign n70 = n69 ^ n54 ;
  assign n71 = x9 & ~n70 ;
  assign n72 = ~x9 & ~n56 ;
  assign n73 = ~x0 & n33 ;
  assign n74 = ~n58 & ~n73 ;
  assign n75 = ~n72 & n74 ;
  assign n76 = ~n71 & ~n75 ;
  assign n77 = x1 & ~n76 ;
  assign n78 = x10 ^ x7 ;
  assign n79 = n78 ^ x10 ;
  assign n80 = n26 & n79 ;
  assign n81 = n80 ^ x10 ;
  assign n82 = x3 & n81 ;
  assign n83 = ~n77 & ~n82 ;
  assign n84 = ~n51 & n83 ;
  assign n85 = ~n52 & ~n56 ;
  assign n86 = n28 & ~n85 ;
  assign n87 = n86 ^ x9 ;
  assign n88 = n86 ^ n56 ;
  assign n89 = n88 ^ n56 ;
  assign n90 = ~x0 & x4 ;
  assign n91 = ~x2 & x6 ;
  assign n92 = ~x3 & x7 ;
  assign n93 = ~n91 & ~n92 ;
  assign n94 = ~n90 & n93 ;
  assign n95 = ~x5 & n94 ;
  assign n96 = ~x8 & ~n95 ;
  assign n97 = n96 ^ n56 ;
  assign n98 = ~n89 & n97 ;
  assign n99 = n98 ^ n56 ;
  assign n100 = n87 & n99 ;
  assign n101 = n100 ^ x9 ;
  assign n102 = n84 & ~n101 ;
  assign y0 = ~n102 ;
endmodule
