module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 ;
  assign n12 = x1 & x5 ;
  assign n13 = ~x10 & n12 ;
  assign n14 = x0 & n13 ;
  assign n15 = ~x6 & ~x8 ;
  assign n17 = x2 & x3 ;
  assign n16 = ~x7 & x9 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = x7 & ~x9 ;
  assign n21 = x4 & n20 ;
  assign n22 = n21 ^ n16 ;
  assign n23 = n19 & n22 ;
  assign n24 = n23 ^ n16 ;
  assign n25 = n15 & n24 ;
  assign n26 = n14 & n25 ;
  assign y0 = n26 ;
endmodule
