module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 ;
  assign n22 = ~x1 & ~x3 ;
  assign n23 = n22 ^ x3 ;
  assign n24 = ~x2 & n23 ;
  assign n25 = n24 ^ x3 ;
  assign n26 = ~x0 & ~x3 ;
  assign n27 = ~x2 & n26 ;
  assign n28 = n27 ^ x1 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ x4 ;
  assign n31 = x5 ^ x0 ;
  assign n32 = x5 & n31 ;
  assign n33 = n32 ^ n27 ;
  assign n34 = n33 ^ x5 ;
  assign n35 = n30 & n34 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ x5 ;
  assign n38 = ~x4 & n37 ;
  assign n39 = ~n25 & n38 ;
  assign n40 = ~x19 & ~x20 ;
  assign n41 = n40 ^ x18 ;
  assign n42 = n41 ^ x18 ;
  assign n43 = x3 & ~x5 ;
  assign n44 = x4 & n43 ;
  assign n45 = x5 ^ x2 ;
  assign n48 = ~x6 & ~x7 ;
  assign n49 = ~x8 & n48 ;
  assign n50 = x10 & ~x11 ;
  assign n51 = n49 & n50 ;
  assign n52 = ~x10 & x11 ;
  assign n53 = x8 & n48 ;
  assign n54 = n52 & n53 ;
  assign n55 = n48 ^ x10 ;
  assign n56 = ~x8 & n55 ;
  assign n57 = n56 ^ x10 ;
  assign n58 = ~x11 & n57 ;
  assign n59 = ~n54 & ~n58 ;
  assign n60 = x9 & ~n59 ;
  assign n61 = ~n51 & ~n60 ;
  assign n62 = n61 ^ x0 ;
  assign n63 = n62 ^ x0 ;
  assign n46 = x3 ^ x0 ;
  assign n47 = n46 ^ x0 ;
  assign n64 = n63 ^ n47 ;
  assign n65 = ~x12 & ~x13 ;
  assign n66 = n65 ^ x0 ;
  assign n67 = n66 ^ x0 ;
  assign n68 = n67 ^ n63 ;
  assign n69 = ~n63 & ~n68 ;
  assign n70 = n69 ^ n63 ;
  assign n71 = n64 & ~n70 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = n72 ^ x0 ;
  assign n74 = n73 ^ n63 ;
  assign n75 = ~x4 & n74 ;
  assign n76 = n75 ^ x0 ;
  assign n77 = n76 ^ x5 ;
  assign n78 = n77 ^ n76 ;
  assign n79 = ~x3 & x13 ;
  assign n80 = ~n26 & ~n79 ;
  assign n81 = n80 ^ n76 ;
  assign n82 = n78 & ~n81 ;
  assign n83 = n82 ^ n76 ;
  assign n84 = n45 & n83 ;
  assign n85 = n84 ^ x2 ;
  assign n86 = ~n44 & ~n85 ;
  assign n87 = x1 & ~n86 ;
  assign n88 = x2 & ~x3 ;
  assign n89 = ~x17 & n49 ;
  assign n90 = x16 & n52 ;
  assign n91 = n89 & n90 ;
  assign n92 = x15 ^ x12 ;
  assign n93 = x13 & n92 ;
  assign n94 = n93 ^ x12 ;
  assign n95 = n91 & ~n94 ;
  assign n96 = n88 & ~n95 ;
  assign n97 = ~x1 & x3 ;
  assign n98 = ~x12 & n79 ;
  assign n99 = ~n97 & ~n98 ;
  assign n100 = ~x2 & ~n99 ;
  assign n101 = ~n96 & ~n100 ;
  assign n102 = ~x8 & ~x11 ;
  assign n103 = n79 & n102 ;
  assign n104 = ~x10 & n103 ;
  assign n105 = x2 & n58 ;
  assign n106 = ~x1 & n53 ;
  assign n107 = n52 & n106 ;
  assign n108 = ~n105 & ~n107 ;
  assign n109 = ~x0 & ~x4 ;
  assign n110 = ~x13 & n109 ;
  assign n111 = ~n108 & n110 ;
  assign n112 = ~x1 & ~x8 ;
  assign n113 = ~x10 & ~n112 ;
  assign n114 = ~x3 & x11 ;
  assign n115 = ~n113 & n114 ;
  assign n116 = ~n111 & ~n115 ;
  assign n117 = ~x12 & ~n116 ;
  assign n118 = ~n88 & ~n117 ;
  assign n119 = ~n104 & n118 ;
  assign n120 = x9 & ~n119 ;
  assign n121 = ~x3 & ~x4 ;
  assign n122 = ~x12 & n48 ;
  assign n123 = ~x13 & ~n122 ;
  assign n124 = n109 & ~n123 ;
  assign n125 = ~x9 & n52 ;
  assign n126 = ~x13 & n50 ;
  assign n127 = ~n125 & ~n126 ;
  assign n128 = x2 & ~x8 ;
  assign n129 = ~n127 & n128 ;
  assign n130 = n124 & n129 ;
  assign n131 = ~n121 & ~n130 ;
  assign n132 = ~n120 & n131 ;
  assign n133 = n101 & n132 ;
  assign n134 = x5 & ~n133 ;
  assign n135 = ~x2 & ~x4 ;
  assign n136 = x9 & n65 ;
  assign n137 = n58 & n97 ;
  assign n138 = n48 & n102 ;
  assign n139 = ~n54 & ~n138 ;
  assign n140 = ~x0 & ~x5 ;
  assign n141 = ~n139 & n140 ;
  assign n142 = ~n137 & ~n141 ;
  assign n143 = n136 & ~n142 ;
  assign n144 = ~x0 & ~x1 ;
  assign n145 = n51 & n144 ;
  assign n146 = n65 & n145 ;
  assign n147 = ~n26 & ~n146 ;
  assign n148 = ~n143 & n147 ;
  assign n149 = n135 & ~n148 ;
  assign n154 = n43 ^ x4 ;
  assign n151 = n106 & n136 ;
  assign n152 = n52 & n151 ;
  assign n150 = n43 ^ x0 ;
  assign n153 = n152 ^ n150 ;
  assign n155 = n154 ^ n153 ;
  assign n156 = n155 ^ n153 ;
  assign n157 = n156 ^ x4 ;
  assign n158 = n157 ^ n150 ;
  assign n161 = n22 ^ x2 ;
  assign n162 = n161 ^ n22 ;
  assign n159 = n22 ^ x5 ;
  assign n160 = n159 ^ n22 ;
  assign n163 = n162 ^ n160 ;
  assign n164 = x13 & n125 ;
  assign n165 = ~x8 & n164 ;
  assign n166 = n49 & n65 ;
  assign n167 = x11 ^ x10 ;
  assign n168 = n166 & n167 ;
  assign n169 = ~n165 & ~n168 ;
  assign n170 = ~n136 & n169 ;
  assign n171 = n170 ^ n22 ;
  assign n172 = n171 ^ n22 ;
  assign n173 = n172 ^ n162 ;
  assign n174 = ~n162 & n173 ;
  assign n175 = n174 ^ n162 ;
  assign n176 = ~n163 & ~n175 ;
  assign n177 = n176 ^ n174 ;
  assign n178 = n177 ^ n22 ;
  assign n179 = n178 ^ n162 ;
  assign n180 = ~x4 & ~n179 ;
  assign n181 = n180 ^ n22 ;
  assign n182 = n181 ^ x4 ;
  assign n183 = ~n158 & n182 ;
  assign n184 = n183 ^ n181 ;
  assign n199 = n158 ^ n150 ;
  assign n185 = n112 & n125 ;
  assign n186 = ~x4 & n57 ;
  assign n187 = x9 & ~x11 ;
  assign n188 = x10 & n102 ;
  assign n189 = ~n187 & ~n188 ;
  assign n190 = n65 & ~n189 ;
  assign n191 = n186 & n190 ;
  assign n192 = ~n152 & ~n191 ;
  assign n193 = ~n185 & n192 ;
  assign n194 = n88 & ~n193 ;
  assign n195 = n194 ^ n153 ;
  assign n196 = ~n153 & n195 ;
  assign n197 = n196 ^ n153 ;
  assign n198 = n197 ^ n158 ;
  assign n200 = n199 ^ n198 ;
  assign n201 = n195 ^ x4 ;
  assign n202 = n201 ^ n158 ;
  assign n203 = n202 ^ n199 ;
  assign n204 = ~n202 & n203 ;
  assign n205 = n204 ^ n194 ;
  assign n206 = n205 ^ n199 ;
  assign n207 = ~n200 & n206 ;
  assign n208 = n207 ^ n158 ;
  assign n209 = n208 ^ n199 ;
  assign n210 = n184 & n209 ;
  assign n211 = n210 ^ n207 ;
  assign n212 = n211 ^ n158 ;
  assign n213 = n212 ^ n199 ;
  assign n214 = n213 ^ x0 ;
  assign n215 = ~n149 & ~n214 ;
  assign n216 = ~n134 & n215 ;
  assign n217 = ~n87 & n216 ;
  assign n218 = n217 ^ x18 ;
  assign n219 = n42 & n218 ;
  assign n220 = n219 ^ x18 ;
  assign n221 = x14 & n220 ;
  assign n222 = ~n39 & n221 ;
  assign y0 = ~n222 ;
endmodule
