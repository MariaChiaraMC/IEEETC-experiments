module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n9 = x3 ^ x1 ;
  assign n10 = x3 ^ x2 ;
  assign n11 = n10 ^ x2 ;
  assign n12 = n11 ^ n9 ;
  assign n13 = x5 & x6 ;
  assign n14 = x2 & ~n13 ;
  assign n15 = x4 & ~n14 ;
  assign n16 = x7 ^ x5 ;
  assign n17 = x7 ^ x6 ;
  assign n18 = x6 ^ x2 ;
  assign n19 = n18 ^ x6 ;
  assign n20 = n17 & n19 ;
  assign n21 = n20 ^ x6 ;
  assign n22 = n16 & ~n21 ;
  assign n23 = n22 ^ x5 ;
  assign n24 = ~x4 & ~n23 ;
  assign n25 = n24 ^ n15 ;
  assign n26 = ~n15 & n25 ;
  assign n27 = n26 ^ x2 ;
  assign n28 = n27 ^ n15 ;
  assign n29 = n12 & ~n28 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n30 ^ n15 ;
  assign n32 = ~n9 & ~n31 ;
  assign n33 = ~x0 & n32 ;
  assign y0 = n33 ;
endmodule
