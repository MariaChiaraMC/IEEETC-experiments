// Benchmark "./pla/dc2.pla_dbb_orig_6NonExact" written by ABC on Fri Nov 20 10:18:47 2020

module \./pla/dc2.pla_dbb_orig_6NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = x0;
endmodule


