module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n13 = x8 ^ x0 ;
  assign n14 = ~x2 & x7 ;
  assign n15 = n14 ^ x8 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = ~x1 & ~x2 ;
  assign n18 = ~x3 & x6 ;
  assign n19 = n17 & n18 ;
  assign n20 = n19 ^ n14 ;
  assign n21 = n20 ^ n13 ;
  assign n22 = ~n16 & n21 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = ~x5 & ~x9 ;
  assign n25 = n19 & n24 ;
  assign n26 = n25 ^ n13 ;
  assign n27 = n23 & ~n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = ~n13 & n28 ;
  assign n30 = n29 ^ n22 ;
  assign n31 = n30 ^ n19 ;
  assign y0 = n31 ;
endmodule
