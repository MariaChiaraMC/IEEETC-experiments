module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n9 = x5 & x6 ;
  assign n10 = ~x3 & ~n9 ;
  assign n11 = x2 & ~n10 ;
  assign n14 = x7 ^ x3 ;
  assign n12 = x5 ^ x3 ;
  assign n13 = n12 ^ x3 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = x6 ^ x2 ;
  assign n17 = n14 ^ x3 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = n16 & n18 ;
  assign n20 = n19 ^ x6 ;
  assign n21 = n14 & ~n20 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = ~n15 & ~n22 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n24 ^ x3 ;
  assign n26 = n25 ^ n14 ;
  assign n27 = n26 ^ n13 ;
  assign n28 = ~x4 & n27 ;
  assign n29 = n28 ^ x3 ;
  assign n30 = ~n11 & n29 ;
  assign y0 = n30 ;
endmodule
