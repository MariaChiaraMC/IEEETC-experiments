module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n9 = x4 & ~x6 ;
  assign n10 = ~x5 & ~x7 ;
  assign n11 = ~n9 & n10 ;
  assign n12 = ~x2 & x3 ;
  assign n13 = ~n11 & n12 ;
  assign n14 = ~x4 & ~x5 ;
  assign n15 = ~x2 & ~x7 ;
  assign n16 = n15 ^ x6 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n15 ^ x3 ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = n19 ^ n15 ;
  assign n21 = n14 & n20 ;
  assign n22 = ~n13 & ~n21 ;
  assign n23 = ~x0 & ~x1 ;
  assign n24 = ~n22 & n23 ;
  assign y0 = n24 ;
endmodule
