module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 ;
  assign n9 = x1 ^ x0 ;
  assign n10 = x7 ^ x6 ;
  assign n11 = ~x5 & ~n10 ;
  assign n12 = n11 ^ x6 ;
  assign n13 = x5 & x7 ;
  assign n14 = x4 & ~n13 ;
  assign n15 = ~x2 & n14 ;
  assign n16 = n15 ^ x4 ;
  assign n17 = ~n12 & n16 ;
  assign n18 = ~x0 & n17 ;
  assign n19 = x4 & x5 ;
  assign n20 = ~x0 & ~x6 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = ~x2 & n21 ;
  assign n23 = x0 & n22 ;
  assign n24 = x5 & ~x6 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = x7 ^ x4 ;
  assign n27 = n26 ^ x4 ;
  assign n28 = n27 ^ n23 ;
  assign n29 = n28 ^ n22 ;
  assign n30 = n25 & n29 ;
  assign n31 = n30 ^ x4 ;
  assign n32 = n23 & n31 ;
  assign n33 = n32 ^ n23 ;
  assign n34 = n33 ^ n22 ;
  assign n35 = ~n18 & ~n34 ;
  assign n36 = ~x3 & ~n35 ;
  assign n37 = n36 ^ n9 ;
  assign n38 = n37 ^ x1 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = x3 ^ x2 ;
  assign n41 = ~x5 & x7 ;
  assign n42 = n41 ^ x6 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = n43 ^ x4 ;
  assign n45 = x5 ^ x1 ;
  assign n46 = ~x5 & n45 ;
  assign n47 = n46 ^ n41 ;
  assign n48 = n47 ^ x5 ;
  assign n49 = n44 & ~n48 ;
  assign n50 = n49 ^ n46 ;
  assign n51 = n50 ^ x5 ;
  assign n52 = ~x4 & ~n51 ;
  assign n53 = n52 ^ x3 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = n54 ^ n40 ;
  assign n56 = ~x1 & x7 ;
  assign n57 = x6 ^ x5 ;
  assign n58 = x4 & ~n57 ;
  assign n59 = n58 ^ x5 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = n56 & n60 ;
  assign n62 = n61 ^ n52 ;
  assign n63 = n62 ^ n56 ;
  assign n64 = n55 & n63 ;
  assign n65 = n64 ^ n61 ;
  assign n66 = n65 ^ n56 ;
  assign n67 = n40 & n66 ;
  assign n68 = n67 ^ n37 ;
  assign n69 = n68 ^ n9 ;
  assign n70 = n39 & ~n69 ;
  assign n71 = n70 ^ n67 ;
  assign n75 = ~x4 & x6 ;
  assign n72 = ~x4 & x5 ;
  assign n73 = ~x2 & ~n72 ;
  assign n74 = ~n14 & n73 ;
  assign n76 = n75 ^ n74 ;
  assign n77 = n76 ^ n74 ;
  assign n78 = ~x2 & ~x7 ;
  assign n79 = n78 ^ n74 ;
  assign n80 = n77 & ~n79 ;
  assign n81 = n80 ^ n74 ;
  assign n82 = x3 & n81 ;
  assign n83 = ~n67 & ~n82 ;
  assign n84 = n83 ^ n9 ;
  assign n85 = ~n71 & n84 ;
  assign n86 = n85 ^ n83 ;
  assign n87 = n9 & n86 ;
  assign n88 = n87 ^ n70 ;
  assign n89 = n88 ^ x0 ;
  assign n90 = n89 ^ n67 ;
  assign y0 = n90 ;
endmodule
