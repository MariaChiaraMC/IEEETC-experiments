module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 ;
  assign n16 = ~x1 & x3 ;
  assign n17 = ~x12 & n16 ;
  assign n18 = ~x14 & n17 ;
  assign n19 = ~x7 & ~x9 ;
  assign n20 = n19 ^ x10 ;
  assign n21 = x2 & ~x6 ;
  assign n22 = x5 & n21 ;
  assign n23 = ~x0 & x4 ;
  assign n24 = n22 & n23 ;
  assign n25 = n24 ^ n19 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n26 ^ n20 ;
  assign n28 = x7 & x9 ;
  assign n29 = x8 & ~n28 ;
  assign n30 = ~x4 & ~x5 ;
  assign n31 = x0 & n30 ;
  assign n32 = x6 & n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n29 & n33 ;
  assign n35 = n34 ^ n24 ;
  assign n36 = n35 ^ n29 ;
  assign n37 = n27 & n36 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = n38 ^ n29 ;
  assign n40 = ~n20 & n39 ;
  assign n41 = n18 & n40 ;
  assign n42 = x10 ^ x2 ;
  assign n43 = x10 ^ x5 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = x6 ^ x3 ;
  assign n46 = ~x5 & n45 ;
  assign n47 = n46 ^ x6 ;
  assign n48 = n44 & n47 ;
  assign n49 = n48 ^ n46 ;
  assign n50 = n49 ^ x6 ;
  assign n51 = n50 ^ x5 ;
  assign n52 = ~n42 & ~n51 ;
  assign n53 = n52 ^ x2 ;
  assign n54 = ~x8 & n53 ;
  assign n64 = x3 ^ x1 ;
  assign n65 = x12 ^ x3 ;
  assign n66 = ~n64 & n65 ;
  assign n68 = ~x7 & x14 ;
  assign n67 = x10 & n21 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = n68 ^ x12 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = n71 ^ n66 ;
  assign n73 = n69 & n72 ;
  assign n74 = n73 ^ n67 ;
  assign n75 = n66 & n74 ;
  assign n55 = ~x1 & ~x3 ;
  assign n56 = x2 & n55 ;
  assign n57 = ~x14 & ~n56 ;
  assign n58 = n32 & n57 ;
  assign n59 = x1 & ~x12 ;
  assign n60 = x7 & ~n59 ;
  assign n61 = n58 & n60 ;
  assign n76 = n75 ^ n61 ;
  assign n77 = n76 ^ n61 ;
  assign n62 = n61 ^ n23 ;
  assign n63 = n62 ^ n61 ;
  assign n78 = n77 ^ n63 ;
  assign n79 = n61 ^ x5 ;
  assign n80 = n79 ^ n61 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n77 & n81 ;
  assign n83 = n82 ^ n77 ;
  assign n84 = n78 & n83 ;
  assign n85 = n84 ^ n82 ;
  assign n86 = n85 ^ n61 ;
  assign n87 = n86 ^ n77 ;
  assign n88 = x9 & n87 ;
  assign n89 = n88 ^ n61 ;
  assign n90 = n54 & n89 ;
  assign n91 = ~n41 & ~n90 ;
  assign n92 = ~x13 & ~n91 ;
  assign n93 = ~x0 & ~x10 ;
  assign n94 = ~x2 & n30 ;
  assign n95 = ~x6 & ~x8 ;
  assign n96 = n55 & n95 ;
  assign n97 = n94 & n96 ;
  assign n98 = ~x9 & ~x12 ;
  assign n99 = x13 & n98 ;
  assign n100 = n97 & n99 ;
  assign n101 = n93 & n100 ;
  assign n102 = n68 & n101 ;
  assign n103 = ~n92 & ~n102 ;
  assign n104 = ~x11 & ~n103 ;
  assign y0 = n104 ;
endmodule
