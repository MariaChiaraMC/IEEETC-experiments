module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 ;
  assign n16 = ~x0 & ~x11 ;
  assign n17 = x7 & ~x14 ;
  assign n18 = x4 & n17 ;
  assign n26 = x8 ^ x1 ;
  assign n27 = n26 ^ x10 ;
  assign n28 = x10 ^ x1 ;
  assign n29 = x10 ^ x9 ;
  assign n30 = n29 ^ x10 ;
  assign n31 = ~x10 & ~n30 ;
  assign n32 = n31 ^ x10 ;
  assign n33 = n28 & ~n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n34 ^ x10 ;
  assign n36 = n35 ^ n29 ;
  assign n37 = n27 & ~n36 ;
  assign n19 = ~x6 & ~x8 ;
  assign n20 = ~x9 & x10 ;
  assign n21 = ~x1 & ~x3 ;
  assign n22 = n20 & n21 ;
  assign n23 = n19 & n22 ;
  assign n38 = n37 ^ n23 ;
  assign n39 = n38 ^ n23 ;
  assign n24 = n23 ^ x6 ;
  assign n25 = n24 ^ n23 ;
  assign n40 = n39 ^ n25 ;
  assign n41 = n23 ^ x3 ;
  assign n42 = n41 ^ n23 ;
  assign n43 = n42 ^ n39 ;
  assign n44 = n39 & n43 ;
  assign n45 = n44 ^ n39 ;
  assign n46 = n40 & n45 ;
  assign n47 = n46 ^ n44 ;
  assign n48 = n47 ^ n23 ;
  assign n49 = n48 ^ n39 ;
  assign n50 = ~x5 & n49 ;
  assign n51 = n50 ^ n23 ;
  assign n52 = n18 & n51 ;
  assign n53 = ~x7 & ~x8 ;
  assign n54 = ~x4 & ~x5 ;
  assign n55 = n53 & n54 ;
  assign n56 = ~x6 & ~x9 ;
  assign n57 = ~x10 & x14 ;
  assign n58 = n56 & n57 ;
  assign n59 = n21 & n58 ;
  assign n60 = n55 & n59 ;
  assign n61 = ~n52 & ~n60 ;
  assign n62 = ~x2 & ~n61 ;
  assign n63 = x9 & n53 ;
  assign n64 = x2 & x10 ;
  assign n65 = ~x14 & n64 ;
  assign n66 = x4 & x5 ;
  assign n67 = ~x1 & x3 ;
  assign n68 = x6 & n67 ;
  assign n69 = n66 & n68 ;
  assign n70 = n65 & n69 ;
  assign n71 = n63 & n70 ;
  assign n72 = ~n62 & ~n71 ;
  assign n73 = ~x12 & ~x13 ;
  assign n74 = ~n72 & n73 ;
  assign n75 = n16 & n74 ;
  assign y0 = n75 ;
endmodule
