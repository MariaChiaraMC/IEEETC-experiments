module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 ;
  assign n41 = ~x13 & ~x14 ;
  assign n78 = x3 & x4 ;
  assign n79 = n41 & n78 ;
  assign n23 = x4 & ~x14 ;
  assign n24 = ~x3 & x13 ;
  assign n25 = n23 & n24 ;
  assign n18 = x5 ^ x4 ;
  assign n19 = x14 ^ x5 ;
  assign n20 = n18 & n19 ;
  assign n21 = n20 ^ x4 ;
  assign n16 = x3 & x13 ;
  assign n27 = ~x3 & ~x13 ;
  assign n75 = ~n16 & ~n27 ;
  assign n76 = ~n21 & ~n75 ;
  assign n77 = ~n25 & ~n76 ;
  assign n80 = n79 ^ n77 ;
  assign n81 = x2 & ~n80 ;
  assign n82 = n81 ^ n79 ;
  assign n17 = ~x6 & n16 ;
  assign n22 = n17 & ~n21 ;
  assign n26 = ~x4 & x14 ;
  assign n28 = n26 & n27 ;
  assign n29 = ~n25 & ~n28 ;
  assign n30 = x14 & n27 ;
  assign n31 = ~x5 & n30 ;
  assign n32 = n29 & ~n31 ;
  assign n33 = ~n22 & n32 ;
  assign n34 = ~x1 & ~x2 ;
  assign n35 = x0 & x6 ;
  assign n36 = n34 & ~n35 ;
  assign n37 = ~n33 & n36 ;
  assign n38 = x11 & n37 ;
  assign n39 = x13 & x14 ;
  assign n40 = x6 & ~n39 ;
  assign n42 = x13 ^ x4 ;
  assign n43 = ~x2 & ~x3 ;
  assign n44 = n43 ^ x4 ;
  assign n45 = x4 & n44 ;
  assign n46 = n45 ^ x4 ;
  assign n47 = ~n18 & n46 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = n48 ^ x4 ;
  assign n50 = n49 ^ n43 ;
  assign n51 = n42 & n50 ;
  assign n52 = n51 ^ n43 ;
  assign n53 = ~x1 & n52 ;
  assign n54 = ~n41 & ~n53 ;
  assign n55 = ~x0 & ~n54 ;
  assign n56 = n55 ^ n40 ;
  assign n57 = x8 & x9 ;
  assign n58 = ~x7 & ~x11 ;
  assign n59 = ~n57 & n58 ;
  assign n60 = n59 ^ n41 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = n59 ^ x11 ;
  assign n63 = ~n61 & n62 ;
  assign n64 = n63 ^ n59 ;
  assign n65 = n64 ^ n40 ;
  assign n66 = ~n56 & n65 ;
  assign n67 = n66 ^ n63 ;
  assign n68 = n67 ^ n59 ;
  assign n69 = n68 ^ n55 ;
  assign n70 = n40 & ~n69 ;
  assign n71 = n70 ^ n40 ;
  assign n72 = ~n38 & ~n71 ;
  assign n83 = n82 ^ n72 ;
  assign n84 = n83 ^ n72 ;
  assign n73 = n72 ^ x1 ;
  assign n74 = n73 ^ n72 ;
  assign n85 = n84 ^ n74 ;
  assign n86 = ~x6 & x11 ;
  assign n87 = n86 ^ n72 ;
  assign n88 = n87 ^ n72 ;
  assign n89 = n88 ^ n84 ;
  assign n90 = n84 & n89 ;
  assign n91 = n90 ^ n84 ;
  assign n92 = ~n85 & n91 ;
  assign n93 = n92 ^ n90 ;
  assign n94 = n93 ^ n72 ;
  assign n95 = n94 ^ n84 ;
  assign n96 = x12 & ~n95 ;
  assign n97 = n96 ^ n72 ;
  assign n98 = ~x10 & ~n97 ;
  assign n99 = x10 & ~x11 ;
  assign n102 = ~x2 & n79 ;
  assign n100 = n26 & ~n75 ;
  assign n101 = ~n25 & ~n100 ;
  assign n103 = n102 ^ n101 ;
  assign n104 = n101 ^ x12 ;
  assign n105 = n104 ^ x2 ;
  assign n106 = n105 ^ n101 ;
  assign n107 = n106 ^ n99 ;
  assign n108 = ~n103 & n107 ;
  assign n109 = n108 ^ n102 ;
  assign n110 = n99 & n109 ;
  assign n111 = ~n98 & ~n110 ;
  assign y0 = ~n111 ;
endmodule
