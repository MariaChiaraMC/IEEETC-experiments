module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 ;
  assign n13 = x9 ^ x7 ;
  assign n14 = x2 & x6 ;
  assign n15 = n14 ^ x7 ;
  assign n16 = ~x10 & ~x11 ;
  assign n17 = n16 ^ x7 ;
  assign n18 = ~x7 & ~n17 ;
  assign n19 = n18 ^ x7 ;
  assign n20 = n15 & ~n19 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n21 ^ x7 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = ~n13 & ~n23 ;
  assign n25 = x7 & ~x9 ;
  assign n50 = n25 ^ x5 ;
  assign n26 = x3 ^ x0 ;
  assign n27 = x11 ^ x10 ;
  assign n28 = x10 ^ x3 ;
  assign n29 = n28 ^ x10 ;
  assign n30 = ~n27 & ~n29 ;
  assign n31 = n30 ^ x10 ;
  assign n32 = n26 & n31 ;
  assign n33 = n25 & n32 ;
  assign n34 = ~x7 & x11 ;
  assign n35 = n34 ^ n16 ;
  assign n36 = n35 ^ x9 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = n37 ^ x0 ;
  assign n39 = n34 ^ x3 ;
  assign n40 = x3 & n39 ;
  assign n41 = n40 ^ n35 ;
  assign n42 = n41 ^ x3 ;
  assign n43 = ~n38 & n42 ;
  assign n44 = n43 ^ n40 ;
  assign n45 = n44 ^ x3 ;
  assign n46 = x0 & n45 ;
  assign n47 = n46 ^ n34 ;
  assign n48 = ~n33 & ~n47 ;
  assign n49 = n48 ^ x5 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = n51 ^ x11 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n51 ^ n49 ;
  assign n55 = n54 ^ x5 ;
  assign n56 = n53 & n55 ;
  assign n57 = n56 ^ n49 ;
  assign n58 = x3 & x10 ;
  assign n59 = ~n49 & n58 ;
  assign n60 = n59 ^ x5 ;
  assign n61 = ~n57 & n60 ;
  assign n62 = n61 ^ n59 ;
  assign n63 = x5 & n62 ;
  assign n64 = n63 ^ n56 ;
  assign n65 = n64 ^ n48 ;
  assign n66 = n65 ^ n49 ;
  assign n67 = ~n24 & ~n66 ;
  assign n68 = n67 ^ x7 ;
  assign n69 = n68 ^ x8 ;
  assign n81 = n69 ^ n68 ;
  assign n70 = ~x3 & x9 ;
  assign n71 = x0 & ~n70 ;
  assign n72 = ~x10 & x11 ;
  assign n73 = ~n71 & n72 ;
  assign n74 = x5 & n73 ;
  assign n75 = n74 ^ n69 ;
  assign n76 = n75 ^ n68 ;
  assign n77 = n69 ^ n67 ;
  assign n78 = n77 ^ n74 ;
  assign n79 = n78 ^ n76 ;
  assign n80 = n76 & n79 ;
  assign n82 = n81 ^ n80 ;
  assign n83 = n82 ^ n76 ;
  assign n84 = x9 & n16 ;
  assign n85 = ~x5 & x6 ;
  assign n86 = n84 & n85 ;
  assign n87 = ~x9 & x10 ;
  assign n88 = x5 & n87 ;
  assign n89 = x0 & n88 ;
  assign n90 = ~n86 & ~n89 ;
  assign n91 = n90 ^ n68 ;
  assign n92 = n80 ^ n76 ;
  assign n93 = n91 & n92 ;
  assign n94 = n93 ^ n68 ;
  assign n95 = ~n83 & n94 ;
  assign n96 = n95 ^ n68 ;
  assign n97 = n96 ^ x7 ;
  assign n98 = n97 ^ n68 ;
  assign n99 = ~x4 & ~n98 ;
  assign n100 = ~x2 & x4 ;
  assign n101 = n100 ^ n72 ;
  assign n102 = ~x8 & n101 ;
  assign n103 = n102 ^ n72 ;
  assign n104 = x9 & n103 ;
  assign n105 = n100 ^ x11 ;
  assign n106 = ~x1 & x9 ;
  assign n107 = x2 & n106 ;
  assign n108 = x8 & ~n107 ;
  assign n109 = n108 ^ n100 ;
  assign n110 = n109 ^ n100 ;
  assign n111 = n110 ^ n105 ;
  assign n112 = x10 ^ x9 ;
  assign n113 = ~n100 & ~n112 ;
  assign n114 = n113 ^ x9 ;
  assign n115 = n111 & ~n114 ;
  assign n116 = n115 ^ n113 ;
  assign n117 = n116 ^ x9 ;
  assign n118 = n117 ^ n100 ;
  assign n119 = n105 & n118 ;
  assign n120 = n119 ^ x11 ;
  assign n121 = ~n104 & ~n120 ;
  assign n122 = ~x7 & ~n121 ;
  assign n123 = ~x8 & n100 ;
  assign n124 = ~n25 & ~n87 ;
  assign n125 = n123 & ~n124 ;
  assign n126 = ~n122 & ~n125 ;
  assign n127 = x5 & ~n126 ;
  assign n128 = ~n99 & ~n127 ;
  assign y0 = ~n128 ;
endmodule
