// Benchmark "./pla/opa.pla_dbb_orig_67NonExact" written by ABC on Fri Nov 20 10:27:44 2020

module \./pla/opa.pla_dbb_orig_67NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = 1'b1;
endmodule


