module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 ;
  assign n33 = x9 & x10 ;
  assign n34 = x5 & ~n33 ;
  assign n35 = x7 & ~n34 ;
  assign n36 = x14 & ~x15 ;
  assign n37 = ~x11 & n36 ;
  assign n38 = ~x8 & n37 ;
  assign n39 = ~n35 & n38 ;
  assign n40 = ~x4 & x5 ;
  assign n41 = ~x7 & ~n40 ;
  assign n42 = ~x6 & ~n41 ;
  assign n43 = ~x9 & ~x10 ;
  assign n44 = ~x12 & ~x13 ;
  assign n45 = ~n43 & n44 ;
  assign n46 = ~x0 & n45 ;
  assign n47 = ~n42 & n46 ;
  assign n48 = n39 & n47 ;
  assign n19 = x6 ^ x4 ;
  assign n20 = n19 ^ x6 ;
  assign n17 = x6 ^ x5 ;
  assign n18 = n17 ^ x6 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = x7 ^ x6 ;
  assign n23 = n22 ^ x6 ;
  assign n24 = n23 ^ n20 ;
  assign n25 = n20 & n24 ;
  assign n26 = n25 ^ n20 ;
  assign n27 = n21 & n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n28 ^ x6 ;
  assign n30 = n29 ^ n20 ;
  assign n31 = ~x0 & n30 ;
  assign n32 = n31 ^ x6 ;
  assign n49 = n48 ^ n32 ;
  assign n50 = x1 & n49 ;
  assign n51 = n50 ^ n32 ;
  assign y0 = n51 ;
endmodule
