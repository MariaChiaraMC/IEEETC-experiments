module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n11 = ~x3 & ~x6 ;
  assign n12 = ~x2 & n11 ;
  assign n13 = ~x0 & n12 ;
  assign n14 = ~x4 & ~n13 ;
  assign n15 = ~x2 & x8 ;
  assign n16 = ~x0 & ~n15 ;
  assign n17 = ~n12 & ~n16 ;
  assign n18 = x9 ^ x8 ;
  assign n19 = x7 & ~n18 ;
  assign n20 = ~n17 & ~n19 ;
  assign n21 = x3 ^ x2 ;
  assign n22 = x6 ^ x2 ;
  assign n23 = n21 & n22 ;
  assign n24 = n23 ^ x2 ;
  assign n25 = ~x1 & ~n24 ;
  assign n26 = ~x5 & n25 ;
  assign n27 = n20 & n26 ;
  assign n28 = n14 & n27 ;
  assign y0 = n28 ;
endmodule
