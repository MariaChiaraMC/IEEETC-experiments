module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n15 = ~x0 & x2 ;
  assign n16 = x1 & x6 ;
  assign n17 = x4 & n16 ;
  assign n18 = x5 & n17 ;
  assign n26 = x6 ^ x1 ;
  assign n27 = ~x5 & n26 ;
  assign n28 = ~x4 & n27 ;
  assign n29 = ~x3 & ~n28 ;
  assign n19 = x3 & ~x12 ;
  assign n20 = ~x9 & ~x11 ;
  assign n21 = x8 & n20 ;
  assign n22 = n19 & n21 ;
  assign n23 = ~x7 & ~x13 ;
  assign n24 = ~x10 & n23 ;
  assign n25 = n22 & n24 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = n18 & n30 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = n15 & n32 ;
  assign y0 = n33 ;
endmodule
