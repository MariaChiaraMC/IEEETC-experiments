module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 ;
  assign n9 = ~x3 & ~x4 ;
  assign n10 = n9 ^ x2 ;
  assign n11 = ~x6 & ~x7 ;
  assign n12 = x5 & ~n11 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = x6 & x7 ;
  assign n16 = ~x3 & ~x5 ;
  assign n17 = ~n15 & n16 ;
  assign n18 = n17 ^ n12 ;
  assign n19 = ~n14 & n18 ;
  assign n20 = n19 ^ n12 ;
  assign n21 = ~n10 & ~n20 ;
  assign n22 = ~x1 & n21 ;
  assign y0 = ~n22 ;
endmodule
