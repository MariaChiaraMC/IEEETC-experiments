module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 ;
  assign n8 = ~x2 & ~x4 ;
  assign n11 = ~x3 & ~x6 ;
  assign n20 = n8 & ~n11 ;
  assign n21 = x4 ^ x3 ;
  assign n22 = x5 ^ x3 ;
  assign n23 = x1 & x6 ;
  assign n24 = n23 ^ x3 ;
  assign n25 = x3 & ~n24 ;
  assign n26 = n25 ^ x3 ;
  assign n27 = ~n22 & n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n28 ^ x3 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = n21 & ~n30 ;
  assign n32 = ~n20 & ~n31 ;
  assign n9 = x4 ^ x1 ;
  assign n10 = n9 ^ n8 ;
  assign n12 = n11 ^ x6 ;
  assign n13 = x4 & n12 ;
  assign n14 = n13 ^ n11 ;
  assign n15 = ~n10 & n14 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = n16 ^ n11 ;
  assign n18 = n17 ^ x4 ;
  assign n19 = ~n8 & n18 ;
  assign n33 = n32 ^ n19 ;
  assign n34 = x1 & ~x6 ;
  assign n35 = x3 & ~n34 ;
  assign n36 = n35 ^ n19 ;
  assign n37 = n19 ^ x5 ;
  assign n38 = ~n19 & n37 ;
  assign n39 = n38 ^ n19 ;
  assign n40 = n36 & ~n39 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n41 ^ n19 ;
  assign n43 = n42 ^ x5 ;
  assign n44 = ~n33 & n43 ;
  assign n45 = n44 ^ n32 ;
  assign n46 = ~x0 & ~n45 ;
  assign y0 = n46 ;
endmodule
