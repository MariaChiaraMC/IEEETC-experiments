module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 ;
  assign n9 = x2 & ~x3 ;
  assign n10 = ~x4 & ~x5 ;
  assign n11 = x7 & n10 ;
  assign n12 = ~x6 & n11 ;
  assign n13 = x5 & x6 ;
  assign n14 = x4 & ~x7 ;
  assign n15 = n13 & n14 ;
  assign n16 = ~n12 & ~n15 ;
  assign n17 = n9 & ~n16 ;
  assign n18 = ~x2 & x4 ;
  assign n19 = x3 & ~x5 ;
  assign n20 = x6 & ~x7 ;
  assign n21 = n19 & n20 ;
  assign n22 = n18 & n21 ;
  assign n23 = ~n17 & ~n22 ;
  assign n24 = ~x0 & ~n23 ;
  assign n25 = x4 & ~x5 ;
  assign n26 = ~x3 & n25 ;
  assign n27 = x0 & ~x2 ;
  assign n28 = n26 & n27 ;
  assign n29 = n20 & n28 ;
  assign n30 = x0 & x2 ;
  assign n31 = n12 & n30 ;
  assign n32 = ~x0 & x5 ;
  assign n33 = ~x6 & n32 ;
  assign n34 = ~x3 & n33 ;
  assign n35 = n18 & n34 ;
  assign n36 = x6 ^ x4 ;
  assign n43 = x2 ^ x0 ;
  assign n44 = n43 ^ x2 ;
  assign n45 = n43 & ~n44 ;
  assign n37 = x5 ^ x0 ;
  assign n38 = n37 ^ x6 ;
  assign n39 = x6 ^ x0 ;
  assign n40 = n39 ^ x2 ;
  assign n41 = n38 & n40 ;
  assign n48 = n45 ^ n41 ;
  assign n42 = n41 ^ n36 ;
  assign n46 = n45 ^ n43 ;
  assign n47 = ~n42 & n46 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = ~n36 & n49 ;
  assign n51 = n50 ^ n41 ;
  assign n52 = n51 ^ n45 ;
  assign n53 = n52 ^ n47 ;
  assign n54 = n53 ^ x3 ;
  assign n55 = n54 ^ n53 ;
  assign n56 = x4 & x6 ;
  assign n57 = x2 & ~n56 ;
  assign n58 = ~x5 & n57 ;
  assign n59 = n13 & n18 ;
  assign n60 = ~n58 & ~n59 ;
  assign n61 = x0 & ~n60 ;
  assign n62 = n61 ^ n53 ;
  assign n63 = ~n55 & n62 ;
  assign n64 = n63 ^ n53 ;
  assign n65 = ~n35 & ~n64 ;
  assign n66 = n65 ^ x7 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = ~x3 & n56 ;
  assign n69 = ~x2 & ~n37 ;
  assign n70 = n69 ^ x0 ;
  assign n71 = n68 & n70 ;
  assign n72 = ~x2 & ~x4 ;
  assign n73 = n33 & n72 ;
  assign n74 = ~n71 & ~n73 ;
  assign n75 = n74 ^ n65 ;
  assign n76 = ~n67 & n75 ;
  assign n77 = n76 ^ n65 ;
  assign n78 = ~n31 & n77 ;
  assign n79 = n78 ^ x1 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = ~n14 & n34 ;
  assign n82 = ~x4 & ~x7 ;
  assign n83 = n19 & n82 ;
  assign n84 = ~x0 & n83 ;
  assign n85 = ~n81 & ~n84 ;
  assign n86 = x4 & n32 ;
  assign n87 = x3 & n86 ;
  assign n88 = x7 & n26 ;
  assign n89 = ~n87 & ~n88 ;
  assign n90 = x7 ^ x6 ;
  assign n91 = ~n89 & ~n90 ;
  assign n92 = n85 & ~n91 ;
  assign n93 = x2 & ~n92 ;
  assign n97 = x3 ^ x2 ;
  assign n94 = x4 ^ x3 ;
  assign n95 = n94 ^ x7 ;
  assign n104 = n97 ^ n95 ;
  assign n96 = n95 ^ x5 ;
  assign n98 = n97 ^ n96 ;
  assign n99 = n97 ^ x4 ;
  assign n100 = n99 ^ x7 ;
  assign n101 = n100 ^ x5 ;
  assign n102 = n101 ^ n98 ;
  assign n103 = ~n98 & ~n102 ;
  assign n105 = n104 ^ n103 ;
  assign n106 = n105 ^ n98 ;
  assign n107 = n97 ^ x7 ;
  assign n108 = n107 ^ n97 ;
  assign n109 = n103 ^ n98 ;
  assign n110 = ~n108 & ~n109 ;
  assign n111 = n110 ^ n97 ;
  assign n112 = ~n106 & n111 ;
  assign n113 = n112 ^ n97 ;
  assign n114 = n113 ^ n97 ;
  assign n115 = x6 & n114 ;
  assign n116 = ~x6 & ~x7 ;
  assign n117 = x5 ^ x3 ;
  assign n118 = x5 ^ x4 ;
  assign n119 = n118 ^ x4 ;
  assign n120 = n72 ^ x4 ;
  assign n121 = n119 & n120 ;
  assign n122 = n121 ^ x4 ;
  assign n123 = ~n117 & n122 ;
  assign n124 = n116 & n123 ;
  assign n125 = ~n115 & ~n124 ;
  assign n126 = n125 ^ x0 ;
  assign n127 = n126 ^ n125 ;
  assign n128 = n127 ^ n93 ;
  assign n129 = x6 & x7 ;
  assign n130 = n72 & n129 ;
  assign n131 = n130 ^ x5 ;
  assign n132 = x5 & n131 ;
  assign n133 = n132 ^ n125 ;
  assign n134 = n133 ^ x5 ;
  assign n135 = n128 & ~n134 ;
  assign n136 = n135 ^ n132 ;
  assign n137 = n136 ^ x5 ;
  assign n138 = ~n93 & n137 ;
  assign n139 = n138 ^ n93 ;
  assign n140 = n139 ^ n78 ;
  assign n141 = n80 & ~n140 ;
  assign n142 = n141 ^ n78 ;
  assign n143 = ~n29 & n142 ;
  assign n144 = ~n24 & n143 ;
  assign y0 = ~n144 ;
endmodule
