module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 ;
  assign n17 = x4 & x13 ;
  assign n18 = ~x4 & ~x13 ;
  assign n19 = ~x0 & n18 ;
  assign n20 = ~n17 & ~n19 ;
  assign n21 = x6 & ~x12 ;
  assign n22 = n21 ^ x5 ;
  assign n23 = x14 & ~x15 ;
  assign n24 = n23 ^ x7 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = ~x14 & x15 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = ~n25 & n27 ;
  assign n29 = n28 ^ n23 ;
  assign n30 = n29 ^ n21 ;
  assign n31 = ~n22 & n30 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = n32 ^ n23 ;
  assign n34 = n33 ^ x5 ;
  assign n35 = n21 & ~n34 ;
  assign n36 = n35 ^ n21 ;
  assign n37 = ~n20 & n36 ;
  assign n63 = x13 ^ x7 ;
  assign n64 = x14 & x15 ;
  assign n65 = n64 ^ x13 ;
  assign n66 = n65 ^ n64 ;
  assign n67 = n66 ^ n63 ;
  assign n68 = ~x14 & ~x15 ;
  assign n69 = n68 ^ x0 ;
  assign n70 = n68 & ~n69 ;
  assign n71 = n70 ^ n64 ;
  assign n72 = n71 ^ n68 ;
  assign n73 = ~n67 & n72 ;
  assign n74 = n73 ^ n70 ;
  assign n75 = n74 ^ n68 ;
  assign n76 = ~n63 & n75 ;
  assign n77 = ~x4 & n76 ;
  assign n78 = ~x7 & n64 ;
  assign n79 = n17 & n78 ;
  assign n80 = ~n77 & ~n79 ;
  assign n38 = x7 & ~x12 ;
  assign n39 = x15 & n38 ;
  assign n40 = ~x15 & ~n38 ;
  assign n41 = x5 & x14 ;
  assign n42 = n17 & n41 ;
  assign n43 = x0 & ~n42 ;
  assign n44 = n40 & ~n43 ;
  assign n45 = ~n39 & ~n44 ;
  assign n46 = n18 & n41 ;
  assign n47 = ~x5 & ~x14 ;
  assign n48 = n17 & n47 ;
  assign n49 = ~n46 & ~n48 ;
  assign n50 = ~n42 & n49 ;
  assign n51 = ~n45 & ~n50 ;
  assign n52 = ~x4 & x13 ;
  assign n53 = x12 & x14 ;
  assign n54 = ~n52 & n53 ;
  assign n55 = n26 & n38 ;
  assign n56 = n18 & n55 ;
  assign n57 = ~n54 & ~n56 ;
  assign n58 = ~x5 & ~n57 ;
  assign n59 = ~x0 & n58 ;
  assign n60 = ~n51 & ~n59 ;
  assign n81 = n80 ^ n60 ;
  assign n82 = n81 ^ n60 ;
  assign n61 = n60 ^ x12 ;
  assign n62 = n61 ^ n60 ;
  assign n83 = n82 ^ n62 ;
  assign n84 = n60 ^ x5 ;
  assign n85 = n84 ^ n60 ;
  assign n86 = n85 ^ n82 ;
  assign n87 = ~n82 & ~n86 ;
  assign n88 = n87 ^ n82 ;
  assign n89 = n83 & ~n88 ;
  assign n90 = n89 ^ n87 ;
  assign n91 = n90 ^ n60 ;
  assign n92 = n91 ^ n82 ;
  assign n93 = x6 & n92 ;
  assign n94 = n93 ^ n60 ;
  assign n95 = ~n37 & n94 ;
  assign n132 = x1 & ~x8 ;
  assign n133 = ~x3 & n132 ;
  assign n96 = n53 ^ x5 ;
  assign n104 = n96 ^ x5 ;
  assign n97 = n96 ^ x15 ;
  assign n98 = n97 ^ n96 ;
  assign n99 = n98 ^ x5 ;
  assign n100 = n96 ^ n38 ;
  assign n101 = n100 ^ n97 ;
  assign n102 = n101 ^ n99 ;
  assign n103 = n99 & ~n102 ;
  assign n105 = n104 ^ n103 ;
  assign n106 = n105 ^ n99 ;
  assign n107 = x14 ^ x5 ;
  assign n108 = n107 ^ x5 ;
  assign n109 = n103 ^ n99 ;
  assign n110 = ~n108 & n109 ;
  assign n111 = n110 ^ x5 ;
  assign n112 = n106 & n111 ;
  assign n113 = n112 ^ x5 ;
  assign n114 = n113 ^ n53 ;
  assign n115 = n114 ^ x5 ;
  assign n116 = ~x6 & n115 ;
  assign n117 = ~n36 & ~n116 ;
  assign n118 = n18 & ~n117 ;
  assign n119 = x13 & n68 ;
  assign n120 = ~n53 & ~n119 ;
  assign n121 = x4 & ~x6 ;
  assign n122 = ~x5 & n121 ;
  assign n123 = ~n38 & n122 ;
  assign n124 = x6 & x7 ;
  assign n125 = n68 & n124 ;
  assign n126 = x5 & ~x12 ;
  assign n127 = n52 & n126 ;
  assign n128 = n125 & n127 ;
  assign n129 = ~n123 & ~n128 ;
  assign n130 = ~n120 & ~n129 ;
  assign n131 = ~n118 & ~n130 ;
  assign n134 = n133 ^ n131 ;
  assign n135 = n134 ^ n131 ;
  assign n136 = n135 ^ x0 ;
  assign n137 = ~x5 & x9 ;
  assign n138 = ~x10 & n137 ;
  assign n139 = n54 & n138 ;
  assign n140 = ~x9 & ~x10 ;
  assign n141 = ~x12 & ~n140 ;
  assign n142 = n40 & ~n49 ;
  assign n143 = ~n141 & n142 ;
  assign n144 = ~n139 & ~n143 ;
  assign n145 = ~x6 & ~n144 ;
  assign n146 = x5 & x6 ;
  assign n147 = x13 & ~n146 ;
  assign n148 = ~x6 & ~x7 ;
  assign n149 = ~n124 & ~n148 ;
  assign n150 = x15 ^ x5 ;
  assign n151 = ~n149 & n150 ;
  assign n152 = n151 ^ x5 ;
  assign n153 = ~n147 & ~n152 ;
  assign n154 = x9 & x11 ;
  assign n155 = x10 & n154 ;
  assign n156 = ~n140 & ~n155 ;
  assign n157 = ~x13 & n68 ;
  assign n158 = x5 & ~x13 ;
  assign n159 = ~n157 & ~n158 ;
  assign n160 = ~n156 & ~n159 ;
  assign n161 = n124 ^ x6 ;
  assign n162 = ~x5 & ~n161 ;
  assign n163 = n162 ^ x6 ;
  assign n164 = x14 & n163 ;
  assign n165 = ~n160 & ~n164 ;
  assign n166 = n153 & n165 ;
  assign n167 = ~x7 & ~x13 ;
  assign n168 = x5 & n23 ;
  assign n169 = n167 & n168 ;
  assign n170 = n155 & n169 ;
  assign n171 = ~x6 & n170 ;
  assign n172 = ~n166 & ~n171 ;
  assign n173 = ~x4 & ~n172 ;
  assign n175 = n68 & n156 ;
  assign n174 = ~x7 & n122 ;
  assign n176 = n175 ^ n174 ;
  assign n177 = x4 & ~x13 ;
  assign n178 = x7 ^ x6 ;
  assign n179 = n158 & n178 ;
  assign n180 = ~n177 & ~n179 ;
  assign n181 = n180 ^ n174 ;
  assign n182 = n181 ^ n180 ;
  assign n183 = n119 & n155 ;
  assign n184 = n183 ^ n180 ;
  assign n185 = n182 & n184 ;
  assign n186 = n185 ^ n180 ;
  assign n187 = n176 & n186 ;
  assign n188 = n187 ^ n175 ;
  assign n189 = ~n173 & ~n188 ;
  assign n190 = ~x12 & ~n189 ;
  assign n191 = n190 ^ n145 ;
  assign n192 = ~n145 & n191 ;
  assign n193 = n192 ^ n131 ;
  assign n194 = n193 ^ n145 ;
  assign n195 = n136 & ~n194 ;
  assign n196 = n195 ^ n192 ;
  assign n197 = n196 ^ n145 ;
  assign n198 = x0 & ~n197 ;
  assign n199 = n198 ^ x0 ;
  assign n200 = n95 & ~n199 ;
  assign n201 = x2 & ~n200 ;
  assign n202 = n26 ^ x13 ;
  assign n203 = n202 ^ n26 ;
  assign n204 = x6 & ~n23 ;
  assign n205 = n204 ^ n26 ;
  assign n206 = n203 & ~n205 ;
  assign n207 = n206 ^ n26 ;
  assign n208 = x4 & n207 ;
  assign n209 = n208 ^ x13 ;
  assign n210 = ~x5 & n209 ;
  assign n228 = x14 & n177 ;
  assign n229 = x15 ^ x4 ;
  assign n230 = ~x14 & ~n229 ;
  assign n231 = n230 ^ x4 ;
  assign n232 = ~n17 & n231 ;
  assign n233 = n232 ^ x5 ;
  assign n234 = n233 ^ n232 ;
  assign n235 = n234 ^ n228 ;
  assign n236 = n18 ^ x15 ;
  assign n237 = x15 & n236 ;
  assign n238 = n237 ^ n232 ;
  assign n239 = n238 ^ x15 ;
  assign n240 = n235 & ~n239 ;
  assign n241 = n240 ^ n237 ;
  assign n242 = n241 ^ x15 ;
  assign n243 = ~n228 & n242 ;
  assign n244 = n243 ^ n228 ;
  assign n211 = ~n46 & ~n47 ;
  assign n212 = ~n42 & n211 ;
  assign n213 = n212 ^ x2 ;
  assign n214 = n212 ^ x15 ;
  assign n215 = n214 ^ x15 ;
  assign n216 = n215 ^ n213 ;
  assign n217 = x0 & n133 ;
  assign n218 = ~x5 & ~n217 ;
  assign n219 = n218 ^ n138 ;
  assign n220 = ~n138 & n219 ;
  assign n221 = n220 ^ x15 ;
  assign n222 = n221 ^ n138 ;
  assign n223 = ~n216 & ~n222 ;
  assign n224 = n223 ^ n220 ;
  assign n225 = n224 ^ n138 ;
  assign n226 = ~n213 & ~n225 ;
  assign n227 = n226 ^ x2 ;
  assign n245 = n244 ^ n227 ;
  assign n246 = n245 ^ n244 ;
  assign n247 = n244 ^ n157 ;
  assign n248 = n247 ^ n244 ;
  assign n249 = ~n246 & ~n248 ;
  assign n250 = n249 ^ n244 ;
  assign n251 = ~x6 & n250 ;
  assign n252 = n251 ^ n244 ;
  assign n253 = ~n210 & ~n252 ;
  assign n256 = n253 ^ n175 ;
  assign n257 = n256 ^ n253 ;
  assign n254 = n253 ^ n217 ;
  assign n255 = n254 ^ n253 ;
  assign n258 = n257 ^ n255 ;
  assign n259 = ~x2 & ~x13 ;
  assign n260 = n259 ^ n253 ;
  assign n261 = n260 ^ n253 ;
  assign n262 = n261 ^ n257 ;
  assign n263 = n257 & n262 ;
  assign n264 = n263 ^ n257 ;
  assign n265 = n258 & n264 ;
  assign n266 = n265 ^ n263 ;
  assign n267 = n266 ^ n253 ;
  assign n268 = n267 ^ n257 ;
  assign n269 = ~x12 & ~n268 ;
  assign n270 = n269 ^ n253 ;
  assign n271 = ~n201 & n270 ;
  assign y0 = ~n271 ;
endmodule
