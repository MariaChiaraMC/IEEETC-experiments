module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 ;
  assign n7 = x3 & x4 ;
  assign n8 = x1 & ~n7 ;
  assign n9 = ~x2 & ~n8 ;
  assign n10 = x3 & x5 ;
  assign n11 = ~n9 & ~n10 ;
  assign n12 = ~x0 & ~n11 ;
  assign n21 = x5 ^ x0 ;
  assign n13 = x5 ^ x1 ;
  assign n14 = n13 ^ x2 ;
  assign n24 = n21 ^ n14 ;
  assign n22 = n21 ^ x5 ;
  assign n23 = n22 ^ n21 ;
  assign n25 = n24 ^ n23 ;
  assign n15 = n14 ^ x4 ;
  assign n16 = n15 ^ x5 ;
  assign n17 = n14 ^ x3 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = ~n16 & n19 ;
  assign n26 = n25 ^ n20 ;
  assign n27 = n26 ^ n16 ;
  assign n28 = n24 ^ n21 ;
  assign n29 = n14 ^ x2 ;
  assign n30 = n29 ^ n21 ;
  assign n31 = n30 ^ n24 ;
  assign n32 = ~n28 & ~n31 ;
  assign n33 = n32 ^ n21 ;
  assign n34 = n31 ^ n25 ;
  assign n35 = n29 ^ n24 ;
  assign n36 = n35 ^ n25 ;
  assign n37 = ~n34 & n36 ;
  assign n38 = n37 ^ n21 ;
  assign n39 = n38 ^ n29 ;
  assign n40 = n39 ^ n25 ;
  assign n41 = ~n33 & ~n40 ;
  assign n42 = n41 ^ n29 ;
  assign n43 = n42 ^ n25 ;
  assign n44 = ~n27 & n43 ;
  assign n45 = n44 ^ n37 ;
  assign n46 = n45 ^ n32 ;
  assign n47 = n46 ^ n20 ;
  assign n48 = n47 ^ n41 ;
  assign n49 = n48 ^ n29 ;
  assign n50 = n49 ^ n24 ;
  assign n51 = n50 ^ n25 ;
  assign n52 = n51 ^ n16 ;
  assign n53 = n52 ^ x5 ;
  assign n54 = n53 ^ n22 ;
  assign n55 = ~n12 & ~n54 ;
  assign y0 = ~n55 ;
endmodule
