module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 ;
  assign n10 = ~x6 & ~x7 ;
  assign n11 = ~x4 & n10 ;
  assign n12 = x1 & n11 ;
  assign n13 = x1 & x7 ;
  assign n14 = x6 & ~x8 ;
  assign n15 = x4 & x5 ;
  assign n16 = n14 & n15 ;
  assign n17 = n13 & n16 ;
  assign n18 = ~n12 & ~n17 ;
  assign n21 = ~x5 & x7 ;
  assign n19 = ~x4 & x6 ;
  assign n20 = ~x1 & n19 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = ~x7 & ~x8 ;
  assign n24 = n23 ^ n20 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = ~x6 & x8 ;
  assign n28 = n27 ^ x4 ;
  assign n29 = x4 & n28 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = n30 ^ x4 ;
  assign n32 = ~n26 & ~n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ x4 ;
  assign n35 = n22 & n34 ;
  assign n36 = n35 ^ n20 ;
  assign n37 = n18 & ~n36 ;
  assign n38 = x2 & ~n37 ;
  assign n39 = ~x2 & x5 ;
  assign n40 = x6 & n39 ;
  assign n41 = x1 & n40 ;
  assign n42 = ~x7 & x8 ;
  assign n43 = n42 ^ x7 ;
  assign n44 = x4 & n43 ;
  assign n45 = n44 ^ x7 ;
  assign n46 = n41 & n45 ;
  assign n47 = ~x4 & ~x5 ;
  assign n48 = x7 & ~x8 ;
  assign n49 = n47 & n48 ;
  assign n53 = ~x4 & x7 ;
  assign n54 = x8 & n53 ;
  assign n55 = x2 & n42 ;
  assign n56 = ~n54 & ~n55 ;
  assign n50 = ~x2 & x4 ;
  assign n51 = x1 & ~x7 ;
  assign n52 = ~n50 & n51 ;
  assign n57 = n56 ^ n52 ;
  assign n58 = ~x5 & ~n57 ;
  assign n59 = n58 ^ n56 ;
  assign n60 = ~n49 & n59 ;
  assign n61 = x6 & ~n60 ;
  assign n62 = x2 & x4 ;
  assign n63 = n23 & n62 ;
  assign n64 = ~x5 & ~n63 ;
  assign n65 = ~x1 & ~n64 ;
  assign n66 = x6 & x7 ;
  assign n67 = ~n19 & ~n66 ;
  assign n68 = x8 ^ x7 ;
  assign n69 = ~n67 & ~n68 ;
  assign n70 = x5 & ~n69 ;
  assign n71 = ~x2 & ~x6 ;
  assign n72 = n53 ^ x8 ;
  assign n73 = n72 ^ n53 ;
  assign n74 = n53 ^ x4 ;
  assign n75 = n73 & n74 ;
  assign n76 = n75 ^ n53 ;
  assign n77 = n71 & n76 ;
  assign n78 = n70 & ~n77 ;
  assign n79 = n65 & ~n78 ;
  assign n80 = ~x5 & ~n14 ;
  assign n81 = n13 & ~n27 ;
  assign n82 = n80 & n81 ;
  assign n83 = x4 & n82 ;
  assign n84 = ~n79 & ~n83 ;
  assign n88 = ~x4 & x8 ;
  assign n89 = x4 & ~x6 ;
  assign n90 = n48 & n89 ;
  assign n91 = ~n88 & ~n90 ;
  assign n92 = n65 & ~n91 ;
  assign n93 = ~x4 & n51 ;
  assign n94 = ~n49 & ~n93 ;
  assign n95 = ~n92 & n94 ;
  assign n85 = ~n13 & ~n14 ;
  assign n86 = ~n66 & ~n85 ;
  assign n87 = ~n80 & n86 ;
  assign n96 = n95 ^ n87 ;
  assign n97 = n96 ^ n95 ;
  assign n98 = n95 ^ x4 ;
  assign n99 = n98 ^ n95 ;
  assign n100 = n97 & n99 ;
  assign n101 = n100 ^ n95 ;
  assign n102 = ~x2 & ~n101 ;
  assign n103 = n102 ^ n95 ;
  assign n104 = n84 & n103 ;
  assign n105 = ~n61 & n104 ;
  assign n106 = n105 ^ x3 ;
  assign n107 = n106 ^ n105 ;
  assign n108 = x5 & n10 ;
  assign n109 = ~n66 & ~n108 ;
  assign n110 = ~x2 & ~x4 ;
  assign n111 = ~x1 & n110 ;
  assign n112 = ~n109 & n111 ;
  assign n155 = x6 & ~x7 ;
  assign n156 = ~n89 & ~n155 ;
  assign n157 = x2 & ~n53 ;
  assign n158 = n156 & n157 ;
  assign n159 = ~x2 & ~n13 ;
  assign n160 = n159 ^ n67 ;
  assign n161 = n159 ^ n53 ;
  assign n162 = n159 ^ x1 ;
  assign n163 = n159 & ~n162 ;
  assign n164 = n163 ^ n159 ;
  assign n165 = n161 & n164 ;
  assign n166 = n165 ^ n163 ;
  assign n167 = n166 ^ n159 ;
  assign n168 = n167 ^ x1 ;
  assign n169 = ~n160 & ~n168 ;
  assign n170 = n169 ^ n159 ;
  assign n171 = ~n158 & ~n170 ;
  assign n172 = ~x5 & ~n171 ;
  assign n173 = n51 ^ x5 ;
  assign n174 = n173 ^ n110 ;
  assign n182 = n174 ^ n173 ;
  assign n175 = n62 & n155 ;
  assign n176 = n175 ^ n174 ;
  assign n177 = n176 ^ n173 ;
  assign n178 = n174 ^ n51 ;
  assign n179 = n178 ^ n175 ;
  assign n180 = n179 ^ n177 ;
  assign n181 = ~n177 & ~n180 ;
  assign n183 = n182 ^ n181 ;
  assign n184 = n183 ^ n177 ;
  assign n185 = ~x6 & n13 ;
  assign n186 = n185 ^ n173 ;
  assign n187 = n181 ^ n177 ;
  assign n188 = ~n186 & ~n187 ;
  assign n189 = n188 ^ n173 ;
  assign n190 = ~n184 & n189 ;
  assign n191 = n190 ^ n173 ;
  assign n192 = n191 ^ x5 ;
  assign n193 = n192 ^ n173 ;
  assign n194 = ~n172 & ~n193 ;
  assign n134 = ~n13 & ~n50 ;
  assign n135 = ~n89 & ~n134 ;
  assign n115 = x4 ^ x2 ;
  assign n113 = x4 ^ x1 ;
  assign n114 = n113 ^ x6 ;
  assign n116 = n115 ^ n114 ;
  assign n117 = n116 ^ x4 ;
  assign n118 = n117 ^ x7 ;
  assign n119 = n118 ^ n117 ;
  assign n122 = n114 ^ x6 ;
  assign n123 = n122 ^ n116 ;
  assign n124 = n123 ^ n117 ;
  assign n125 = ~n117 & ~n124 ;
  assign n120 = ~x6 & n116 ;
  assign n128 = n125 ^ n120 ;
  assign n121 = n120 ^ n119 ;
  assign n126 = n125 ^ n117 ;
  assign n127 = ~n121 & ~n126 ;
  assign n129 = n128 ^ n127 ;
  assign n130 = ~n119 & n129 ;
  assign n131 = n130 ^ n125 ;
  assign n132 = n131 ^ n127 ;
  assign n133 = n132 ^ n114 ;
  assign n136 = n135 ^ n133 ;
  assign n137 = n136 ^ x5 ;
  assign n144 = n137 ^ n136 ;
  assign n138 = n137 ^ n110 ;
  assign n139 = n138 ^ n136 ;
  assign n140 = n137 ^ n133 ;
  assign n141 = n140 ^ n110 ;
  assign n142 = n141 ^ n139 ;
  assign n143 = n139 & ~n142 ;
  assign n145 = n144 ^ n143 ;
  assign n146 = n145 ^ n139 ;
  assign n147 = n136 ^ x4 ;
  assign n148 = n143 ^ n139 ;
  assign n149 = n147 & n148 ;
  assign n150 = n149 ^ n136 ;
  assign n151 = ~n146 & ~n150 ;
  assign n152 = n151 ^ n136 ;
  assign n153 = n152 ^ n135 ;
  assign n154 = n153 ^ n136 ;
  assign n195 = n194 ^ n154 ;
  assign n196 = ~x8 & ~n195 ;
  assign n197 = n196 ^ n154 ;
  assign n198 = ~n112 & ~n197 ;
  assign n199 = n198 ^ n105 ;
  assign n200 = n107 & n199 ;
  assign n201 = n200 ^ n105 ;
  assign n202 = ~n46 & n201 ;
  assign n203 = ~n38 & n202 ;
  assign n204 = ~x0 & ~n203 ;
  assign n213 = n27 & n47 ;
  assign n205 = n47 ^ x0 ;
  assign n206 = n205 ^ x0 ;
  assign n207 = x8 ^ x0 ;
  assign n208 = n207 ^ x0 ;
  assign n209 = ~n206 & ~n208 ;
  assign n210 = n209 ^ x0 ;
  assign n211 = x6 & ~n210 ;
  assign n212 = n211 ^ x0 ;
  assign n214 = n213 ^ n212 ;
  assign n215 = n214 ^ n213 ;
  assign n216 = ~x4 & ~n14 ;
  assign n217 = n216 ^ n213 ;
  assign n218 = n217 ^ n213 ;
  assign n219 = n215 & ~n218 ;
  assign n220 = n219 ^ n213 ;
  assign n221 = x7 & n220 ;
  assign n222 = n221 ^ n213 ;
  assign n223 = x0 & x5 ;
  assign n224 = n88 & n223 ;
  assign n225 = n15 ^ n14 ;
  assign n226 = n225 ^ n15 ;
  assign n227 = n226 ^ n224 ;
  assign n228 = ~x5 & x6 ;
  assign n229 = ~n23 & ~n228 ;
  assign n230 = n229 ^ x0 ;
  assign n231 = ~n229 & ~n230 ;
  assign n232 = n231 ^ n15 ;
  assign n233 = n232 ^ n229 ;
  assign n234 = n227 & ~n233 ;
  assign n235 = n234 ^ n231 ;
  assign n236 = n235 ^ n229 ;
  assign n237 = ~n224 & ~n236 ;
  assign n238 = n237 ^ n224 ;
  assign n239 = ~n222 & ~n238 ;
  assign n240 = ~x2 & ~x3 ;
  assign n241 = ~n239 & n240 ;
  assign n242 = ~x1 & n241 ;
  assign n243 = ~n204 & ~n242 ;
  assign y0 = ~n243 ;
endmodule
