module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 ;
  assign n22 = x15 ^ x12 ;
  assign n23 = n22 ^ x13 ;
  assign n30 = n23 ^ n22 ;
  assign n24 = n23 ^ x14 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n23 ^ x15 ;
  assign n27 = n26 ^ x14 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = ~n25 & ~n28 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n31 ^ n25 ;
  assign n33 = x15 & ~x16 ;
  assign n34 = x17 & n33 ;
  assign n35 = n34 ^ n22 ;
  assign n36 = n29 ^ n25 ;
  assign n37 = n35 & ~n36 ;
  assign n38 = n37 ^ n22 ;
  assign n39 = ~n32 & n38 ;
  assign n40 = n39 ^ n22 ;
  assign n41 = n40 ^ x12 ;
  assign n42 = n41 ^ n22 ;
  assign n43 = x11 & n42 ;
  assign n44 = ~x1 & ~x8 ;
  assign n45 = ~x0 & n44 ;
  assign n46 = ~x2 & ~x7 ;
  assign n47 = x10 & x20 ;
  assign n48 = ~x5 & ~x6 ;
  assign n49 = n47 & n48 ;
  assign n50 = ~x3 & ~x4 ;
  assign n51 = ~x9 & ~x19 ;
  assign n52 = n50 & n51 ;
  assign n53 = n49 & n52 ;
  assign n54 = x11 & ~x13 ;
  assign n55 = ~x18 & n54 ;
  assign n56 = ~x12 & ~n55 ;
  assign n57 = n53 & ~n56 ;
  assign n58 = n46 & n57 ;
  assign n59 = n45 & n58 ;
  assign n60 = ~n43 & n59 ;
  assign y0 = n60 ;
endmodule
