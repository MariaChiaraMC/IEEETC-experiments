module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n12 = ~x0 & ~x1 ;
  assign n13 = x9 & ~x10 ;
  assign n14 = x8 & n13 ;
  assign n15 = ~x4 & ~n14 ;
  assign n16 = ~x3 & ~n15 ;
  assign n17 = x9 ^ x8 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = ~x7 & ~n18 ;
  assign n20 = n19 ^ n13 ;
  assign n21 = ~x6 & n20 ;
  assign n22 = ~n16 & ~n21 ;
  assign n23 = x5 & ~n22 ;
  assign n24 = ~x4 & ~x6 ;
  assign n25 = x3 & ~n24 ;
  assign n26 = ~n15 & n25 ;
  assign n27 = x2 & n26 ;
  assign n28 = ~n23 & ~n27 ;
  assign n29 = ~n12 & ~n28 ;
  assign y0 = n29 ;
endmodule
