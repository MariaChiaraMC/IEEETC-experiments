module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 ;
  output y0 ;
  wire n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 ;
  assign n29 = x14 ^ x4 ;
  assign n30 = x14 ^ x3 ;
  assign n31 = n30 ^ x14 ;
  assign n32 = n31 ^ n29 ;
  assign n41 = x16 ^ x15 ;
  assign n42 = x18 ^ x16 ;
  assign n43 = ~n41 & ~n42 ;
  assign n44 = x24 & n43 ;
  assign n33 = x21 & x22 ;
  assign n34 = x17 & ~x19 ;
  assign n35 = x18 & n34 ;
  assign n36 = x20 & ~n35 ;
  assign n37 = ~n33 & ~n36 ;
  assign n38 = n37 ^ x13 ;
  assign n39 = ~x16 & ~n38 ;
  assign n40 = n39 ^ x13 ;
  assign n45 = n44 ^ n40 ;
  assign n46 = ~x14 & ~n45 ;
  assign n47 = n46 ^ n44 ;
  assign n48 = ~n32 & ~n47 ;
  assign n49 = n48 ^ n46 ;
  assign n50 = n49 ^ n44 ;
  assign n51 = n50 ^ x14 ;
  assign n52 = n29 & n51 ;
  assign n53 = x2 & n52 ;
  assign n54 = x2 ^ x0 ;
  assign n55 = x4 ^ x2 ;
  assign n56 = n55 ^ x4 ;
  assign n57 = ~x3 & ~x4 ;
  assign n58 = ~x10 & x12 ;
  assign n59 = ~x11 & n58 ;
  assign n60 = ~x9 & ~n59 ;
  assign n61 = ~x8 & ~n60 ;
  assign n62 = x10 & ~x11 ;
  assign n63 = ~x13 & n62 ;
  assign n64 = x7 & ~n63 ;
  assign n65 = ~n61 & n64 ;
  assign n66 = x6 & ~n65 ;
  assign n67 = n57 & n66 ;
  assign n68 = x4 & ~x14 ;
  assign n70 = x16 & ~x19 ;
  assign n71 = x20 & ~n70 ;
  assign n72 = n68 & ~n71 ;
  assign n73 = x26 & x27 ;
  assign n74 = ~n33 & ~n73 ;
  assign n75 = x4 & x25 ;
  assign n76 = x14 & n75 ;
  assign n77 = x18 & n76 ;
  assign n78 = n74 & n77 ;
  assign n79 = ~n72 & ~n78 ;
  assign n69 = x15 & n68 ;
  assign n80 = n79 ^ n69 ;
  assign n81 = ~x3 & ~n80 ;
  assign n82 = n81 ^ n79 ;
  assign n83 = ~n67 & n82 ;
  assign n84 = n83 ^ x4 ;
  assign n85 = ~n56 & ~n84 ;
  assign n86 = n85 ^ x4 ;
  assign n87 = ~n54 & n86 ;
  assign n88 = n87 ^ x0 ;
  assign n89 = ~n53 & ~n88 ;
  assign n90 = ~x5 & ~n89 ;
  assign n91 = x14 & n57 ;
  assign n92 = ~n68 & ~n91 ;
  assign n93 = x0 & ~n92 ;
  assign n96 = n68 ^ x0 ;
  assign n97 = n96 ^ x0 ;
  assign n94 = x5 ^ x0 ;
  assign n95 = n94 ^ x0 ;
  assign n98 = n97 ^ n95 ;
  assign n99 = x22 & ~x23 ;
  assign n100 = n99 ^ x0 ;
  assign n101 = n100 ^ x0 ;
  assign n102 = n101 ^ n97 ;
  assign n103 = n97 & n102 ;
  assign n104 = n103 ^ n97 ;
  assign n105 = n98 & n104 ;
  assign n106 = n105 ^ n103 ;
  assign n107 = n106 ^ x0 ;
  assign n108 = n107 ^ n97 ;
  assign n109 = x2 & n108 ;
  assign n110 = n109 ^ x0 ;
  assign n111 = n110 ^ x3 ;
  assign n112 = n111 ^ n110 ;
  assign n113 = x2 & x5 ;
  assign n114 = x14 & ~n113 ;
  assign n115 = x0 & ~n114 ;
  assign n116 = x5 & n34 ;
  assign n117 = ~x4 & ~x14 ;
  assign n118 = ~x16 & n117 ;
  assign n119 = n116 & n118 ;
  assign n120 = ~x21 & ~x22 ;
  assign n121 = ~x13 & x16 ;
  assign n122 = n68 & n121 ;
  assign n123 = ~n120 & n122 ;
  assign n124 = ~n119 & ~n123 ;
  assign n125 = x2 & ~n124 ;
  assign n126 = ~n115 & ~n125 ;
  assign n127 = n126 ^ n110 ;
  assign n128 = n112 & ~n127 ;
  assign n129 = n128 ^ n110 ;
  assign n130 = ~n93 & ~n129 ;
  assign n131 = ~n90 & n130 ;
  assign n132 = x1 & ~n131 ;
  assign y0 = n132 ;
endmodule
