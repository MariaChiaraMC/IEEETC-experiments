// Benchmark "./pla/xparc.pla_dbb_orig_1NonExact" written by ABC on Fri Nov 20 10:30:38 2020

module \./pla/xparc.pla_dbb_orig_1NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = 1'b1;
endmodule


