module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 ;
  assign n16 = x12 ^ x11 ;
  assign n17 = x9 & x10 ;
  assign n18 = ~x13 & x14 ;
  assign n19 = n17 & ~n18 ;
  assign n77 = ~x0 & x1 ;
  assign n108 = x3 & ~x10 ;
  assign n109 = n77 & n108 ;
  assign n110 = x2 & n109 ;
  assign n112 = n110 ^ x9 ;
  assign n122 = n112 ^ n110 ;
  assign n123 = n122 ^ n110 ;
  assign n124 = ~n122 & ~n123 ;
  assign n96 = ~x2 & ~x3 ;
  assign n97 = x0 & ~n96 ;
  assign n98 = ~x1 & n97 ;
  assign n114 = x14 & ~n98 ;
  assign n115 = x10 & ~n114 ;
  assign n20 = x2 & x7 ;
  assign n21 = ~x3 & ~x4 ;
  assign n22 = ~x0 & ~x2 ;
  assign n23 = n21 & n22 ;
  assign n24 = x9 & n23 ;
  assign n25 = ~x6 & n24 ;
  assign n26 = ~n20 & ~n25 ;
  assign n27 = ~x1 & ~n26 ;
  assign n28 = x9 ^ x7 ;
  assign n29 = n28 ^ x7 ;
  assign n30 = ~x3 & x4 ;
  assign n31 = x6 & x7 ;
  assign n32 = n30 & n31 ;
  assign n33 = x2 & x6 ;
  assign n34 = ~x0 & ~x1 ;
  assign n35 = ~n33 & n34 ;
  assign n36 = ~n32 & n35 ;
  assign n37 = ~x0 & ~n30 ;
  assign n38 = ~n22 & ~n37 ;
  assign n40 = x4 ^ x3 ;
  assign n39 = x4 ^ x2 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = n42 ^ n40 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = n44 ^ x1 ;
  assign n46 = ~n43 & ~n45 ;
  assign n47 = n46 ^ n42 ;
  assign n48 = n47 ^ n43 ;
  assign n52 = n43 ^ x6 ;
  assign n53 = ~n43 & n52 ;
  assign n49 = n42 ^ x2 ;
  assign n50 = n49 ^ n43 ;
  assign n51 = x7 & n50 ;
  assign n54 = n53 ^ n51 ;
  assign n55 = n54 ^ n42 ;
  assign n56 = n55 ^ x2 ;
  assign n57 = n56 ^ n43 ;
  assign n58 = n57 ^ x1 ;
  assign n59 = x2 & ~n58 ;
  assign n60 = n59 ^ n51 ;
  assign n61 = n60 ^ n42 ;
  assign n62 = n61 ^ n43 ;
  assign n63 = n62 ^ x1 ;
  assign n64 = n48 & ~n63 ;
  assign n65 = n64 ^ n51 ;
  assign n66 = n65 ^ n46 ;
  assign n67 = n66 ^ n59 ;
  assign n68 = n67 ^ x1 ;
  assign n69 = n68 ^ x1 ;
  assign n70 = n38 & n69 ;
  assign n71 = ~n36 & ~n70 ;
  assign n72 = n71 ^ x7 ;
  assign n73 = ~n29 & n72 ;
  assign n74 = n73 ^ x7 ;
  assign n75 = ~n27 & n74 ;
  assign n76 = x5 & ~n75 ;
  assign n78 = ~x5 & n21 ;
  assign n79 = x2 & ~n78 ;
  assign n80 = n77 & ~n79 ;
  assign n81 = ~n20 & n80 ;
  assign n82 = x1 & ~x3 ;
  assign n83 = x4 & ~n33 ;
  assign n84 = n83 ^ x6 ;
  assign n85 = n84 ^ n82 ;
  assign n86 = x0 & ~x5 ;
  assign n87 = n86 ^ x5 ;
  assign n88 = x6 & n87 ;
  assign n89 = n88 ^ x5 ;
  assign n90 = n85 & ~n89 ;
  assign n91 = n90 ^ n88 ;
  assign n92 = n91 ^ x5 ;
  assign n93 = n92 ^ x6 ;
  assign n94 = n82 & ~n93 ;
  assign n95 = ~n81 & ~n94 ;
  assign n99 = x9 & ~n23 ;
  assign n100 = x3 & ~x4 ;
  assign n101 = n86 & ~n100 ;
  assign n102 = x2 & n101 ;
  assign n103 = ~n99 & ~n102 ;
  assign n104 = ~x10 & n103 ;
  assign n105 = ~n98 & n104 ;
  assign n106 = n95 & n105 ;
  assign n107 = ~n76 & n106 ;
  assign n111 = n110 ^ n107 ;
  assign n113 = n112 ^ n111 ;
  assign n116 = n115 ^ n113 ;
  assign n117 = n116 ^ n113 ;
  assign n118 = n113 ^ n112 ;
  assign n119 = n118 ^ n110 ;
  assign n120 = ~n117 & ~n119 ;
  assign n127 = n124 ^ n120 ;
  assign n121 = n120 ^ x13 ;
  assign n125 = n124 ^ n122 ;
  assign n126 = n121 & ~n125 ;
  assign n128 = n127 ^ n126 ;
  assign n129 = x13 & n128 ;
  assign n130 = n129 ^ n120 ;
  assign n131 = n130 ^ n124 ;
  assign n132 = n131 ^ n126 ;
  assign n133 = n132 ^ x9 ;
  assign n134 = ~n19 & n133 ;
  assign n135 = n134 ^ x12 ;
  assign n136 = n135 ^ n134 ;
  assign n137 = n136 ^ n16 ;
  assign n138 = n17 ^ x13 ;
  assign n139 = n17 & ~n138 ;
  assign n140 = n139 ^ n134 ;
  assign n141 = n140 ^ n17 ;
  assign n142 = ~n137 & ~n141 ;
  assign n143 = n142 ^ n139 ;
  assign n144 = n143 ^ n17 ;
  assign n145 = ~n16 & n144 ;
  assign y0 = n145 ;
endmodule
