// Benchmark "./pla/add6.pla_res_0NonExact" written by ABC on Fri Nov 20 10:16:55 2020

module \./pla/add6.pla_res_0NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = x0;
endmodule


