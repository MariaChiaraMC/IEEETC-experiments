module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 ;
  assign n8 = x1 & ~x5 ;
  assign n9 = ~x2 & ~n8 ;
  assign n10 = ~x3 & n9 ;
  assign n11 = ~x5 & ~x6 ;
  assign n12 = x1 & x2 ;
  assign n13 = n11 & n12 ;
  assign n14 = ~n10 & ~n13 ;
  assign n15 = x4 & ~n14 ;
  assign n16 = x4 & ~x6 ;
  assign n17 = ~x1 & x5 ;
  assign n18 = x3 & ~n17 ;
  assign n19 = ~n16 & ~n18 ;
  assign n20 = x4 ^ x2 ;
  assign n21 = n19 & n20 ;
  assign n22 = ~n15 & ~n21 ;
  assign n23 = ~x0 & ~n22 ;
  assign n24 = x0 & ~x2 ;
  assign n25 = n8 & n16 ;
  assign n26 = n24 & n25 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = n8 ^ x2 ;
  assign n29 = n28 ^ n8 ;
  assign n30 = n29 ^ n17 ;
  assign n31 = ~x1 & x6 ;
  assign n32 = n31 ^ x0 ;
  assign n33 = ~n31 & ~n32 ;
  assign n34 = n33 ^ n8 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = n30 & n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ n31 ;
  assign n39 = ~n17 & ~n38 ;
  assign n40 = n39 ^ x2 ;
  assign n41 = ~x4 & n40 ;
  assign n42 = ~x1 & x4 ;
  assign n43 = x5 ^ x2 ;
  assign n44 = n43 ^ x5 ;
  assign n45 = x5 ^ x0 ;
  assign n46 = n44 & n45 ;
  assign n47 = n46 ^ x5 ;
  assign n48 = n42 & n47 ;
  assign n49 = ~n41 & ~n48 ;
  assign n50 = n49 ^ x3 ;
  assign n51 = n50 ^ n49 ;
  assign n60 = n20 ^ x2 ;
  assign n52 = x2 ^ x1 ;
  assign n53 = n52 ^ x4 ;
  assign n54 = n53 ^ n20 ;
  assign n55 = n54 ^ n20 ;
  assign n56 = n55 ^ x2 ;
  assign n57 = n54 ^ n43 ;
  assign n58 = n57 ^ n56 ;
  assign n59 = n56 & ~n58 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = n61 ^ n56 ;
  assign n63 = x6 ^ x2 ;
  assign n64 = n63 ^ x2 ;
  assign n65 = n59 ^ n56 ;
  assign n66 = n64 & n65 ;
  assign n67 = n66 ^ x2 ;
  assign n68 = n62 & n67 ;
  assign n69 = n68 ^ x2 ;
  assign n70 = n69 ^ n53 ;
  assign n71 = n70 ^ x2 ;
  assign n72 = x0 & ~n71 ;
  assign n73 = x2 & x5 ;
  assign n74 = ~x4 & ~x6 ;
  assign n75 = n73 & ~n74 ;
  assign n76 = ~n31 & n75 ;
  assign n77 = ~x1 & ~x2 ;
  assign n78 = n77 ^ n74 ;
  assign n79 = n78 ^ n74 ;
  assign n80 = ~x0 & ~n20 ;
  assign n81 = n80 ^ n74 ;
  assign n82 = ~n79 & n81 ;
  assign n83 = n82 ^ n74 ;
  assign n84 = ~x5 & n83 ;
  assign n85 = ~n76 & ~n84 ;
  assign n86 = ~n72 & n85 ;
  assign n87 = n86 ^ n49 ;
  assign n88 = n51 & n87 ;
  assign n89 = n88 ^ n49 ;
  assign n90 = n89 ^ n23 ;
  assign n91 = n27 & ~n90 ;
  assign n92 = n91 ^ n88 ;
  assign n93 = n92 ^ n49 ;
  assign n94 = n93 ^ n26 ;
  assign n95 = ~n23 & ~n94 ;
  assign n96 = n95 ^ n23 ;
  assign y0 = n96 ;
endmodule
