module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 ;
  assign n9 = x7 ^ x3 ;
  assign n20 = x7 ^ x2 ;
  assign n10 = x5 ^ x1 ;
  assign n11 = x5 ^ x0 ;
  assign n12 = n11 ^ x5 ;
  assign n13 = x5 ^ x4 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = n12 & n14 ;
  assign n16 = n15 ^ x5 ;
  assign n17 = n10 & ~n16 ;
  assign n18 = n17 ^ x1 ;
  assign n19 = n18 ^ x7 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = x7 ^ x6 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n21 & n23 ;
  assign n25 = n24 ^ n20 ;
  assign n26 = n9 & ~n25 ;
  assign n27 = n26 ^ x3 ;
  assign y0 = n27 ;
endmodule
