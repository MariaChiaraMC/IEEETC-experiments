module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 ;
  assign n10 = x3 & ~x8 ;
  assign n11 = ~x2 & n10 ;
  assign n12 = x2 & x3 ;
  assign n13 = ~x6 & ~x8 ;
  assign n14 = ~n12 & ~n13 ;
  assign n15 = ~x1 & ~n14 ;
  assign n16 = ~n11 & ~n15 ;
  assign n17 = ~x0 & x4 ;
  assign n18 = x5 & n17 ;
  assign n19 = ~n16 & n18 ;
  assign n20 = x5 & x6 ;
  assign n21 = x0 & ~x4 ;
  assign n22 = ~x1 & ~x3 ;
  assign n23 = n21 & n22 ;
  assign n24 = ~x2 & n23 ;
  assign n25 = x2 & ~x8 ;
  assign n26 = ~x3 & n25 ;
  assign n27 = n26 ^ x4 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = x1 & x8 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = ~n28 & n30 ;
  assign n32 = n31 ^ n26 ;
  assign n33 = ~x0 & n32 ;
  assign n34 = ~n24 & ~n33 ;
  assign n35 = ~n20 & ~n34 ;
  assign n36 = ~x0 & ~x4 ;
  assign n37 = n12 & n29 ;
  assign n38 = ~x2 & ~x5 ;
  assign n39 = n38 ^ x3 ;
  assign n40 = n38 ^ x1 ;
  assign n41 = n40 ^ x1 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = ~x1 & ~x2 ;
  assign n44 = ~x5 & x8 ;
  assign n45 = ~n43 & ~n44 ;
  assign n46 = n45 ^ x6 ;
  assign n47 = ~x6 & n46 ;
  assign n48 = n47 ^ x1 ;
  assign n49 = n48 ^ x6 ;
  assign n50 = ~n42 & n49 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = n51 ^ x6 ;
  assign n53 = n39 & ~n52 ;
  assign n54 = n53 ^ n38 ;
  assign n55 = ~n37 & ~n54 ;
  assign n56 = n36 & ~n55 ;
  assign n57 = ~n35 & ~n56 ;
  assign n58 = ~x5 & ~x6 ;
  assign n59 = x4 & ~n58 ;
  assign n60 = x8 & n43 ;
  assign n61 = ~n59 & n60 ;
  assign n62 = n36 & ~n43 ;
  assign n63 = x8 ^ x1 ;
  assign n64 = n63 ^ x8 ;
  assign n65 = n58 ^ x8 ;
  assign n66 = n64 & ~n65 ;
  assign n67 = n66 ^ x8 ;
  assign n68 = n62 & ~n67 ;
  assign n69 = ~n61 & ~n68 ;
  assign n70 = n20 ^ x4 ;
  assign n71 = x8 ^ x0 ;
  assign n72 = n71 ^ x0 ;
  assign n73 = n43 ^ x0 ;
  assign n74 = ~n72 & ~n73 ;
  assign n75 = n74 ^ x0 ;
  assign n76 = n75 ^ n20 ;
  assign n77 = n70 & ~n76 ;
  assign n78 = n77 ^ n74 ;
  assign n79 = n78 ^ x0 ;
  assign n80 = n79 ^ x4 ;
  assign n81 = n20 & ~n80 ;
  assign n82 = n81 ^ n20 ;
  assign n83 = n69 & ~n82 ;
  assign n84 = ~x3 & ~n83 ;
  assign n85 = n57 & ~n84 ;
  assign n86 = ~n19 & n85 ;
  assign n87 = x7 & ~n86 ;
  assign n88 = n12 & n13 ;
  assign n89 = ~x1 & ~x5 ;
  assign n90 = x2 & n89 ;
  assign n91 = ~x3 & x8 ;
  assign n92 = n58 & n91 ;
  assign n93 = ~n90 & ~n92 ;
  assign n94 = ~n88 & n93 ;
  assign n95 = x4 & ~n94 ;
  assign n96 = x6 & ~x8 ;
  assign n97 = n43 & n96 ;
  assign n98 = ~x4 & n97 ;
  assign n99 = x3 & ~n96 ;
  assign n100 = ~x4 & x5 ;
  assign n101 = x1 & ~n91 ;
  assign n102 = n100 & ~n101 ;
  assign n103 = ~n99 & n102 ;
  assign n104 = n103 ^ n98 ;
  assign n105 = ~x3 & ~x6 ;
  assign n106 = n100 & n105 ;
  assign n107 = ~x1 & x8 ;
  assign n108 = x1 & ~x5 ;
  assign n109 = x4 ^ x3 ;
  assign n110 = n109 ^ x4 ;
  assign n111 = n96 ^ x4 ;
  assign n112 = n110 & ~n111 ;
  assign n113 = n112 ^ x4 ;
  assign n114 = n108 & ~n113 ;
  assign n115 = ~n107 & ~n114 ;
  assign n116 = ~n106 & n115 ;
  assign n117 = n116 ^ x2 ;
  assign n118 = n117 ^ n116 ;
  assign n119 = n116 ^ n29 ;
  assign n120 = ~n118 & ~n119 ;
  assign n121 = n120 ^ n116 ;
  assign n122 = n121 ^ n98 ;
  assign n123 = n104 & ~n122 ;
  assign n124 = n123 ^ n120 ;
  assign n125 = n124 ^ n116 ;
  assign n126 = n125 ^ n103 ;
  assign n127 = ~n98 & ~n126 ;
  assign n128 = n127 ^ n98 ;
  assign n129 = ~n95 & ~n128 ;
  assign n130 = ~x7 & ~n129 ;
  assign n131 = n10 & n100 ;
  assign n132 = x2 ^ x1 ;
  assign n133 = n131 & ~n132 ;
  assign n134 = x8 & n22 ;
  assign n135 = n134 ^ x4 ;
  assign n136 = n135 ^ n133 ;
  assign n137 = x7 & ~n20 ;
  assign n138 = x1 & ~x2 ;
  assign n139 = x3 & n58 ;
  assign n140 = n138 & ~n139 ;
  assign n141 = ~n137 & n140 ;
  assign n142 = n141 ^ x5 ;
  assign n143 = n11 ^ x1 ;
  assign n144 = n143 ^ n11 ;
  assign n145 = n88 ^ n11 ;
  assign n146 = n144 & n145 ;
  assign n147 = n146 ^ n11 ;
  assign n148 = n147 ^ n141 ;
  assign n149 = n142 & ~n148 ;
  assign n150 = n149 ^ n146 ;
  assign n151 = n150 ^ n11 ;
  assign n152 = n151 ^ x5 ;
  assign n153 = ~n141 & ~n152 ;
  assign n154 = n153 ^ n141 ;
  assign n155 = n154 ^ n141 ;
  assign n156 = n155 ^ n20 ;
  assign n157 = ~n134 & n156 ;
  assign n158 = n157 ^ n20 ;
  assign n159 = ~n136 & ~n158 ;
  assign n160 = n159 ^ n157 ;
  assign n161 = n160 ^ n20 ;
  assign n162 = n161 ^ n134 ;
  assign n163 = ~n133 & n162 ;
  assign n164 = ~n130 & n163 ;
  assign n165 = ~x0 & ~n164 ;
  assign n166 = ~x4 & ~x5 ;
  assign n167 = ~x7 & ~n166 ;
  assign n168 = x6 & n21 ;
  assign n169 = ~n167 & ~n168 ;
  assign n170 = n91 & ~n169 ;
  assign n171 = n43 & n170 ;
  assign n172 = ~n165 & ~n171 ;
  assign n173 = ~n87 & n172 ;
  assign y0 = ~n173 ;
endmodule
