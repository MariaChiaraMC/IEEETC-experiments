module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 ;
  assign n9 = ~x4 & ~x5 ;
  assign n10 = ~x6 & ~x7 ;
  assign n11 = ~x4 & n10 ;
  assign n12 = x0 & ~n11 ;
  assign n13 = ~n9 & n12 ;
  assign n14 = x5 & ~x7 ;
  assign n15 = ~x0 & ~n14 ;
  assign n20 = n15 ^ x3 ;
  assign n28 = n20 ^ n15 ;
  assign n16 = x6 & ~x7 ;
  assign n17 = x5 & ~x6 ;
  assign n18 = ~n16 & ~n17 ;
  assign n19 = n18 ^ n15 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n22 ^ n15 ;
  assign n24 = n21 ^ x4 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n23 & n26 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = ~x5 & x7 ;
  assign n32 = n31 ^ n15 ;
  assign n33 = n27 ^ n23 ;
  assign n34 = ~n32 & n33 ;
  assign n35 = n34 ^ n15 ;
  assign n36 = n30 & n35 ;
  assign n37 = n36 ^ n15 ;
  assign n38 = n37 ^ x3 ;
  assign n39 = n38 ^ n15 ;
  assign n40 = ~n13 & ~n39 ;
  assign n41 = ~x2 & ~n40 ;
  assign n42 = x4 & ~x5 ;
  assign n43 = x2 & ~x6 ;
  assign n44 = ~n42 & ~n43 ;
  assign n45 = x0 & ~n44 ;
  assign n46 = x4 & x5 ;
  assign n47 = n46 ^ x6 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = n48 ^ x2 ;
  assign n50 = n31 ^ x4 ;
  assign n51 = ~n31 & ~n50 ;
  assign n52 = n51 ^ n46 ;
  assign n53 = n52 ^ n31 ;
  assign n54 = n49 & n53 ;
  assign n55 = n54 ^ n51 ;
  assign n56 = n55 ^ n31 ;
  assign n57 = x2 & ~n56 ;
  assign n58 = n57 ^ x2 ;
  assign n59 = ~n45 & ~n58 ;
  assign n60 = n59 ^ x3 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = n61 ^ n41 ;
  assign n64 = x4 ^ x2 ;
  assign n65 = n64 ^ x2 ;
  assign n63 = x6 ^ x2 ;
  assign n66 = n65 ^ n63 ;
  assign n67 = x7 ^ x2 ;
  assign n68 = n67 ^ x2 ;
  assign n69 = n68 ^ n65 ;
  assign n70 = ~n65 & n69 ;
  assign n71 = n70 ^ n65 ;
  assign n72 = ~n66 & ~n71 ;
  assign n73 = n72 ^ n70 ;
  assign n74 = n73 ^ x2 ;
  assign n75 = n74 ^ n65 ;
  assign n76 = ~x5 & ~n75 ;
  assign n77 = n76 ^ x0 ;
  assign n78 = n76 & ~n77 ;
  assign n79 = n78 ^ n59 ;
  assign n80 = n79 ^ n76 ;
  assign n81 = ~n62 & ~n80 ;
  assign n82 = n81 ^ n78 ;
  assign n83 = n82 ^ n76 ;
  assign n84 = ~n41 & n83 ;
  assign n85 = n84 ^ n41 ;
  assign n86 = ~x1 & n85 ;
  assign n87 = x1 & n17 ;
  assign n88 = ~n14 & ~n87 ;
  assign n89 = ~x4 & ~n88 ;
  assign n90 = ~x3 & ~x6 ;
  assign n91 = n90 ^ x1 ;
  assign n92 = n9 & n91 ;
  assign n93 = ~n89 & ~n92 ;
  assign n94 = ~x2 & ~n93 ;
  assign n95 = x1 & ~x3 ;
  assign n96 = n95 ^ n63 ;
  assign n97 = n46 ^ n9 ;
  assign n98 = x6 & n97 ;
  assign n99 = n98 ^ n9 ;
  assign n100 = n96 & ~n99 ;
  assign n101 = n100 ^ n98 ;
  assign n102 = n101 ^ n9 ;
  assign n103 = n102 ^ x6 ;
  assign n104 = n95 & ~n103 ;
  assign n105 = ~n94 & ~n104 ;
  assign n106 = ~x0 & ~n105 ;
  assign n107 = ~n86 & ~n106 ;
  assign y0 = ~n107 ;
endmodule
