module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 ;
  assign n13 = ~x1 & x9 ;
  assign n14 = x0 & n13 ;
  assign n16 = x5 & x8 ;
  assign n15 = x2 & x7 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = x8 ^ x5 ;
  assign n19 = x8 ^ x4 ;
  assign n20 = n19 ^ x4 ;
  assign n21 = x3 & x4 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = ~n20 & ~n22 ;
  assign n24 = n23 ^ x4 ;
  assign n25 = ~n18 & ~n24 ;
  assign n26 = x6 & n25 ;
  assign n27 = n26 ^ n17 ;
  assign n28 = n27 ^ n15 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = ~x6 & ~x7 ;
  assign n31 = ~x11 & n30 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = n32 ^ n17 ;
  assign n34 = n29 & ~n33 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = ~x6 & ~x10 ;
  assign n37 = x11 & ~n36 ;
  assign n38 = n21 & ~n37 ;
  assign n39 = ~n31 & ~n38 ;
  assign n40 = n39 ^ n17 ;
  assign n41 = ~n35 & ~n40 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = ~n17 & n42 ;
  assign n44 = n43 ^ n34 ;
  assign n45 = n44 ^ n16 ;
  assign n46 = n45 ^ n31 ;
  assign n47 = n14 & ~n46 ;
  assign y0 = n47 ;
endmodule
