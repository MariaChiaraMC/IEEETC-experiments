module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 ;
  assign n16 = ~x11 & ~x12 ;
  assign n17 = ~x5 & x7 ;
  assign n18 = x1 & ~x14 ;
  assign n19 = n17 & n18 ;
  assign n20 = x5 & ~x7 ;
  assign n21 = x14 ^ x13 ;
  assign n22 = ~n20 & ~n21 ;
  assign n23 = ~n19 & ~n22 ;
  assign n24 = n16 & ~n23 ;
  assign n25 = ~x13 & x14 ;
  assign n26 = ~x12 & ~n25 ;
  assign n27 = x10 & ~n26 ;
  assign n28 = ~x11 & x12 ;
  assign n29 = x12 & ~x13 ;
  assign n30 = x2 & n29 ;
  assign n31 = ~n28 & ~n30 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = x5 & x6 ;
  assign n34 = x1 & x5 ;
  assign n35 = ~n33 & ~n34 ;
  assign n36 = n35 ^ x13 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = n35 ^ n19 ;
  assign n39 = n37 & ~n38 ;
  assign n40 = n39 ^ n35 ;
  assign n41 = n40 ^ n27 ;
  assign n42 = n32 & ~n41 ;
  assign n43 = n42 ^ n39 ;
  assign n44 = n43 ^ n35 ;
  assign n45 = n44 ^ n31 ;
  assign n46 = n27 & ~n45 ;
  assign n47 = n46 ^ n27 ;
  assign n48 = ~n24 & ~n47 ;
  assign n49 = ~x0 & ~n48 ;
  assign n50 = n16 & n33 ;
  assign n51 = ~n21 & n50 ;
  assign n52 = x7 & n51 ;
  assign n53 = ~n49 & ~n52 ;
  assign n56 = n53 ^ x5 ;
  assign n57 = n56 ^ n53 ;
  assign n54 = n53 ^ x14 ;
  assign n55 = n54 ^ n53 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = ~x6 & n28 ;
  assign n60 = x8 ^ x7 ;
  assign n61 = x13 ^ x8 ;
  assign n62 = n60 & ~n61 ;
  assign n63 = n59 & n62 ;
  assign n64 = n63 ^ n53 ;
  assign n65 = n64 ^ n53 ;
  assign n66 = n65 ^ n57 ;
  assign n67 = ~n57 & ~n66 ;
  assign n68 = n67 ^ n57 ;
  assign n69 = ~n58 & ~n68 ;
  assign n70 = n69 ^ n67 ;
  assign n71 = n70 ^ n53 ;
  assign n72 = n71 ^ n57 ;
  assign n73 = ~x4 & n72 ;
  assign n74 = n73 ^ n53 ;
  assign n75 = ~x9 & ~n74 ;
  assign n76 = ~x4 & ~x5 ;
  assign n77 = x6 & ~x7 ;
  assign n78 = n76 & n77 ;
  assign n79 = x11 & ~x12 ;
  assign n80 = x9 & x10 ;
  assign n81 = n79 & n80 ;
  assign n82 = ~x0 & ~x13 ;
  assign n83 = ~x8 & n82 ;
  assign n84 = n81 & n83 ;
  assign n85 = n78 & n84 ;
  assign n86 = ~n75 & ~n85 ;
  assign n87 = x3 & ~n86 ;
  assign n88 = x12 ^ x11 ;
  assign n89 = n88 ^ x0 ;
  assign n90 = n89 ^ x12 ;
  assign n91 = n90 ^ n89 ;
  assign n92 = n89 ^ n25 ;
  assign n93 = n92 ^ n88 ;
  assign n94 = ~n91 & ~n93 ;
  assign n95 = n94 ^ n25 ;
  assign n96 = x1 & n25 ;
  assign n97 = n96 ^ n88 ;
  assign n98 = n95 & n97 ;
  assign n99 = n98 ^ n96 ;
  assign n100 = n88 & n99 ;
  assign n101 = n100 ^ n94 ;
  assign n102 = n101 ^ x11 ;
  assign n103 = n102 ^ n25 ;
  assign n104 = ~n82 & n103 ;
  assign n105 = ~x3 & x11 ;
  assign n106 = x14 & ~n77 ;
  assign n107 = n105 & n106 ;
  assign n108 = n29 & ~n107 ;
  assign n109 = x9 & ~n108 ;
  assign n110 = ~n104 & n109 ;
  assign n111 = x4 & x12 ;
  assign n112 = ~x3 & x14 ;
  assign n113 = ~n111 & n112 ;
  assign n114 = ~x11 & ~n113 ;
  assign n115 = x12 ^ x9 ;
  assign n116 = x11 ^ x3 ;
  assign n117 = n116 ^ x3 ;
  assign n118 = x1 & x13 ;
  assign n119 = n118 ^ x3 ;
  assign n120 = ~n117 & n119 ;
  assign n121 = n120 ^ x3 ;
  assign n122 = n121 ^ x12 ;
  assign n123 = n115 & n122 ;
  assign n124 = n123 ^ n120 ;
  assign n125 = n124 ^ x3 ;
  assign n126 = n125 ^ x9 ;
  assign n127 = ~x12 & n126 ;
  assign n128 = n127 ^ x12 ;
  assign n129 = n128 ^ x9 ;
  assign n130 = ~n114 & n129 ;
  assign n131 = ~n110 & ~n130 ;
  assign n132 = ~x10 & n131 ;
  assign n133 = ~n87 & ~n132 ;
  assign y0 = ~n133 ;
endmodule
