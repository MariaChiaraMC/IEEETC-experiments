module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n10 = x7 & x8 ;
  assign n11 = x4 & ~x5 ;
  assign n12 = x1 & ~n11 ;
  assign n13 = n10 & ~n12 ;
  assign n14 = ~x6 & n13 ;
  assign n15 = x3 & ~n14 ;
  assign n16 = ~x0 & ~n15 ;
  assign n17 = x4 & ~x8 ;
  assign n18 = n17 ^ x2 ;
  assign n19 = x3 ^ x1 ;
  assign n20 = n11 ^ x3 ;
  assign n21 = n20 ^ n11 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n10 ^ x6 ;
  assign n24 = ~n10 & ~n23 ;
  assign n25 = n24 ^ n11 ;
  assign n26 = n25 ^ n10 ;
  assign n27 = ~n22 & ~n26 ;
  assign n28 = n27 ^ n24 ;
  assign n29 = n28 ^ n10 ;
  assign n30 = n19 & ~n29 ;
  assign n31 = n30 ^ x3 ;
  assign n32 = ~n18 & n31 ;
  assign n33 = n16 & n32 ;
  assign y0 = n33 ;
endmodule
