module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 ;
  assign n9 = ~x0 & ~x2 ;
  assign n10 = x1 & n9 ;
  assign n12 = x7 ^ x5 ;
  assign n11 = x7 ^ x3 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n14 ^ x7 ;
  assign n16 = x7 ^ x6 ;
  assign n17 = x4 & ~n16 ;
  assign n18 = n12 ^ x7 ;
  assign n19 = n14 & ~n18 ;
  assign n20 = n19 ^ n15 ;
  assign n21 = n17 & n20 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n15 & n22 ;
  assign n24 = n23 ^ n19 ;
  assign n25 = n10 & n24 ;
  assign y0 = n25 ;
endmodule
