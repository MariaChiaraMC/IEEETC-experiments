module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 ;
  assign n30 = x1 & ~x5 ;
  assign n31 = x2 & n30 ;
  assign n32 = ~x2 & ~n30 ;
  assign n33 = ~n31 & ~n32 ;
  assign n11 = x3 ^ x0 ;
  assign n9 = x5 ^ x3 ;
  assign n18 = n11 ^ n9 ;
  assign n7 = x3 ^ x2 ;
  assign n8 = n7 ^ x5 ;
  assign n10 = n9 ^ n8 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = n9 ^ x1 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = n14 ^ n8 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = n12 & n16 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = n19 ^ n12 ;
  assign n21 = n11 ^ x5 ;
  assign n22 = n21 ^ n11 ;
  assign n23 = n17 ^ n12 ;
  assign n24 = n22 & n23 ;
  assign n25 = n24 ^ n11 ;
  assign n26 = n20 & ~n25 ;
  assign n27 = n26 ^ n11 ;
  assign n28 = n27 ^ n7 ;
  assign n29 = n28 ^ n11 ;
  assign n34 = n33 ^ n29 ;
  assign n35 = n34 ^ x4 ;
  assign n44 = n35 ^ n34 ;
  assign n36 = ~x0 & ~x1 ;
  assign n37 = ~x5 & n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = n38 ^ n34 ;
  assign n40 = n37 ^ n33 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = ~n39 & ~n42 ;
  assign n45 = n44 ^ n43 ;
  assign n46 = n45 ^ n39 ;
  assign n47 = x0 & ~x5 ;
  assign n48 = ~x3 & ~n47 ;
  assign n49 = n48 ^ n34 ;
  assign n50 = n43 ^ n39 ;
  assign n51 = n49 & ~n50 ;
  assign n52 = n51 ^ n34 ;
  assign n53 = ~n46 & n52 ;
  assign n54 = n53 ^ n34 ;
  assign n55 = n54 ^ n33 ;
  assign n56 = n55 ^ n34 ;
  assign y0 = n56 ;
endmodule
