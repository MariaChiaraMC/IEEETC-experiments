module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 ;
  assign n9 = ~x1 & x2 ;
  assign n10 = ~x6 & x7 ;
  assign n11 = x3 & n10 ;
  assign n12 = ~x5 & n11 ;
  assign n13 = n9 & n12 ;
  assign n14 = ~x0 & n13 ;
  assign n116 = x2 & ~x6 ;
  assign n117 = x1 & x5 ;
  assign n19 = ~x6 & ~x7 ;
  assign n118 = x2 & x3 ;
  assign n119 = ~n19 & ~n118 ;
  assign n120 = n117 & ~n119 ;
  assign n121 = x6 & ~x7 ;
  assign n49 = ~x1 & ~x2 ;
  assign n122 = ~x3 & ~x5 ;
  assign n123 = ~n49 & n122 ;
  assign n124 = ~n121 & n123 ;
  assign n125 = ~n120 & ~n124 ;
  assign n126 = ~n116 & ~n125 ;
  assign n85 = x3 ^ x1 ;
  assign n127 = n85 ^ x5 ;
  assign n77 = x3 ^ x2 ;
  assign n128 = x7 ^ x3 ;
  assign n129 = n128 ^ n77 ;
  assign n130 = ~n77 & n129 ;
  assign n131 = n130 ^ x3 ;
  assign n132 = n131 ^ n77 ;
  assign n133 = n127 & ~n132 ;
  assign n134 = n133 ^ n130 ;
  assign n135 = n134 ^ n77 ;
  assign n136 = ~x5 & ~n135 ;
  assign n137 = ~x6 & n136 ;
  assign n138 = ~n126 & ~n137 ;
  assign n73 = x7 ^ x5 ;
  assign n68 = x5 ^ x3 ;
  assign n69 = n68 ^ x7 ;
  assign n70 = n69 ^ x6 ;
  assign n71 = n70 ^ x7 ;
  assign n72 = n71 ^ n69 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = n74 ^ n69 ;
  assign n76 = n75 ^ n72 ;
  assign n78 = n77 ^ x5 ;
  assign n79 = n78 ^ x7 ;
  assign n80 = n79 ^ n75 ;
  assign n81 = ~n76 & ~n80 ;
  assign n82 = n81 ^ n72 ;
  assign n83 = n82 ^ n69 ;
  assign n84 = n83 ^ n79 ;
  assign n86 = n85 ^ x6 ;
  assign n87 = n86 ^ x7 ;
  assign n88 = n87 ^ x7 ;
  assign n89 = n88 ^ n71 ;
  assign n90 = n89 ^ n87 ;
  assign n91 = n90 ^ n79 ;
  assign n92 = n91 ^ n72 ;
  assign n93 = n92 ^ n69 ;
  assign n94 = n93 ^ n87 ;
  assign n95 = n94 ^ n79 ;
  assign n96 = n94 & ~n95 ;
  assign n97 = n96 ^ n87 ;
  assign n98 = n97 ^ n79 ;
  assign n99 = n91 ^ n76 ;
  assign n100 = n92 ^ n87 ;
  assign n101 = n100 ^ n79 ;
  assign n102 = ~n99 & n101 ;
  assign n103 = n102 ^ n75 ;
  assign n104 = n103 ^ n91 ;
  assign n105 = n104 ^ n69 ;
  assign n106 = n105 ^ n87 ;
  assign n107 = ~n98 & ~n106 ;
  assign n108 = n107 ^ n87 ;
  assign n109 = ~n84 & n108 ;
  assign n110 = n109 ^ n81 ;
  assign n111 = n110 ^ n107 ;
  assign n112 = n111 ^ n72 ;
  assign n113 = n112 ^ n69 ;
  assign n114 = n113 ^ n87 ;
  assign n115 = n114 ^ n79 ;
  assign n139 = n138 ^ n115 ;
  assign n140 = ~x0 & ~n139 ;
  assign n141 = n140 ^ n115 ;
  assign n142 = ~n13 & ~n141 ;
  assign n15 = x0 & x3 ;
  assign n16 = x5 & x7 ;
  assign n17 = n9 & n16 ;
  assign n18 = n15 & n17 ;
  assign n20 = x1 & x2 ;
  assign n23 = x3 & ~x7 ;
  assign n24 = x0 & n10 ;
  assign n25 = ~n23 & ~n24 ;
  assign n26 = ~n15 & ~n25 ;
  assign n27 = n20 & n26 ;
  assign n28 = ~x2 & ~x7 ;
  assign n29 = n28 ^ x3 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = n28 ^ x7 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = ~n30 & n32 ;
  assign n34 = n33 ^ n28 ;
  assign n35 = ~x1 & n34 ;
  assign n36 = n35 ^ n28 ;
  assign n37 = n36 ^ x0 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = ~x1 & x7 ;
  assign n40 = ~n23 & ~n39 ;
  assign n41 = ~x2 & ~n40 ;
  assign n42 = n41 ^ n36 ;
  assign n43 = ~n38 & n42 ;
  assign n44 = n43 ^ n36 ;
  assign n45 = x6 & n44 ;
  assign n46 = ~n27 & ~n45 ;
  assign n21 = n19 & ~n20 ;
  assign n22 = ~x3 & n21 ;
  assign n47 = n46 ^ n22 ;
  assign n48 = n47 ^ x5 ;
  assign n56 = n48 ^ n47 ;
  assign n50 = n49 ^ n48 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = n49 ^ n22 ;
  assign n53 = n52 ^ n49 ;
  assign n54 = n53 ^ n51 ;
  assign n55 = n51 & n54 ;
  assign n57 = n56 ^ n55 ;
  assign n58 = n57 ^ n51 ;
  assign n59 = n47 ^ x0 ;
  assign n60 = n55 ^ n51 ;
  assign n61 = ~n59 & n60 ;
  assign n62 = n61 ^ n47 ;
  assign n63 = ~n58 & ~n62 ;
  assign n64 = n63 ^ n47 ;
  assign n65 = n64 ^ n22 ;
  assign n66 = n65 ^ n47 ;
  assign n67 = ~n18 & ~n66 ;
  assign n143 = n142 ^ n67 ;
  assign n144 = ~x4 & n143 ;
  assign n145 = n144 ^ n142 ;
  assign n146 = ~n14 & n145 ;
  assign y0 = ~n146 ;
endmodule
