module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 ;
  assign n47 = x3 ^ x0 ;
  assign n48 = x5 ^ x3 ;
  assign n49 = n48 ^ x5 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = x7 ^ x5 ;
  assign n52 = x6 ^ x5 ;
  assign n53 = ~x4 & ~n52 ;
  assign n54 = n53 ^ n47 ;
  assign n55 = ~n51 & ~n54 ;
  assign n56 = n55 ^ x5 ;
  assign n57 = n50 & n56 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = ~n47 & n58 ;
  assign n60 = n59 ^ n55 ;
  assign n61 = n60 ^ n57 ;
  assign n62 = n61 ^ n47 ;
  assign n15 = x5 & x7 ;
  assign n16 = x1 & n15 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = ~x6 & ~n17 ;
  assign n25 = x1 & ~x5 ;
  assign n26 = ~x4 & ~n25 ;
  assign n27 = x0 & ~n26 ;
  assign n28 = ~x8 & n27 ;
  assign n19 = ~x3 & x8 ;
  assign n20 = ~x4 & ~x6 ;
  assign n21 = ~x0 & n20 ;
  assign n22 = n19 & n21 ;
  assign n23 = n22 ^ x1 ;
  assign n24 = n23 ^ x3 ;
  assign n29 = n28 ^ n24 ;
  assign n30 = n29 ^ n24 ;
  assign n31 = n24 ^ n23 ;
  assign n32 = n31 ^ x1 ;
  assign n33 = n30 & n32 ;
  assign n34 = n33 ^ n23 ;
  assign n35 = ~x5 & ~x7 ;
  assign n36 = ~n23 & n35 ;
  assign n37 = n36 ^ x1 ;
  assign n38 = ~n34 & ~n37 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = ~x1 & n39 ;
  assign n41 = n40 ^ n33 ;
  assign n42 = n41 ^ n22 ;
  assign n43 = n42 ^ n23 ;
  assign n44 = ~n18 & ~n43 ;
  assign n63 = n62 ^ n44 ;
  assign n64 = n63 ^ n44 ;
  assign n45 = n44 ^ x8 ;
  assign n46 = n45 ^ n44 ;
  assign n65 = n64 ^ n46 ;
  assign n66 = n44 ^ x1 ;
  assign n67 = n66 ^ n44 ;
  assign n68 = n67 ^ n64 ;
  assign n69 = n64 & n68 ;
  assign n70 = n69 ^ n64 ;
  assign n71 = ~n65 & n70 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = n72 ^ n44 ;
  assign n74 = n73 ^ n64 ;
  assign n75 = x2 & n74 ;
  assign n76 = n75 ^ n44 ;
  assign n12 = ~x8 & x10 ;
  assign n13 = x3 ^ x2 ;
  assign n14 = n12 & n13 ;
  assign n77 = n76 ^ n14 ;
  assign n78 = x9 & n77 ;
  assign n79 = n78 ^ n76 ;
  assign y0 = n79 ;
endmodule
