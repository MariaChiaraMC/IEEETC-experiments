module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n10 = x7 ^ x3 ;
  assign n11 = n10 ^ x8 ;
  assign n12 = n11 ^ x1 ;
  assign n13 = x4 & ~x5 ;
  assign n14 = n13 ^ x3 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = x8 & n15 ;
  assign n17 = n16 ^ x3 ;
  assign n18 = n17 ^ x8 ;
  assign n19 = n18 ^ n11 ;
  assign n20 = n19 ^ x1 ;
  assign n21 = n12 & ~n20 ;
  assign n22 = n21 ^ n16 ;
  assign n23 = n22 ^ x3 ;
  assign n24 = n23 ^ n11 ;
  assign n25 = ~x1 & n24 ;
  assign n26 = n25 ^ x1 ;
  assign n27 = n26 ^ x1 ;
  assign n28 = ~x2 & n27 ;
  assign n29 = ~x0 & ~n28 ;
  assign n30 = x6 ^ x0 ;
  assign n31 = x6 ^ x4 ;
  assign n32 = n31 ^ x4 ;
  assign n33 = x5 ^ x4 ;
  assign n34 = ~n32 & n33 ;
  assign n35 = n34 ^ x4 ;
  assign n36 = n30 & n35 ;
  assign n37 = n36 ^ x0 ;
  assign n38 = ~n29 & ~n37 ;
  assign y0 = n38 ;
endmodule
