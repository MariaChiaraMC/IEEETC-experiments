module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n10 = ~x2 & ~x5 ;
  assign n11 = x1 & x3 ;
  assign n12 = x0 & n11 ;
  assign n13 = n10 & n12 ;
  assign n14 = x6 ^ x4 ;
  assign n19 = n14 ^ x4 ;
  assign n16 = x8 ^ x4 ;
  assign n15 = n14 ^ x7 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n17 ^ x4 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = n15 ^ n14 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = n22 ^ x4 ;
  assign n24 = n17 & ~n23 ;
  assign n25 = n24 ^ n17 ;
  assign n26 = ~n22 & n25 ;
  assign n27 = n26 ^ x4 ;
  assign n28 = n20 & n27 ;
  assign n29 = n28 ^ n24 ;
  assign n30 = n29 ^ x4 ;
  assign n31 = n30 ^ n19 ;
  assign n32 = n13 & n31 ;
  assign y0 = n32 ;
endmodule
