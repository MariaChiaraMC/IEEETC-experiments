module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 ;
  assign n17 = ~x8 & ~x12 ;
  assign n18 = ~x11 & n17 ;
  assign n19 = x10 ^ x9 ;
  assign n20 = n18 & n19 ;
  assign n21 = ~x14 & ~x15 ;
  assign n22 = n21 ^ x13 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = x15 ^ x14 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = ~n23 & n25 ;
  assign n27 = n26 ^ n21 ;
  assign n28 = n20 & n27 ;
  assign n29 = n28 ^ x5 ;
  assign n30 = n28 ^ x7 ;
  assign n31 = n30 ^ x7 ;
  assign n32 = x7 ^ x6 ;
  assign n33 = n31 & ~n32 ;
  assign n34 = n33 ^ x7 ;
  assign n35 = x4 & ~x7 ;
  assign n36 = n35 ^ n29 ;
  assign n37 = ~n34 & ~n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = ~n29 & n38 ;
  assign n40 = n39 ^ n28 ;
  assign n41 = n40 ^ n29 ;
  assign n42 = ~x0 & n41 ;
  assign y0 = ~n42 ;
endmodule
