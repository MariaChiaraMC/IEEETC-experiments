module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 ;
  assign n8 = x5 & x6 ;
  assign n9 = ~x1 & ~n8 ;
  assign n10 = x5 & ~x6 ;
  assign n11 = x4 & ~n10 ;
  assign n12 = x3 & ~n11 ;
  assign n13 = ~n9 & n12 ;
  assign n14 = x1 & x2 ;
  assign n18 = x4 & ~x6 ;
  assign n15 = x2 & ~x4 ;
  assign n16 = n15 ^ x3 ;
  assign n17 = x6 & n16 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = ~n14 & n19 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = ~x5 & n21 ;
  assign n23 = ~x3 & n10 ;
  assign n24 = ~x2 & x4 ;
  assign n25 = ~n23 & ~n24 ;
  assign n26 = ~x1 & ~n25 ;
  assign n27 = x4 & x6 ;
  assign n28 = ~x3 & x5 ;
  assign n29 = n27 & n28 ;
  assign n30 = ~n26 & ~n29 ;
  assign n31 = ~n22 & n30 ;
  assign n32 = ~n13 & n31 ;
  assign n33 = x0 & ~n32 ;
  assign n34 = ~x4 & n28 ;
  assign n35 = ~x0 & x6 ;
  assign n36 = ~x5 & n35 ;
  assign n37 = ~n34 & ~n36 ;
  assign n38 = n14 & ~n37 ;
  assign n39 = ~x4 & x6 ;
  assign n40 = ~x0 & n39 ;
  assign n41 = ~x1 & n18 ;
  assign n42 = ~n40 & ~n41 ;
  assign n43 = n28 & ~n42 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = x4 ^ x3 ;
  assign n46 = n45 ^ x5 ;
  assign n47 = n46 ^ x4 ;
  assign n48 = n47 ^ x5 ;
  assign n49 = n48 ^ x0 ;
  assign n52 = n46 ^ x5 ;
  assign n50 = n46 ^ x6 ;
  assign n51 = n50 ^ x0 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n52 ^ n48 ;
  assign n55 = n54 ^ x0 ;
  assign n56 = n55 ^ n46 ;
  assign n57 = n56 ^ n49 ;
  assign n58 = n53 & ~n57 ;
  assign n59 = n58 ^ x0 ;
  assign n60 = ~n49 & ~n59 ;
  assign n61 = n60 ^ x0 ;
  assign n62 = n46 ^ x1 ;
  assign n63 = n58 ^ n53 ;
  assign n64 = ~n62 & n63 ;
  assign n65 = n64 ^ n46 ;
  assign n66 = ~n61 & n65 ;
  assign n67 = n66 ^ x2 ;
  assign n68 = n67 ^ n66 ;
  assign n69 = n39 ^ x0 ;
  assign n70 = n69 ^ n39 ;
  assign n76 = n70 ^ n69 ;
  assign n73 = n69 ^ x3 ;
  assign n77 = n76 ^ n73 ;
  assign n78 = n77 ^ n73 ;
  assign n79 = n69 ^ x1 ;
  assign n80 = n79 ^ n73 ;
  assign n81 = n78 & ~n80 ;
  assign n71 = n69 ^ n18 ;
  assign n72 = n71 ^ n70 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = ~n70 & ~n74 ;
  assign n82 = n81 ^ n75 ;
  assign n83 = n82 ^ n70 ;
  assign n84 = n75 ^ n73 ;
  assign n85 = n84 ^ n77 ;
  assign n86 = n73 & n85 ;
  assign n87 = n86 ^ n75 ;
  assign n88 = ~n83 & n87 ;
  assign n89 = n88 ^ n81 ;
  assign n90 = n89 ^ n86 ;
  assign n91 = n90 ^ n70 ;
  assign n92 = n91 ^ n73 ;
  assign n93 = n92 ^ n77 ;
  assign n94 = n93 ^ x0 ;
  assign n95 = ~x5 & n94 ;
  assign n96 = ~n18 & ~n23 ;
  assign n97 = ~x1 & ~n96 ;
  assign n98 = ~n95 & ~n97 ;
  assign n99 = n98 ^ n66 ;
  assign n100 = ~n68 & ~n99 ;
  assign n101 = n100 ^ n66 ;
  assign n102 = n101 ^ n38 ;
  assign n103 = n44 & n102 ;
  assign n104 = n103 ^ n100 ;
  assign n105 = n104 ^ n66 ;
  assign n106 = n105 ^ n43 ;
  assign n107 = ~n38 & n106 ;
  assign n108 = n107 ^ n38 ;
  assign n109 = ~n33 & ~n108 ;
  assign y0 = ~n109 ;
endmodule
