module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 ;
  output y0 ;
  wire n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 ;
  assign n21 = x2 & x10 ;
  assign n27 = ~x14 & x15 ;
  assign n28 = x7 ^ x6 ;
  assign n29 = x3 & n28 ;
  assign n30 = n29 ^ x6 ;
  assign n31 = ~n27 & n30 ;
  assign n32 = ~x3 & x13 ;
  assign n33 = x11 & n32 ;
  assign n34 = x4 & ~n33 ;
  assign n35 = n27 ^ x12 ;
  assign n36 = n35 ^ n27 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = x11 & x13 ;
  assign n39 = x14 & ~n38 ;
  assign n40 = ~x15 & ~n39 ;
  assign n41 = n40 ^ n32 ;
  assign n42 = ~n32 & n41 ;
  assign n43 = n42 ^ n27 ;
  assign n44 = n43 ^ n32 ;
  assign n45 = n37 & ~n44 ;
  assign n46 = n45 ^ n42 ;
  assign n47 = n46 ^ n32 ;
  assign n48 = n34 & ~n47 ;
  assign n49 = n48 ^ n34 ;
  assign n50 = ~n31 & ~n49 ;
  assign n22 = x0 & x3 ;
  assign n23 = x9 & n22 ;
  assign n24 = x8 & n23 ;
  assign n51 = n50 ^ n24 ;
  assign n52 = n51 ^ n24 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = n25 ^ n24 ;
  assign n53 = n52 ^ n26 ;
  assign n54 = n24 ^ x0 ;
  assign n55 = n54 ^ n24 ;
  assign n56 = n55 ^ n52 ;
  assign n57 = ~n52 & n56 ;
  assign n58 = n57 ^ n52 ;
  assign n59 = ~n53 & ~n58 ;
  assign n60 = n59 ^ n57 ;
  assign n61 = n60 ^ n24 ;
  assign n62 = n61 ^ n52 ;
  assign n63 = x1 & ~n62 ;
  assign n64 = n63 ^ n24 ;
  assign n65 = n21 & n64 ;
  assign n66 = ~x10 & x18 ;
  assign n67 = x16 & n66 ;
  assign n68 = x19 ^ x17 ;
  assign n69 = n67 & n68 ;
  assign n70 = ~n65 & ~n69 ;
  assign y0 = ~n70 ;
endmodule
