module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
  assign n11 = ~x5 & ~x9 ;
  assign n12 = ~x8 & ~n11 ;
  assign n13 = x4 & x6 ;
  assign n14 = ~x1 & ~x3 ;
  assign n15 = ~x2 & n14 ;
  assign n16 = n13 & n15 ;
  assign n17 = ~n12 & n16 ;
  assign n18 = n17 ^ x0 ;
  assign n26 = n18 ^ n17 ;
  assign n19 = ~x2 & x7 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n19 ^ x8 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n21 & ~n24 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = n17 ^ x4 ;
  assign n30 = n25 ^ n21 ;
  assign n31 = ~n29 & n30 ;
  assign n32 = n31 ^ n17 ;
  assign n33 = ~n28 & n32 ;
  assign n34 = n33 ^ n17 ;
  assign n35 = n34 ^ n17 ;
  assign y0 = n35 ;
endmodule
