module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 ;
  assign n17 = x12 ^ x11 ;
  assign n15 = x10 ^ x0 ;
  assign n16 = n15 ^ x9 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = n15 ^ x10 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = n21 ^ n15 ;
  assign n24 = n22 ^ n15 ;
  assign n23 = n22 ^ n16 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n18 & ~n25 ;
  assign n27 = n26 ^ n22 ;
  assign n28 = n27 ^ n24 ;
  assign n29 = n15 ^ x12 ;
  assign n30 = n29 ^ n16 ;
  assign n31 = n30 ^ n20 ;
  assign n32 = n31 ^ n22 ;
  assign n33 = n32 ^ n24 ;
  assign n34 = n31 ^ n17 ;
  assign n35 = n34 ^ n24 ;
  assign n36 = n33 & n35 ;
  assign n37 = n36 ^ n22 ;
  assign n38 = n37 ^ n16 ;
  assign n39 = n38 ^ n31 ;
  assign n40 = n39 ^ n24 ;
  assign n41 = n31 ^ n23 ;
  assign n42 = n41 ^ n24 ;
  assign n43 = ~x13 & ~n42 ;
  assign n44 = n43 ^ x13 ;
  assign n45 = n44 ^ n16 ;
  assign n46 = n45 ^ n31 ;
  assign n47 = n46 ^ n24 ;
  assign n48 = ~n40 & ~n47 ;
  assign n49 = n48 ^ n16 ;
  assign n50 = n49 ^ n24 ;
  assign n51 = n28 & n50 ;
  assign n52 = n51 ^ n48 ;
  assign n53 = n52 ^ n16 ;
  assign n54 = n53 ^ n24 ;
  assign n55 = n54 ^ x10 ;
  assign n56 = x13 ^ x9 ;
  assign n57 = n56 ^ x9 ;
  assign n58 = ~x11 & ~x12 ;
  assign n59 = n58 ^ x0 ;
  assign n60 = n59 ^ x0 ;
  assign n61 = x9 ^ x0 ;
  assign n62 = n61 ^ x0 ;
  assign n63 = n60 & ~n62 ;
  assign n64 = n63 ^ x0 ;
  assign n65 = ~x10 & n64 ;
  assign n66 = n65 ^ x0 ;
  assign n67 = n66 ^ x9 ;
  assign n68 = ~n57 & n67 ;
  assign n69 = n68 ^ x9 ;
  assign n70 = x9 & x11 ;
  assign n71 = n70 ^ n55 ;
  assign n72 = n69 & ~n71 ;
  assign n73 = n72 ^ n70 ;
  assign n74 = ~n55 & n73 ;
  assign n75 = n74 ^ n55 ;
  assign y0 = ~n75 ;
endmodule
