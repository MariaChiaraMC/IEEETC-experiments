module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 ;
  assign n13 = x5 ^ x1 ;
  assign n14 = x5 ^ x3 ;
  assign n22 = n14 ^ x5 ;
  assign n23 = n22 ^ x5 ;
  assign n24 = n22 & ~n23 ;
  assign n15 = n14 ^ x4 ;
  assign n16 = n15 ^ x0 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n15 ^ n14 ;
  assign n19 = n18 ^ x5 ;
  assign n20 = n17 & ~n19 ;
  assign n27 = n24 ^ n20 ;
  assign n21 = n20 ^ n13 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = ~n21 & n25 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = ~n13 & n28 ;
  assign n30 = n29 ^ n20 ;
  assign n31 = n30 ^ n24 ;
  assign n32 = n31 ^ n26 ;
  assign n33 = n32 ^ x3 ;
  assign n34 = x2 & n33 ;
  assign n35 = ~x4 & ~x5 ;
  assign n8 = ~x2 & x4 ;
  assign n9 = ~x1 & n8 ;
  assign n36 = n35 ^ n9 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = ~x0 & ~x1 ;
  assign n39 = x2 & ~n38 ;
  assign n40 = x5 & ~n39 ;
  assign n41 = n40 ^ n35 ;
  assign n42 = n41 ^ n35 ;
  assign n43 = ~n37 & ~n42 ;
  assign n44 = n43 ^ n35 ;
  assign n45 = ~x3 & ~n44 ;
  assign n46 = n45 ^ n35 ;
  assign n47 = ~n34 & ~n46 ;
  assign n10 = x4 ^ x3 ;
  assign n11 = ~n9 & ~n10 ;
  assign n12 = x5 & ~n11 ;
  assign n48 = n47 ^ n12 ;
  assign n49 = ~x6 & ~n48 ;
  assign n50 = n49 ^ n47 ;
  assign y0 = ~n50 ;
endmodule
