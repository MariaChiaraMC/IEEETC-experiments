module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 ;
  assign n9 = x0 & x4 ;
  assign n10 = ~x0 & ~x4 ;
  assign n11 = ~n9 & ~n10 ;
  assign n12 = x3 ^ x1 ;
  assign n13 = x5 ^ x3 ;
  assign n14 = n12 & n13 ;
  assign n15 = n13 ^ x7 ;
  assign n16 = ~x2 & ~x6 ;
  assign n17 = x2 & x6 ;
  assign n18 = ~n16 & ~n17 ;
  assign n19 = x5 & n18 ;
  assign n20 = n19 ^ n14 ;
  assign n21 = ~n15 & n20 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n14 & n22 ;
  assign n24 = n11 & n23 ;
  assign n25 = ~x3 & x5 ;
  assign n26 = x2 & x7 ;
  assign n27 = n26 ^ x4 ;
  assign n28 = ~x1 & ~n27 ;
  assign n29 = n28 ^ x4 ;
  assign n30 = n29 ^ x0 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = x1 & ~x2 ;
  assign n33 = x1 & x4 ;
  assign n34 = ~x2 & x7 ;
  assign n35 = ~n33 & ~n34 ;
  assign n36 = ~n32 & ~n35 ;
  assign n37 = n36 ^ n29 ;
  assign n38 = n31 & ~n37 ;
  assign n39 = n38 ^ n29 ;
  assign n40 = n25 & ~n39 ;
  assign n41 = ~n24 & ~n40 ;
  assign n42 = ~x3 & ~x7 ;
  assign n43 = x4 ^ x0 ;
  assign n44 = x6 ^ x2 ;
  assign n45 = x1 & ~x5 ;
  assign n46 = n45 ^ x6 ;
  assign n47 = n46 ^ n45 ;
  assign n48 = ~x1 & x5 ;
  assign n49 = n48 ^ n45 ;
  assign n50 = ~n47 & n49 ;
  assign n51 = n50 ^ n45 ;
  assign n52 = n44 & n51 ;
  assign n53 = n52 ^ x4 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = x5 ^ x1 ;
  assign n56 = ~x2 & x6 ;
  assign n57 = n56 ^ x5 ;
  assign n58 = n57 ^ n56 ;
  assign n59 = x2 & ~x6 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = ~n58 & n60 ;
  assign n62 = n61 ^ n56 ;
  assign n63 = n55 & n62 ;
  assign n64 = n63 ^ n52 ;
  assign n65 = n54 & n64 ;
  assign n66 = n65 ^ n52 ;
  assign n67 = n43 & n66 ;
  assign n68 = ~n42 & n67 ;
  assign n69 = ~x2 & x4 ;
  assign n70 = x0 & x1 ;
  assign n71 = n69 & n70 ;
  assign n72 = x5 & n71 ;
  assign n73 = ~n68 & ~n72 ;
  assign n74 = n41 & n73 ;
  assign n75 = n17 & n33 ;
  assign n76 = x7 & n75 ;
  assign n77 = x2 & ~x4 ;
  assign n78 = ~x1 & n77 ;
  assign n79 = n78 ^ x2 ;
  assign n80 = x5 & n79 ;
  assign n81 = ~n32 & ~n80 ;
  assign n82 = ~n76 & n81 ;
  assign n83 = ~x0 & ~n82 ;
  assign n86 = ~x0 & x4 ;
  assign n84 = x4 ^ x2 ;
  assign n85 = n84 ^ x7 ;
  assign n87 = n86 ^ n85 ;
  assign n96 = n87 ^ n85 ;
  assign n88 = x0 & ~x4 ;
  assign n89 = n17 & n88 ;
  assign n90 = n89 ^ n87 ;
  assign n91 = n90 ^ n85 ;
  assign n92 = n87 ^ n84 ;
  assign n93 = n92 ^ n89 ;
  assign n94 = n93 ^ n91 ;
  assign n95 = n91 & ~n94 ;
  assign n97 = n96 ^ n95 ;
  assign n98 = n97 ^ n91 ;
  assign n99 = n85 ^ n16 ;
  assign n100 = n95 ^ n91 ;
  assign n101 = n99 & n100 ;
  assign n102 = n101 ^ n85 ;
  assign n103 = ~n98 & ~n102 ;
  assign n104 = n103 ^ n85 ;
  assign n105 = n104 ^ x7 ;
  assign n106 = n105 ^ n85 ;
  assign n107 = n48 & n106 ;
  assign n108 = ~x5 & x7 ;
  assign n109 = ~x1 & n108 ;
  assign n110 = ~n18 & n109 ;
  assign n111 = ~n11 & n110 ;
  assign n112 = ~x6 & x7 ;
  assign n113 = ~x2 & ~x5 ;
  assign n114 = ~n112 & n113 ;
  assign n115 = n70 & ~n114 ;
  assign n116 = ~n69 & n115 ;
  assign n117 = ~n111 & ~n116 ;
  assign n118 = ~n107 & n117 ;
  assign n119 = ~n83 & n118 ;
  assign n120 = x3 & ~n119 ;
  assign n121 = n17 ^ n16 ;
  assign n122 = n16 ^ x4 ;
  assign n123 = n122 ^ n16 ;
  assign n124 = n121 & ~n123 ;
  assign n125 = n124 ^ n16 ;
  assign n126 = ~n43 & n125 ;
  assign n127 = x3 & n126 ;
  assign n128 = x3 ^ x2 ;
  assign n129 = n128 ^ x6 ;
  assign n130 = n129 ^ x7 ;
  assign n131 = n10 ^ n9 ;
  assign n132 = n128 ^ n9 ;
  assign n133 = n132 ^ n9 ;
  assign n134 = n131 & ~n133 ;
  assign n135 = n134 ^ n9 ;
  assign n136 = n135 ^ n129 ;
  assign n137 = ~n130 & ~n136 ;
  assign n138 = n137 ^ n134 ;
  assign n139 = n138 ^ n9 ;
  assign n140 = n139 ^ x7 ;
  assign n141 = ~n129 & n140 ;
  assign n142 = n141 ^ n129 ;
  assign n143 = ~n127 & n142 ;
  assign n144 = n143 ^ n45 ;
  assign n145 = n143 ^ n48 ;
  assign n146 = n145 ^ n48 ;
  assign n147 = n146 ^ n144 ;
  assign n148 = ~x3 & x7 ;
  assign n149 = n148 ^ n84 ;
  assign n150 = n84 & n149 ;
  assign n151 = n150 ^ n48 ;
  assign n152 = n151 ^ n84 ;
  assign n153 = ~n147 & ~n152 ;
  assign n154 = n153 ^ n150 ;
  assign n155 = n154 ^ n84 ;
  assign n156 = ~n144 & n155 ;
  assign n157 = n156 ^ n143 ;
  assign n158 = ~n120 & n157 ;
  assign n159 = n74 & n158 ;
  assign y0 = ~n159 ;
endmodule
