module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 ;
  output y0 ;
  wire n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 ;
  assign n28 = x8 ^ x7 ;
  assign n29 = x8 & ~n28 ;
  assign n30 = x6 & n29 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = x13 ^ x5 ;
  assign n33 = x0 & n32 ;
  assign n34 = n33 ^ x5 ;
  assign n35 = ~n31 & n34 ;
  assign n36 = ~x6 & ~x10 ;
  assign n37 = ~x11 & n36 ;
  assign n38 = x14 ^ x9 ;
  assign n39 = x0 & n38 ;
  assign n40 = n39 ^ x9 ;
  assign n41 = n37 & n40 ;
  assign n42 = ~x7 & ~x8 ;
  assign n43 = x15 ^ x12 ;
  assign n44 = x0 & n43 ;
  assign n45 = n44 ^ x12 ;
  assign n46 = x6 & n45 ;
  assign n47 = ~n42 & n46 ;
  assign n48 = ~n41 & ~n47 ;
  assign n49 = ~n35 & n48 ;
  assign y0 = ~n49 ;
endmodule
