module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n11 = x1 & x3 ;
  assign n12 = x0 & ~n11 ;
  assign n9 = ~x1 & ~x3 ;
  assign n10 = x2 & ~n9 ;
  assign n13 = n12 ^ n10 ;
  assign n23 = n13 ^ n12 ;
  assign n14 = x7 & ~n12 ;
  assign n15 = x6 & ~n14 ;
  assign n16 = ~x5 & ~n15 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n17 ^ n12 ;
  assign n19 = n16 ^ x4 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n18 & ~n21 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ n18 ;
  assign n26 = n12 ^ x6 ;
  assign n27 = n22 ^ n18 ;
  assign n28 = n26 & n27 ;
  assign n29 = n28 ^ n12 ;
  assign n30 = n25 & n29 ;
  assign n31 = n30 ^ n12 ;
  assign n32 = n31 ^ n12 ;
  assign y0 = ~n32 ;
endmodule
