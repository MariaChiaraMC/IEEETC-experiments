module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 ;
  assign n10 = x1 & x3 ;
  assign n11 = ~x7 & ~x8 ;
  assign n12 = ~x3 & n11 ;
  assign n13 = ~x1 & x2 ;
  assign n14 = n12 & n13 ;
  assign n15 = ~n10 & ~n14 ;
  assign n16 = ~x5 & ~n15 ;
  assign n17 = x3 & x7 ;
  assign n18 = ~x4 & x5 ;
  assign n19 = ~x2 & n18 ;
  assign n20 = ~n17 & n19 ;
  assign n21 = ~n11 & n20 ;
  assign n22 = ~n16 & ~n21 ;
  assign n23 = ~x6 & ~n22 ;
  assign n24 = x2 & x3 ;
  assign n25 = n18 & n24 ;
  assign n34 = x5 ^ x4 ;
  assign n35 = n34 ^ x4 ;
  assign n36 = x6 & ~n11 ;
  assign n37 = n36 ^ x4 ;
  assign n38 = ~n35 & n37 ;
  assign n39 = n38 ^ x4 ;
  assign n40 = x3 & n39 ;
  assign n26 = x1 & ~x2 ;
  assign n29 = x5 & x8 ;
  assign n30 = x7 & n29 ;
  assign n31 = n26 & ~n30 ;
  assign n32 = n31 ^ x4 ;
  assign n27 = ~n13 & ~n26 ;
  assign n28 = n27 ^ x4 ;
  assign n33 = n32 ^ n28 ;
  assign n41 = n40 ^ n33 ;
  assign n42 = n41 ^ n33 ;
  assign n43 = n33 ^ n28 ;
  assign n44 = n43 ^ x4 ;
  assign n45 = ~n42 & ~n44 ;
  assign n46 = n45 ^ n28 ;
  assign n47 = ~x1 & ~n28 ;
  assign n48 = n47 ^ x4 ;
  assign n49 = ~n46 & n48 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = x4 & n50 ;
  assign n52 = n51 ^ n45 ;
  assign n53 = n52 ^ n27 ;
  assign n54 = n53 ^ n28 ;
  assign n55 = ~n25 & n54 ;
  assign n56 = ~n23 & n55 ;
  assign n57 = x0 & ~n56 ;
  assign n66 = x3 ^ x2 ;
  assign n67 = ~x5 & n26 ;
  assign n68 = n67 ^ n66 ;
  assign n69 = x7 ^ x1 ;
  assign n70 = x7 ^ x3 ;
  assign n71 = n70 ^ x7 ;
  assign n72 = n69 & n71 ;
  assign n73 = n72 ^ x7 ;
  assign n74 = n73 ^ n66 ;
  assign n75 = n68 & n74 ;
  assign n76 = n75 ^ n72 ;
  assign n77 = n76 ^ x7 ;
  assign n78 = n77 ^ n67 ;
  assign n79 = ~n66 & n78 ;
  assign n80 = n79 ^ n66 ;
  assign n81 = n80 ^ n67 ;
  assign n82 = ~x0 & ~n81 ;
  assign n83 = x2 & ~x5 ;
  assign n84 = ~x1 & ~x3 ;
  assign n85 = n83 & n84 ;
  assign n58 = x2 & x5 ;
  assign n86 = x1 & ~x7 ;
  assign n87 = n58 & n86 ;
  assign n88 = x6 & n87 ;
  assign n89 = ~n85 & ~n88 ;
  assign n90 = ~n82 & n89 ;
  assign n59 = ~x0 & ~x3 ;
  assign n60 = n58 & n59 ;
  assign n61 = x5 & n27 ;
  assign n62 = n61 ^ n13 ;
  assign n63 = x3 & ~n62 ;
  assign n64 = ~n31 & n63 ;
  assign n65 = ~n60 & ~n64 ;
  assign n91 = n90 ^ n65 ;
  assign n92 = ~x4 & n91 ;
  assign n93 = n92 ^ n90 ;
  assign n94 = ~n57 & n93 ;
  assign n95 = ~x2 & x3 ;
  assign n96 = ~n17 & ~n95 ;
  assign n97 = x4 & ~x5 ;
  assign n98 = n96 & n97 ;
  assign n99 = ~x3 & x5 ;
  assign n100 = ~x8 & n19 ;
  assign n101 = ~n99 & ~n100 ;
  assign n102 = ~x0 & ~n101 ;
  assign n103 = ~x4 & n95 ;
  assign n104 = ~x7 & n103 ;
  assign n105 = ~n102 & ~n104 ;
  assign n106 = ~n98 & n105 ;
  assign n107 = ~x1 & ~n106 ;
  assign n108 = ~x2 & ~x3 ;
  assign n109 = x7 & x8 ;
  assign n110 = n24 & n109 ;
  assign n111 = ~n108 & ~n110 ;
  assign n112 = ~x0 & ~n111 ;
  assign n113 = n112 ^ x2 ;
  assign n114 = n12 ^ x5 ;
  assign n115 = n114 ^ n12 ;
  assign n116 = n12 ^ n10 ;
  assign n117 = n115 & n116 ;
  assign n118 = n117 ^ n12 ;
  assign n119 = n118 ^ n112 ;
  assign n120 = ~n113 & ~n119 ;
  assign n121 = n120 ^ n117 ;
  assign n122 = n121 ^ n12 ;
  assign n123 = n122 ^ x2 ;
  assign n124 = ~n112 & n123 ;
  assign n125 = n124 ^ n112 ;
  assign n126 = n125 ^ n112 ;
  assign n127 = x4 & ~n126 ;
  assign n128 = ~n107 & ~n127 ;
  assign n129 = n128 ^ x6 ;
  assign n130 = n129 ^ n128 ;
  assign n131 = x0 & ~n29 ;
  assign n132 = n108 & ~n131 ;
  assign n133 = ~x1 & n132 ;
  assign n134 = n59 ^ n29 ;
  assign n135 = n134 ^ x4 ;
  assign n136 = n13 ^ x2 ;
  assign n137 = n59 & ~n136 ;
  assign n138 = n137 ^ n13 ;
  assign n139 = ~n135 & n138 ;
  assign n140 = n139 ^ n137 ;
  assign n141 = n140 ^ n13 ;
  assign n142 = n141 ^ n59 ;
  assign n143 = ~x4 & n142 ;
  assign n144 = ~n133 & ~n143 ;
  assign n145 = x7 & ~n144 ;
  assign n146 = x7 & n99 ;
  assign n147 = ~x4 & ~x5 ;
  assign n148 = x8 & n147 ;
  assign n149 = ~x0 & n148 ;
  assign n150 = ~n146 & ~n149 ;
  assign n151 = x1 & x2 ;
  assign n152 = ~n150 & n151 ;
  assign n153 = x3 ^ x1 ;
  assign n154 = n18 ^ x3 ;
  assign n155 = n154 ^ n18 ;
  assign n156 = ~n19 & ~n83 ;
  assign n157 = n156 ^ n18 ;
  assign n158 = n155 & ~n157 ;
  assign n159 = n158 ^ n18 ;
  assign n160 = ~n153 & n159 ;
  assign n161 = ~n152 & ~n160 ;
  assign n162 = ~n145 & n161 ;
  assign n163 = n162 ^ n128 ;
  assign n164 = n130 & n163 ;
  assign n165 = n164 ^ n128 ;
  assign n166 = n94 & n165 ;
  assign y0 = ~n166 ;
endmodule
