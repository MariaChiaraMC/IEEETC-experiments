module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 ;
  assign n36 = ~x1 & x5 ;
  assign n32 = ~x0 & x4 ;
  assign n33 = ~x2 & ~x3 ;
  assign n34 = n32 & n33 ;
  assign n7 = x4 ^ x2 ;
  assign n8 = x4 ^ x0 ;
  assign n9 = n8 ^ x2 ;
  assign n10 = ~n7 & ~n9 ;
  assign n11 = n10 ^ x2 ;
  assign n12 = n11 ^ x3 ;
  assign n13 = x5 ^ x4 ;
  assign n14 = ~x1 & n13 ;
  assign n15 = n14 ^ x1 ;
  assign n16 = n15 ^ x4 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = n17 ^ n9 ;
  assign n19 = n18 ^ x3 ;
  assign n20 = n13 ^ x3 ;
  assign n21 = n7 ^ x5 ;
  assign n22 = n21 ^ n9 ;
  assign n23 = n22 ^ x3 ;
  assign n24 = n20 & ~n23 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = n25 ^ x5 ;
  assign n27 = n19 & n26 ;
  assign n28 = n27 ^ x3 ;
  assign n29 = n12 & n28 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n30 ^ x3 ;
  assign n35 = n34 ^ n31 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = n37 ^ n31 ;
  assign n44 = n38 ^ n35 ;
  assign n45 = n44 ^ n31 ;
  assign n46 = n45 ^ n31 ;
  assign n47 = ~x1 & ~x2 ;
  assign n48 = ~x0 & ~n47 ;
  assign n49 = ~x4 & ~n48 ;
  assign n50 = n49 ^ n35 ;
  assign n51 = n50 ^ n35 ;
  assign n52 = n51 ^ n31 ;
  assign n53 = n46 & n52 ;
  assign n39 = x1 & ~x5 ;
  assign n40 = n39 ^ n35 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n41 ^ n31 ;
  assign n43 = n38 & n42 ;
  assign n54 = n53 ^ n43 ;
  assign n55 = n54 ^ n38 ;
  assign n56 = n43 ^ n31 ;
  assign n57 = n56 ^ n45 ;
  assign n58 = ~n31 & n57 ;
  assign n59 = n58 ^ n43 ;
  assign n60 = n55 & n59 ;
  assign n61 = n60 ^ n53 ;
  assign n62 = n61 ^ n58 ;
  assign n63 = n62 ^ n38 ;
  assign n64 = n63 ^ n31 ;
  assign n65 = n64 ^ n45 ;
  assign n66 = n65 ^ n34 ;
  assign y0 = n66 ;
endmodule
