module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 ;
  assign n8 = x1 & x6 ;
  assign n9 = x4 & x5 ;
  assign n10 = ~x2 & n9 ;
  assign n11 = x0 & x2 ;
  assign n12 = ~x4 & ~x5 ;
  assign n13 = n11 & n12 ;
  assign n14 = ~n10 & ~n13 ;
  assign n15 = n8 & ~n14 ;
  assign n16 = ~x6 & ~n12 ;
  assign n17 = ~x0 & n16 ;
  assign n18 = n17 ^ n12 ;
  assign n19 = x2 ^ x1 ;
  assign n20 = x3 & ~n19 ;
  assign n21 = n18 & n20 ;
  assign n22 = ~n15 & ~n21 ;
  assign n23 = x0 & n10 ;
  assign n24 = ~x6 & n23 ;
  assign n25 = ~n11 & n19 ;
  assign n26 = ~x4 & x6 ;
  assign n27 = x5 & n26 ;
  assign n28 = ~n25 & n27 ;
  assign n29 = ~n24 & ~n28 ;
  assign n30 = x6 ^ x5 ;
  assign n31 = n30 ^ x2 ;
  assign n32 = n31 ^ x1 ;
  assign n35 = x6 ^ x0 ;
  assign n36 = n35 ^ n31 ;
  assign n33 = x2 ^ x0 ;
  assign n34 = n33 ^ x0 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = n37 ^ x1 ;
  assign n39 = ~n32 & n38 ;
  assign n40 = n39 ^ x0 ;
  assign n41 = n40 ^ n31 ;
  assign n42 = n41 ^ x1 ;
  assign n43 = n31 ^ x0 ;
  assign n44 = n43 ^ n36 ;
  assign n45 = x1 & n44 ;
  assign n46 = n45 ^ x0 ;
  assign n47 = n46 ^ n31 ;
  assign n48 = n47 ^ n33 ;
  assign n49 = n48 ^ n36 ;
  assign n50 = x6 ^ x4 ;
  assign n51 = n50 ^ x6 ;
  assign n52 = n51 ^ x0 ;
  assign n53 = n52 ^ n31 ;
  assign n54 = n53 ^ n33 ;
  assign n55 = n54 ^ n36 ;
  assign n56 = ~n53 & ~n55 ;
  assign n57 = n56 ^ x0 ;
  assign n58 = n57 ^ n33 ;
  assign n59 = n58 ^ n36 ;
  assign n60 = ~n49 & n59 ;
  assign n61 = n60 ^ n31 ;
  assign n62 = n61 ^ n33 ;
  assign n63 = n62 ^ n36 ;
  assign n64 = n63 ^ x1 ;
  assign n65 = ~n42 & ~n64 ;
  assign n66 = n65 ^ n45 ;
  assign n67 = n66 ^ n60 ;
  assign n68 = n67 ^ n31 ;
  assign n69 = n68 ^ n33 ;
  assign n70 = n69 ^ n36 ;
  assign n71 = n29 & n70 ;
  assign n72 = ~x1 & x2 ;
  assign n73 = x4 & x6 ;
  assign n74 = n73 ^ x5 ;
  assign n75 = x5 ^ x0 ;
  assign n76 = ~n74 & n75 ;
  assign n77 = n76 ^ x5 ;
  assign n78 = n72 & ~n77 ;
  assign n79 = n71 & ~n78 ;
  assign n80 = n79 ^ x3 ;
  assign n81 = n80 ^ n79 ;
  assign n82 = ~x5 & n73 ;
  assign n83 = x0 & x1 ;
  assign n84 = n82 & n83 ;
  assign n85 = ~n12 & n72 ;
  assign n86 = ~n73 & n85 ;
  assign n87 = ~n84 & ~n86 ;
  assign n88 = n73 ^ x0 ;
  assign n89 = x5 ^ x1 ;
  assign n90 = n89 ^ x1 ;
  assign n91 = n90 ^ n88 ;
  assign n92 = n73 ^ n8 ;
  assign n93 = ~n73 & ~n92 ;
  assign n94 = n93 ^ x1 ;
  assign n95 = n94 ^ n73 ;
  assign n96 = n91 & n95 ;
  assign n97 = n96 ^ n93 ;
  assign n98 = n97 ^ n73 ;
  assign n99 = n88 & ~n98 ;
  assign n100 = n99 ^ n73 ;
  assign n101 = ~x2 & n100 ;
  assign n102 = n87 & ~n101 ;
  assign n103 = ~n13 & n102 ;
  assign n104 = n103 ^ n79 ;
  assign n105 = n81 & n104 ;
  assign n106 = n105 ^ n79 ;
  assign n107 = n22 & n106 ;
  assign y0 = ~n107 ;
endmodule
