module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 ;
  assign n9 = x7 ^ x1 ;
  assign n10 = n9 ^ x1 ;
  assign n11 = n10 ^ x5 ;
  assign n12 = x2 ^ x0 ;
  assign n13 = x0 & n12 ;
  assign n14 = n13 ^ x1 ;
  assign n15 = n14 ^ x0 ;
  assign n16 = n11 & n15 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n17 ^ x0 ;
  assign n19 = x5 & n18 ;
  assign n20 = n19 ^ x5 ;
  assign n21 = x6 & ~n20 ;
  assign n22 = ~x2 & x7 ;
  assign n23 = n22 ^ x1 ;
  assign n24 = n23 ^ x1 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = x6 ^ x0 ;
  assign n27 = ~x6 & n26 ;
  assign n28 = n27 ^ x1 ;
  assign n29 = n28 ^ x6 ;
  assign n30 = ~n25 & ~n29 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n31 ^ x6 ;
  assign n33 = x5 & ~n32 ;
  assign n34 = ~n21 & ~n33 ;
  assign n35 = ~x4 & ~n34 ;
  assign n36 = x5 & ~x6 ;
  assign n37 = ~x1 & ~n36 ;
  assign n38 = ~x2 & ~n37 ;
  assign n39 = x4 ^ x0 ;
  assign n40 = x5 ^ x1 ;
  assign n41 = n40 ^ x1 ;
  assign n42 = x2 & x7 ;
  assign n43 = ~x1 & n42 ;
  assign n44 = ~x6 & ~n43 ;
  assign n45 = n44 ^ x1 ;
  assign n46 = ~n41 & ~n45 ;
  assign n47 = n46 ^ x1 ;
  assign n48 = n47 ^ x4 ;
  assign n49 = n39 & ~n48 ;
  assign n50 = n49 ^ n46 ;
  assign n51 = n50 ^ x1 ;
  assign n52 = n51 ^ x0 ;
  assign n53 = x4 & ~n52 ;
  assign n54 = n53 ^ x4 ;
  assign n55 = ~n38 & n54 ;
  assign n56 = ~n35 & ~n55 ;
  assign n57 = ~x3 & ~n56 ;
  assign n58 = x2 & x6 ;
  assign n59 = x0 & ~x1 ;
  assign n60 = ~n58 & n59 ;
  assign n61 = x3 & ~x4 ;
  assign n62 = ~n42 & n61 ;
  assign n63 = n60 & n62 ;
  assign n64 = ~x5 & n63 ;
  assign n65 = ~n57 & ~n64 ;
  assign y0 = ~n65 ;
endmodule
