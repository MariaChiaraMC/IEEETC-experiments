module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 ;
  assign n15 = x6 & x7 ;
  assign n16 = ~x8 & n15 ;
  assign n17 = ~x10 & ~n16 ;
  assign n18 = x0 & x1 ;
  assign n19 = ~x11 & ~n18 ;
  assign n20 = ~x3 & ~x9 ;
  assign n21 = x2 & ~n20 ;
  assign n22 = ~n19 & n21 ;
  assign n23 = ~n17 & ~n22 ;
  assign n24 = x7 ^ x6 ;
  assign n25 = n24 ^ x8 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n24 ^ x7 ;
  assign n28 = n27 ^ n24 ;
  assign n29 = ~n26 & n28 ;
  assign n30 = n29 ^ n24 ;
  assign n31 = x5 & ~n30 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = ~x4 & ~n32 ;
  assign n34 = ~n23 & ~n33 ;
  assign n35 = x12 & ~n34 ;
  assign n36 = ~x4 & ~x10 ;
  assign n37 = x13 & ~n36 ;
  assign n38 = ~n17 & n37 ;
  assign n39 = x11 & n38 ;
  assign n40 = ~n35 & ~n39 ;
  assign y0 = ~n40 ;
endmodule
