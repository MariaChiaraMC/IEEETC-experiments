module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 ;
  output y0 ;
  wire n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 ;
  assign n28 = ~x0 & ~x3 ;
  assign n29 = ~x16 & n28 ;
  assign n30 = ~x2 & ~x23 ;
  assign n31 = ~x1 & n30 ;
  assign n32 = n29 & n31 ;
  assign n33 = x5 & n32 ;
  assign n34 = n33 ^ x13 ;
  assign n35 = n34 ^ n33 ;
  assign n36 = x0 & x3 ;
  assign n37 = x16 & n36 ;
  assign n38 = x2 & x23 ;
  assign n39 = x1 & n38 ;
  assign n40 = n37 & n39 ;
  assign n41 = n40 ^ n33 ;
  assign n42 = n41 ^ n33 ;
  assign n43 = n35 & n42 ;
  assign n44 = n43 ^ n33 ;
  assign n45 = x4 & n44 ;
  assign n46 = n45 ^ n33 ;
  assign n47 = x8 ^ x7 ;
  assign n48 = x8 & ~n47 ;
  assign n49 = x6 & n48 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = n46 & ~n50 ;
  assign n52 = ~x6 & ~x9 ;
  assign n53 = ~x4 & ~n52 ;
  assign n54 = n32 & n53 ;
  assign n55 = n40 ^ x4 ;
  assign n56 = x14 ^ x6 ;
  assign n57 = n56 ^ x14 ;
  assign n58 = x15 ^ x14 ;
  assign n59 = n57 & n58 ;
  assign n60 = n59 ^ x14 ;
  assign n61 = n60 ^ n40 ;
  assign n62 = n55 & n61 ;
  assign n63 = n62 ^ n59 ;
  assign n64 = n63 ^ x14 ;
  assign n65 = n64 ^ x4 ;
  assign n66 = n40 & n65 ;
  assign n67 = n66 ^ n40 ;
  assign n68 = ~n54 & ~n67 ;
  assign n69 = ~x7 & ~x8 ;
  assign n70 = ~x4 & ~x12 ;
  assign n71 = ~n69 & ~n70 ;
  assign n72 = n71 ^ x6 ;
  assign n73 = n72 ^ n71 ;
  assign n74 = ~x10 & ~x11 ;
  assign n75 = n74 ^ n71 ;
  assign n76 = ~n73 & n75 ;
  assign n77 = n76 ^ n71 ;
  assign n78 = ~n68 & n77 ;
  assign n79 = ~n51 & ~n78 ;
  assign y0 = ~n79 ;
endmodule
