module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 ;
  assign n9 = x0 & ~x3 ;
  assign n10 = ~x3 & ~x6 ;
  assign n11 = ~x7 & n10 ;
  assign n12 = ~n9 & ~n11 ;
  assign n13 = x5 ^ x1 ;
  assign n14 = n13 ^ n12 ;
  assign n16 = x2 & x7 ;
  assign n15 = x6 & x7 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = x5 & ~n17 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = ~n14 & n19 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n21 ^ n16 ;
  assign n23 = n22 ^ x5 ;
  assign n24 = n12 & n23 ;
  assign n25 = ~x4 & ~n24 ;
  assign n26 = x3 & x5 ;
  assign n27 = x7 & n26 ;
  assign n28 = ~x0 & x3 ;
  assign n29 = ~n27 & ~n28 ;
  assign n30 = ~n25 & n29 ;
  assign n31 = ~n10 & ~n26 ;
  assign n32 = x2 & ~n31 ;
  assign n33 = x6 ^ x4 ;
  assign n34 = n33 ^ x2 ;
  assign n35 = n34 ^ x6 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = ~x5 & ~x7 ;
  assign n38 = ~x3 & n37 ;
  assign n39 = n38 ^ n34 ;
  assign n40 = n39 ^ n33 ;
  assign n41 = n36 & ~n40 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = x0 & n38 ;
  assign n44 = n43 ^ n33 ;
  assign n45 = n42 & ~n44 ;
  assign n46 = n45 ^ n43 ;
  assign n47 = ~n33 & n46 ;
  assign n48 = n47 ^ n41 ;
  assign n49 = n48 ^ x4 ;
  assign n50 = n49 ^ n38 ;
  assign n51 = ~n32 & ~n50 ;
  assign n52 = ~x4 & ~n15 ;
  assign n53 = ~x1 & ~n52 ;
  assign n54 = n51 & ~n53 ;
  assign n55 = n30 & n54 ;
  assign y0 = n55 ;
endmodule
