module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 ;
  assign n10 = ~x7 & x8 ;
  assign n11 = x1 & ~x2 ;
  assign n12 = n10 & n11 ;
  assign n13 = x4 & n12 ;
  assign n14 = ~x1 & ~x4 ;
  assign n16 = x7 & x8 ;
  assign n15 = ~x7 & ~x8 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n16 ^ x2 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n17 & n19 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = n14 & n21 ;
  assign n23 = ~n13 & ~n22 ;
  assign n24 = ~x3 & x6 ;
  assign n25 = ~x5 & n24 ;
  assign n26 = ~n23 & n25 ;
  assign n73 = ~x1 & ~x2 ;
  assign n48 = x8 ^ x5 ;
  assign n74 = ~x3 & x4 ;
  assign n75 = n74 ^ x8 ;
  assign n76 = n75 ^ n74 ;
  assign n77 = x3 & ~x4 ;
  assign n78 = n77 ^ n74 ;
  assign n79 = ~n76 & n78 ;
  assign n80 = n79 ^ n74 ;
  assign n81 = ~n48 & n80 ;
  assign n82 = n73 & n81 ;
  assign n83 = ~x3 & x8 ;
  assign n84 = n14 ^ x4 ;
  assign n85 = n84 ^ n14 ;
  assign n60 = x1 & x2 ;
  assign n86 = n60 ^ n14 ;
  assign n87 = n86 ^ n14 ;
  assign n88 = ~n85 & n87 ;
  assign n89 = n88 ^ n14 ;
  assign n90 = x5 & n89 ;
  assign n91 = n90 ^ n14 ;
  assign n92 = n83 & n91 ;
  assign n27 = x3 & x8 ;
  assign n65 = x4 & ~x5 ;
  assign n93 = n60 & n65 ;
  assign n94 = n27 & n93 ;
  assign n95 = x5 & ~x8 ;
  assign n96 = ~x1 & x2 ;
  assign n97 = n95 & n96 ;
  assign n98 = x4 ^ x3 ;
  assign n99 = n97 & ~n98 ;
  assign n100 = ~n94 & ~n99 ;
  assign n101 = ~n92 & n100 ;
  assign n102 = ~n82 & n101 ;
  assign n41 = x1 & ~x3 ;
  assign n42 = ~n10 & n41 ;
  assign n28 = ~x4 & x5 ;
  assign n43 = ~x7 & ~n28 ;
  assign n44 = ~x5 & n43 ;
  assign n45 = n44 ^ n28 ;
  assign n46 = n42 & n45 ;
  assign n47 = x5 ^ x3 ;
  assign n49 = n47 & n48 ;
  assign n50 = n49 ^ x1 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = x5 & x8 ;
  assign n53 = n52 ^ n49 ;
  assign n54 = n51 & n53 ;
  assign n55 = n54 ^ n49 ;
  assign n56 = x4 & n55 ;
  assign n57 = ~x7 & n56 ;
  assign n58 = ~n46 & ~n57 ;
  assign n59 = ~x2 & ~n58 ;
  assign n61 = x3 & n60 ;
  assign n62 = ~x8 & n61 ;
  assign n63 = n28 ^ x7 ;
  assign n64 = n63 ^ n28 ;
  assign n66 = n65 ^ n28 ;
  assign n67 = n64 & n66 ;
  assign n68 = n67 ^ n28 ;
  assign n69 = n62 & n68 ;
  assign n70 = ~n59 & ~n69 ;
  assign n29 = n11 & n28 ;
  assign n30 = x5 ^ x4 ;
  assign n31 = x4 ^ x2 ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = ~x1 & n32 ;
  assign n34 = ~n29 & ~n33 ;
  assign n35 = n27 & ~n34 ;
  assign n36 = ~x2 & ~x4 ;
  assign n37 = ~x5 & ~x8 ;
  assign n38 = n36 & n37 ;
  assign n39 = ~x3 & n38 ;
  assign n40 = ~n35 & ~n39 ;
  assign n71 = n70 ^ n40 ;
  assign n72 = n71 ^ n40 ;
  assign n103 = n102 ^ n72 ;
  assign n104 = n103 ^ n71 ;
  assign n105 = n71 ^ x7 ;
  assign n106 = n105 ^ n71 ;
  assign n107 = n104 & n106 ;
  assign n108 = n107 ^ n71 ;
  assign n109 = x6 & n108 ;
  assign n110 = n109 ^ n70 ;
  assign n111 = n110 ^ x0 ;
  assign n112 = n111 ^ n110 ;
  assign n159 = n16 & n74 ;
  assign n116 = x6 & ~x8 ;
  assign n117 = n36 & n116 ;
  assign n118 = n117 ^ x3 ;
  assign n113 = n27 & n36 ;
  assign n114 = ~x6 & n113 ;
  assign n115 = n114 ^ x7 ;
  assign n119 = n118 ^ n115 ;
  assign n120 = n118 ^ n114 ;
  assign n121 = n120 ^ x3 ;
  assign n122 = ~n119 & ~n121 ;
  assign n123 = n122 ^ n114 ;
  assign n124 = x4 & ~x8 ;
  assign n125 = ~x6 & n124 ;
  assign n126 = ~x4 & x6 ;
  assign n127 = x8 & n126 ;
  assign n128 = ~n125 & ~n127 ;
  assign n129 = x2 & ~n128 ;
  assign n130 = ~n114 & ~n129 ;
  assign n131 = n130 ^ x3 ;
  assign n132 = ~n123 & ~n131 ;
  assign n133 = n132 ^ n130 ;
  assign n134 = ~x3 & n133 ;
  assign n135 = n134 ^ n122 ;
  assign n136 = n135 ^ x7 ;
  assign n137 = n136 ^ n114 ;
  assign n160 = n159 ^ n137 ;
  assign n138 = x8 ^ x4 ;
  assign n139 = x8 ^ x6 ;
  assign n147 = n139 ^ x8 ;
  assign n148 = n147 ^ x8 ;
  assign n149 = ~n147 & ~n148 ;
  assign n140 = n139 ^ x3 ;
  assign n141 = n140 ^ x7 ;
  assign n142 = n141 ^ n140 ;
  assign n143 = n140 ^ n139 ;
  assign n144 = n143 ^ x8 ;
  assign n145 = ~n142 & ~n144 ;
  assign n152 = n149 ^ n145 ;
  assign n146 = n145 ^ n138 ;
  assign n150 = n149 ^ n147 ;
  assign n151 = ~n146 & ~n150 ;
  assign n153 = n152 ^ n151 ;
  assign n154 = ~n138 & n153 ;
  assign n155 = n154 ^ n145 ;
  assign n156 = n155 ^ n149 ;
  assign n157 = n156 ^ n151 ;
  assign n158 = n157 ^ n137 ;
  assign n161 = n160 ^ n158 ;
  assign n162 = n158 ^ x2 ;
  assign n163 = n162 ^ n158 ;
  assign n164 = n161 & ~n163 ;
  assign n165 = n164 ^ n158 ;
  assign n166 = x1 & n165 ;
  assign n167 = n166 ^ n137 ;
  assign n168 = x5 & n167 ;
  assign n169 = x4 & x6 ;
  assign n170 = n27 & n73 ;
  assign n171 = n169 & n170 ;
  assign n172 = x7 & n171 ;
  assign n173 = x3 & ~x5 ;
  assign n174 = x7 ^ x6 ;
  assign n175 = n174 ^ x8 ;
  assign n176 = n10 & ~n175 ;
  assign n177 = n176 ^ n175 ;
  assign n178 = n96 & ~n177 ;
  assign n179 = ~x4 & n178 ;
  assign n180 = n127 ^ n125 ;
  assign n181 = n125 ^ x7 ;
  assign n182 = n181 ^ n125 ;
  assign n183 = n180 & n182 ;
  assign n184 = n183 ^ n125 ;
  assign n185 = n11 & n184 ;
  assign n186 = ~n179 & ~n185 ;
  assign n187 = n173 & ~n186 ;
  assign n188 = n65 & n83 ;
  assign n189 = ~x6 & x7 ;
  assign n190 = n96 & n189 ;
  assign n191 = n188 & n190 ;
  assign n192 = ~n187 & ~n191 ;
  assign n193 = ~n172 & n192 ;
  assign n194 = ~n168 & n193 ;
  assign n195 = n194 ^ n110 ;
  assign n196 = n112 & n195 ;
  assign n197 = n196 ^ n110 ;
  assign n198 = ~n26 & n197 ;
  assign y0 = ~n198 ;
endmodule
