module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ;
  assign n17 = x12 & ~x15 ;
  assign n18 = x10 & n17 ;
  assign n19 = ~x10 & ~x13 ;
  assign n20 = x9 & n19 ;
  assign n21 = ~x0 & ~x14 ;
  assign n22 = ~x7 & ~x8 ;
  assign n23 = ~x6 & n22 ;
  assign n24 = ~x2 & ~n23 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n24 ^ x1 ;
  assign n28 = n26 & n27 ;
  assign n29 = n28 ^ n24 ;
  assign n30 = n21 & n29 ;
  assign n31 = n30 ^ x11 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = x3 & x4 ;
  assign n34 = x0 & n33 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = ~n32 & n35 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = n20 & n37 ;
  assign n39 = ~n18 & ~n38 ;
  assign y0 = n39 ;
endmodule
