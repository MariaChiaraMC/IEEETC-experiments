module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n9 = x3 ^ x2 ;
  assign n10 = n9 ^ x3 ;
  assign n11 = n10 ^ x0 ;
  assign n12 = x5 ^ x4 ;
  assign n13 = n12 ^ x6 ;
  assign n14 = x6 ^ x5 ;
  assign n15 = n14 ^ x6 ;
  assign n16 = x7 ^ x6 ;
  assign n17 = n15 & ~n16 ;
  assign n18 = n17 ^ x6 ;
  assign n19 = n13 & n18 ;
  assign n20 = ~x1 & n19 ;
  assign n21 = n20 ^ x1 ;
  assign n22 = ~x3 & ~n21 ;
  assign n23 = n22 ^ x1 ;
  assign n24 = n11 & n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n25 ^ x1 ;
  assign n27 = n26 ^ x3 ;
  assign n28 = ~x0 & ~n27 ;
  assign y0 = n28 ;
endmodule
