module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 ;
  output y0 ;
  wire n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 ;
  assign n19 = ~x13 & x14 ;
  assign n20 = ~x3 & ~x13 ;
  assign n21 = x4 & x6 ;
  assign n22 = x7 & x8 ;
  assign n23 = n21 & ~n22 ;
  assign n24 = x15 ^ x5 ;
  assign n25 = n23 & ~n24 ;
  assign n26 = n20 & ~n25 ;
  assign n27 = ~x14 & ~n26 ;
  assign n28 = ~n19 & ~n27 ;
  assign n29 = x17 & ~n28 ;
  assign n30 = ~x5 & ~x15 ;
  assign n31 = x14 ^ x13 ;
  assign n32 = x14 ^ x6 ;
  assign n33 = n32 ^ x6 ;
  assign n34 = ~x2 & ~x9 ;
  assign n35 = n34 ^ x6 ;
  assign n36 = n33 & ~n35 ;
  assign n37 = n36 ^ x6 ;
  assign n38 = n31 & ~n37 ;
  assign n39 = ~x7 & ~x8 ;
  assign n40 = n39 ^ x7 ;
  assign n41 = x6 & n40 ;
  assign n42 = n41 ^ x7 ;
  assign n43 = n38 & n42 ;
  assign n44 = n30 & n43 ;
  assign n45 = ~n29 & ~n44 ;
  assign n46 = n45 ^ x17 ;
  assign n47 = n46 ^ x16 ;
  assign n56 = n47 ^ n46 ;
  assign n48 = x5 & x15 ;
  assign n49 = n43 & n48 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = n50 ^ n46 ;
  assign n52 = n47 ^ n45 ;
  assign n53 = n52 ^ n49 ;
  assign n54 = n53 ^ n51 ;
  assign n55 = ~n51 & n54 ;
  assign n57 = n56 ^ n55 ;
  assign n58 = n57 ^ n51 ;
  assign n59 = x5 & n39 ;
  assign n60 = ~x6 & n59 ;
  assign n61 = x4 & n60 ;
  assign n62 = ~x5 & x7 ;
  assign n63 = x6 & n62 ;
  assign n64 = n63 ^ x3 ;
  assign n65 = n64 ^ n63 ;
  assign n66 = n21 & n62 ;
  assign n67 = n66 ^ n63 ;
  assign n68 = n67 ^ n63 ;
  assign n69 = ~n65 & ~n68 ;
  assign n70 = n69 ^ n63 ;
  assign n71 = ~x13 & n70 ;
  assign n72 = n71 ^ n63 ;
  assign n73 = ~n61 & n72 ;
  assign n74 = ~x14 & ~n73 ;
  assign n75 = n19 & n34 ;
  assign n76 = n63 ^ n34 ;
  assign n77 = n75 ^ n59 ;
  assign n78 = ~n76 & n77 ;
  assign n79 = n78 ^ n59 ;
  assign n80 = n75 & n79 ;
  assign n81 = n80 ^ n19 ;
  assign n82 = ~n74 & ~n81 ;
  assign n83 = x15 & ~n82 ;
  assign n84 = x1 & ~x15 ;
  assign n85 = ~x13 & ~x14 ;
  assign n86 = n85 ^ n84 ;
  assign n87 = ~x10 & x11 ;
  assign n88 = n87 ^ x12 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = n87 ^ x10 ;
  assign n91 = ~n89 & n90 ;
  assign n92 = n91 ^ n87 ;
  assign n93 = n92 ^ n84 ;
  assign n94 = n86 & n93 ;
  assign n95 = n94 ^ n91 ;
  assign n96 = n95 ^ n87 ;
  assign n97 = n96 ^ n85 ;
  assign n98 = n84 & n97 ;
  assign n99 = n98 ^ n84 ;
  assign n100 = ~n83 & ~n99 ;
  assign n101 = n100 ^ n46 ;
  assign n102 = n55 ^ n51 ;
  assign n103 = n101 & ~n102 ;
  assign n104 = n103 ^ n46 ;
  assign n105 = ~n58 & n104 ;
  assign n106 = n105 ^ n46 ;
  assign n107 = n106 ^ x17 ;
  assign n108 = n107 ^ n46 ;
  assign n109 = ~x0 & ~n108 ;
  assign y0 = n109 ;
endmodule
