module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n11 = ~x5 & ~x7 ;
  assign n12 = ~x4 & x9 ;
  assign n13 = ~x1 & n12 ;
  assign n14 = n11 & n13 ;
  assign n15 = x2 ^ x0 ;
  assign n16 = n15 ^ x3 ;
  assign n17 = n16 ^ x6 ;
  assign n18 = x6 ^ x3 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = x8 ^ x2 ;
  assign n21 = ~x2 & n20 ;
  assign n22 = n21 ^ x3 ;
  assign n23 = n22 ^ x2 ;
  assign n24 = n19 & n23 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ x2 ;
  assign n27 = n17 & ~n26 ;
  assign n28 = n14 & n27 ;
  assign y0 = n28 ;
endmodule
