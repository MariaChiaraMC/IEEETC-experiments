module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n23 = ~x1 & ~x2 ;
  assign n10 = x8 ^ x7 ;
  assign n11 = ~x2 & n10 ;
  assign n12 = n11 ^ x7 ;
  assign n14 = n12 ^ x5 ;
  assign n13 = n12 ^ x6 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = n14 ^ x2 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = n15 & ~n17 ;
  assign n19 = n18 ^ n14 ;
  assign n20 = x1 & n19 ;
  assign n21 = n20 ^ n12 ;
  assign n22 = n21 ^ x3 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n21 ^ x4 ;
  assign n27 = n26 ^ n22 ;
  assign n28 = n25 & n27 ;
  assign n29 = n28 ^ n22 ;
  assign n30 = x0 & n29 ;
  assign n31 = n30 ^ n21 ;
  assign y0 = n31 ;
endmodule
