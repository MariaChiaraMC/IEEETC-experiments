module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 ;
  assign n15 = x4 ^ x3 ;
  assign n22 = n15 ^ x5 ;
  assign n16 = n15 ^ x1 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = x4 ^ x1 ;
  assign n19 = n18 ^ x1 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = ~n17 & n20 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n23 ^ n17 ;
  assign n25 = x6 ^ x5 ;
  assign n26 = n25 ^ x5 ;
  assign n27 = n21 ^ n17 ;
  assign n28 = n26 & ~n27 ;
  assign n29 = n28 ^ x5 ;
  assign n30 = n24 & ~n29 ;
  assign n31 = n30 ^ x5 ;
  assign n32 = n31 ^ x5 ;
  assign n33 = ~x2 & n32 ;
  assign n34 = ~x10 & ~x11 ;
  assign n35 = x5 & ~x13 ;
  assign n36 = n34 & n35 ;
  assign n37 = x2 & n36 ;
  assign n38 = x9 ^ x8 ;
  assign n39 = x8 ^ x7 ;
  assign n40 = n38 & ~n39 ;
  assign n41 = n40 ^ x8 ;
  assign n42 = ~x12 & ~n41 ;
  assign n43 = n37 & n42 ;
  assign n44 = x1 & x6 ;
  assign n45 = ~n43 & n44 ;
  assign n46 = x5 & ~x6 ;
  assign n47 = ~x4 & ~n46 ;
  assign n48 = ~x1 & x2 ;
  assign n49 = ~x4 & ~n48 ;
  assign n50 = ~n47 & ~n49 ;
  assign n51 = ~n45 & n50 ;
  assign n52 = x3 & n51 ;
  assign n53 = ~n33 & ~n52 ;
  assign n54 = ~x0 & ~n53 ;
  assign y0 = n54 ;
endmodule
