// Benchmark "./pla/adr4.pla_res_4NonExact" written by ABC on Fri Nov 20 10:16:57 2020

module \./pla/adr4.pla_res_4NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = x0;
endmodule


