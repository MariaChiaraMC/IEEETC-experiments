module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 ;
  assign n9 = x5 ^ x1 ;
  assign n10 = x6 & ~x7 ;
  assign n11 = x2 & ~x3 ;
  assign n12 = n10 & n11 ;
  assign n13 = ~x0 & n12 ;
  assign n14 = n13 ^ x4 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = x0 & ~x2 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n15 & n17 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = n19 ^ x5 ;
  assign n21 = n9 & ~n20 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = n22 ^ n13 ;
  assign n24 = n23 ^ x1 ;
  assign n25 = ~x5 & ~n24 ;
  assign n26 = n25 ^ x5 ;
  assign y0 = n26 ;
endmodule
