module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 ;
  output y0 ;
  wire n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 ;
  assign n28 = x24 & x25 ;
  assign n29 = ~x7 & ~x8 ;
  assign n30 = n29 ^ x6 ;
  assign n31 = x12 ^ x0 ;
  assign n32 = n31 ^ x12 ;
  assign n33 = x15 ^ x12 ;
  assign n34 = n32 & n33 ;
  assign n35 = n34 ^ x12 ;
  assign n36 = n35 ^ n29 ;
  assign n37 = ~n30 & ~n36 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = n38 ^ x12 ;
  assign n40 = n39 ^ x6 ;
  assign n41 = ~n29 & n40 ;
  assign n42 = n41 ^ n29 ;
  assign n44 = x13 ^ x5 ;
  assign n45 = x5 ^ x0 ;
  assign n46 = n45 ^ x5 ;
  assign n47 = n44 & n46 ;
  assign n43 = x6 & x8 ;
  assign n48 = n47 ^ n43 ;
  assign n49 = n48 ^ x5 ;
  assign n50 = x8 ^ x7 ;
  assign n51 = n47 ^ x5 ;
  assign n52 = n50 & n51 ;
  assign n53 = n52 ^ n47 ;
  assign n54 = n53 ^ x5 ;
  assign n55 = n49 & n54 ;
  assign n56 = n42 & ~n55 ;
  assign n57 = ~x6 & ~x10 ;
  assign n58 = n57 ^ x11 ;
  assign n59 = x14 ^ x0 ;
  assign n60 = n59 ^ x14 ;
  assign n61 = x14 ^ x9 ;
  assign n62 = ~n60 & n61 ;
  assign n63 = n62 ^ x14 ;
  assign n64 = n63 ^ n57 ;
  assign n65 = ~n58 & n64 ;
  assign n66 = n65 ^ n62 ;
  assign n67 = n66 ^ x14 ;
  assign n68 = n67 ^ x11 ;
  assign n69 = n57 & ~n68 ;
  assign n70 = n69 ^ n57 ;
  assign n71 = n56 & ~n70 ;
  assign n72 = ~n28 & ~n71 ;
  assign y0 = n72 ;
endmodule
