module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n17 = x13 ^ x10 ;
  assign n18 = n17 ^ x12 ;
  assign n25 = n18 ^ n17 ;
  assign n21 = n17 ^ x14 ;
  assign n22 = n21 ^ n18 ;
  assign n19 = n18 ^ x13 ;
  assign n20 = n19 ^ x15 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n23 ^ n17 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n22 ^ n18 ;
  assign n28 = n27 ^ n17 ;
  assign n29 = n28 ^ n17 ;
  assign n30 = ~n23 & n29 ;
  assign n31 = n30 ^ n23 ;
  assign n32 = n28 & ~n31 ;
  assign n33 = n32 ^ n17 ;
  assign n34 = ~n26 & n33 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n35 ^ n17 ;
  assign n37 = n36 ^ x12 ;
  assign n38 = n37 ^ n25 ;
  assign y0 = n38 ;
endmodule
