module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 ;
  output y0 ;
  wire n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 ;
  assign n32 = ~x7 & ~x8 ;
  assign n33 = ~x23 & ~x24 ;
  assign n34 = ~x29 & ~x30 ;
  assign n35 = ~x28 & ~n34 ;
  assign n36 = ~x27 & ~n35 ;
  assign n37 = ~x25 & ~x26 ;
  assign n38 = ~n36 & n37 ;
  assign n39 = n33 & ~n38 ;
  assign n40 = ~x21 & ~x22 ;
  assign n41 = ~n39 & n40 ;
  assign n42 = ~x20 & ~n41 ;
  assign n43 = ~x19 & ~n42 ;
  assign n44 = ~x17 & ~x18 ;
  assign n45 = ~n43 & n44 ;
  assign n46 = ~x16 & ~n45 ;
  assign n47 = ~x15 & ~n46 ;
  assign n48 = ~x13 & ~x14 ;
  assign n49 = ~n47 & n48 ;
  assign n50 = ~x12 & ~n49 ;
  assign n51 = ~x11 & ~n50 ;
  assign n52 = ~x9 & ~x10 ;
  assign n53 = ~n51 & n52 ;
  assign n54 = n32 & ~n53 ;
  assign n55 = ~x5 & ~x6 ;
  assign n56 = ~n54 & n55 ;
  assign n57 = ~x4 & ~n56 ;
  assign n58 = ~x3 & ~n57 ;
  assign n59 = ~x1 & ~x2 ;
  assign n60 = ~n58 & n59 ;
  assign n61 = ~x0 & ~n60 ;
  assign y0 = n61 ;
endmodule
