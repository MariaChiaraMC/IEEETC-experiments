module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n17 = ~x8 & ~x15 ;
  assign n18 = x14 & ~n17 ;
  assign n19 = ~x11 & ~n18 ;
  assign n20 = ~x14 & n17 ;
  assign n21 = n20 ^ x13 ;
  assign n22 = x10 ^ x9 ;
  assign n23 = n22 ^ x8 ;
  assign n24 = n23 ^ x12 ;
  assign n25 = x15 ^ x9 ;
  assign n26 = ~x8 & n25 ;
  assign n27 = n26 ^ x15 ;
  assign n28 = n24 & ~n27 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = n29 ^ x15 ;
  assign n31 = n30 ^ x8 ;
  assign n32 = ~x12 & n31 ;
  assign n33 = ~n21 & n32 ;
  assign n34 = n19 & n33 ;
  assign n35 = ~x7 & ~n34 ;
  assign n36 = ~x5 & ~n35 ;
  assign n37 = ~x0 & ~n36 ;
  assign y0 = ~n37 ;
endmodule
