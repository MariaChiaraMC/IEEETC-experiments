module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 ;
  assign n11 = x3 & ~x5 ;
  assign n12 = x2 ^ x1 ;
  assign n13 = ~x6 & ~x8 ;
  assign n14 = ~x5 & ~n13 ;
  assign n15 = n14 ^ x2 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n16 ^ n12 ;
  assign n18 = x5 & x9 ;
  assign n19 = x5 & ~x6 ;
  assign n20 = ~n18 & ~n19 ;
  assign n21 = n20 ^ x8 ;
  assign n22 = ~n20 & n21 ;
  assign n23 = n22 ^ n14 ;
  assign n24 = n23 ^ n20 ;
  assign n25 = ~n17 & ~n24 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = n26 ^ n20 ;
  assign n28 = n12 & ~n27 ;
  assign n29 = n28 ^ x3 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = n30 ^ n11 ;
  assign n32 = x6 & x9 ;
  assign n33 = x2 & n13 ;
  assign n34 = x1 & n33 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = ~n32 & n35 ;
  assign n37 = n36 ^ n28 ;
  assign n38 = n37 ^ n32 ;
  assign n39 = ~n31 & n38 ;
  assign n40 = n39 ^ n36 ;
  assign n41 = n40 ^ n32 ;
  assign n42 = ~n11 & ~n41 ;
  assign n43 = n42 ^ n11 ;
  assign n44 = ~x0 & n43 ;
  assign n45 = ~x2 & ~x3 ;
  assign n46 = x1 & x8 ;
  assign n47 = ~x5 & ~x6 ;
  assign n48 = n46 & n47 ;
  assign n49 = n45 & n48 ;
  assign n50 = ~x1 & x3 ;
  assign n51 = ~x5 & ~x8 ;
  assign n52 = ~x2 & n51 ;
  assign n53 = ~n18 & ~n52 ;
  assign n54 = n50 & ~n53 ;
  assign n55 = x6 & n54 ;
  assign n56 = x0 & ~n55 ;
  assign n62 = x2 & ~x3 ;
  assign n57 = ~x1 & x8 ;
  assign n58 = n32 ^ x6 ;
  assign n59 = ~x5 & ~n58 ;
  assign n60 = n59 ^ x6 ;
  assign n61 = n57 & ~n60 ;
  assign n63 = n62 ^ n61 ;
  assign n64 = n63 ^ n61 ;
  assign n65 = n64 ^ n56 ;
  assign n66 = n32 & n51 ;
  assign n67 = ~n18 & ~n66 ;
  assign n68 = x2 & ~x8 ;
  assign n69 = ~x6 & ~n68 ;
  assign n70 = ~n11 & ~n69 ;
  assign n71 = x1 & n70 ;
  assign n72 = n71 ^ n67 ;
  assign n73 = ~n67 & ~n72 ;
  assign n74 = n73 ^ n61 ;
  assign n75 = n74 ^ n67 ;
  assign n76 = ~n65 & ~n75 ;
  assign n77 = n76 ^ n73 ;
  assign n78 = n77 ^ n67 ;
  assign n79 = n56 & ~n78 ;
  assign n80 = n79 ^ n56 ;
  assign n81 = ~n49 & n80 ;
  assign n82 = ~n44 & ~n81 ;
  assign n83 = ~x3 & x5 ;
  assign n84 = ~n11 & ~n83 ;
  assign n85 = n32 & ~n50 ;
  assign n86 = ~n84 & n85 ;
  assign n87 = x2 & n86 ;
  assign n88 = ~n82 & ~n87 ;
  assign n89 = ~x4 & ~n88 ;
  assign n90 = x6 ^ x4 ;
  assign n91 = ~x1 & ~x2 ;
  assign n92 = x4 & n91 ;
  assign n93 = ~x0 & ~x3 ;
  assign n94 = n92 & n93 ;
  assign n95 = ~n51 & n94 ;
  assign n96 = n95 ^ n90 ;
  assign n97 = n96 ^ x6 ;
  assign n98 = n97 ^ n96 ;
  assign n99 = x1 & ~x2 ;
  assign n100 = x3 & n99 ;
  assign n101 = x0 & ~x2 ;
  assign n102 = n50 & n101 ;
  assign n105 = x1 & ~x3 ;
  assign n103 = x8 & n50 ;
  assign n104 = x2 & ~n103 ;
  assign n106 = n105 ^ n104 ;
  assign n107 = ~x2 & ~x8 ;
  assign n108 = n107 ^ n104 ;
  assign n109 = n108 ^ n107 ;
  assign n110 = n107 ^ x0 ;
  assign n111 = n109 & ~n110 ;
  assign n112 = n111 ^ n107 ;
  assign n113 = n106 & ~n112 ;
  assign n114 = n113 ^ n105 ;
  assign n115 = ~n102 & ~n114 ;
  assign n116 = n115 ^ x6 ;
  assign n117 = n116 ^ n115 ;
  assign n118 = ~n50 & ~n105 ;
  assign n119 = ~n68 & ~n118 ;
  assign n120 = ~n101 & n119 ;
  assign n121 = ~x0 & x2 ;
  assign n122 = ~x1 & ~n121 ;
  assign n123 = n101 ^ x3 ;
  assign n124 = x8 & ~n123 ;
  assign n125 = n124 ^ x3 ;
  assign n126 = n122 & ~n125 ;
  assign n127 = ~n120 & ~n126 ;
  assign n128 = n127 ^ n115 ;
  assign n129 = n117 & n128 ;
  assign n130 = n129 ^ n115 ;
  assign n131 = ~n100 & n130 ;
  assign n132 = n131 ^ x3 ;
  assign n133 = n132 ^ n131 ;
  assign n134 = ~x0 & ~x8 ;
  assign n135 = n91 & n134 ;
  assign n136 = n135 ^ n131 ;
  assign n137 = n136 ^ n131 ;
  assign n138 = ~n133 & n137 ;
  assign n139 = n138 ^ n131 ;
  assign n140 = x5 & ~n139 ;
  assign n141 = n140 ^ n131 ;
  assign n142 = n141 ^ n96 ;
  assign n143 = n142 ^ n90 ;
  assign n144 = ~n98 & n143 ;
  assign n145 = n144 ^ n141 ;
  assign n146 = x3 ^ x2 ;
  assign n147 = n51 ^ x2 ;
  assign n148 = n147 ^ x2 ;
  assign n149 = n146 & ~n148 ;
  assign n150 = n149 ^ x2 ;
  assign n151 = ~x1 & n150 ;
  assign n152 = ~x0 & n151 ;
  assign n153 = x3 & ~x8 ;
  assign n154 = n101 & ~n153 ;
  assign n155 = n118 ^ x0 ;
  assign n156 = n155 ^ n118 ;
  assign n157 = ~n62 & ~n100 ;
  assign n158 = ~n46 & n157 ;
  assign n159 = n158 ^ n118 ;
  assign n160 = ~n156 & n159 ;
  assign n161 = n160 ^ n118 ;
  assign n162 = ~n154 & n161 ;
  assign n163 = n162 ^ x3 ;
  assign n164 = n163 ^ n162 ;
  assign n165 = n162 ^ n121 ;
  assign n166 = n165 ^ n162 ;
  assign n167 = n164 & n166 ;
  assign n168 = n167 ^ n162 ;
  assign n169 = ~x5 & ~n168 ;
  assign n170 = n169 ^ n162 ;
  assign n171 = ~n152 & n170 ;
  assign n172 = n141 & n171 ;
  assign n173 = n172 ^ n90 ;
  assign n174 = n145 & ~n173 ;
  assign n175 = n174 ^ n172 ;
  assign n176 = ~n90 & n175 ;
  assign n177 = n176 ^ n144 ;
  assign n178 = n177 ^ x4 ;
  assign n179 = n178 ^ n141 ;
  assign n180 = n179 ^ x9 ;
  assign n181 = n180 ^ n179 ;
  assign n182 = n181 ^ n89 ;
  assign n183 = n94 ^ x6 ;
  assign n184 = x6 & n183 ;
  assign n185 = n184 ^ n179 ;
  assign n186 = n185 ^ x6 ;
  assign n187 = ~n182 & ~n186 ;
  assign n188 = n187 ^ n184 ;
  assign n189 = n188 ^ x6 ;
  assign n190 = ~n89 & n189 ;
  assign n191 = n190 ^ n89 ;
  assign n192 = ~x7 & n191 ;
  assign n193 = ~x9 & ~n122 ;
  assign n194 = x8 & ~n193 ;
  assign n195 = ~x3 & x7 ;
  assign n196 = n47 & n195 ;
  assign n197 = ~x4 & n196 ;
  assign n198 = ~n194 & n197 ;
  assign n199 = n121 ^ x1 ;
  assign n200 = n199 ^ n12 ;
  assign n201 = n200 ^ n134 ;
  assign n202 = n201 ^ n200 ;
  assign n203 = n200 ^ n199 ;
  assign n204 = n203 ^ x1 ;
  assign n205 = ~n202 & ~n204 ;
  assign n206 = n205 ^ n199 ;
  assign n207 = ~x9 & ~n199 ;
  assign n208 = n207 ^ x1 ;
  assign n209 = ~n206 & ~n208 ;
  assign n210 = n209 ^ n207 ;
  assign n211 = ~x1 & n210 ;
  assign n212 = n211 ^ n205 ;
  assign n213 = n212 ^ n121 ;
  assign n214 = n213 ^ n199 ;
  assign n215 = n198 & ~n214 ;
  assign n216 = ~n192 & ~n215 ;
  assign y0 = ~n216 ;
endmodule
