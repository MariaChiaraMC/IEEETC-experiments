module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 ;
  assign n11 = ~x0 & ~x1 ;
  assign n12 = ~x2 & x4 ;
  assign n13 = ~x8 & n12 ;
  assign n14 = n11 & n13 ;
  assign n15 = x5 ^ x3 ;
  assign n16 = x9 ^ x5 ;
  assign n17 = ~n15 & ~n16 ;
  assign n18 = n14 & n17 ;
  assign n19 = ~x4 & x8 ;
  assign n20 = x2 ^ x1 ;
  assign n21 = ~x5 & ~x9 ;
  assign n22 = ~x3 & n21 ;
  assign n23 = n22 ^ x2 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ n20 ;
  assign n26 = x5 & x9 ;
  assign n27 = ~x0 & x3 ;
  assign n28 = x0 & ~x3 ;
  assign n29 = ~n27 & ~n28 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n26 & ~n30 ;
  assign n32 = n31 ^ n22 ;
  assign n33 = n32 ^ n26 ;
  assign n34 = ~n25 & n33 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = n35 ^ n26 ;
  assign n37 = ~n20 & n36 ;
  assign n38 = n19 & n37 ;
  assign n39 = ~n18 & ~n38 ;
  assign n40 = ~x7 & ~n39 ;
  assign n41 = x0 & ~x5 ;
  assign n42 = x3 & n41 ;
  assign n43 = x8 & x9 ;
  assign n44 = n12 & n43 ;
  assign n45 = n44 ^ x2 ;
  assign n46 = n45 ^ n44 ;
  assign n47 = ~x8 & ~x9 ;
  assign n48 = ~x4 & n47 ;
  assign n49 = n48 ^ n44 ;
  assign n50 = n49 ^ n44 ;
  assign n51 = n46 & n50 ;
  assign n52 = n51 ^ n44 ;
  assign n53 = ~x1 & n52 ;
  assign n54 = n53 ^ n44 ;
  assign n55 = n42 & n54 ;
  assign n56 = ~x0 & n48 ;
  assign n57 = ~x2 & x5 ;
  assign n58 = x1 & n57 ;
  assign n59 = ~x1 & x2 ;
  assign n60 = ~x5 & n59 ;
  assign n61 = ~n58 & ~n60 ;
  assign n62 = n56 & ~n61 ;
  assign n63 = x4 & x8 ;
  assign n64 = ~x1 & ~x2 ;
  assign n65 = x0 & n64 ;
  assign n66 = n26 & n65 ;
  assign n67 = n63 & n66 ;
  assign n68 = ~n62 & ~n67 ;
  assign n69 = ~x3 & ~n68 ;
  assign n70 = x0 & x5 ;
  assign n71 = ~x3 & x8 ;
  assign n72 = x4 & ~x9 ;
  assign n73 = n71 & n72 ;
  assign n74 = ~x2 & ~x9 ;
  assign n75 = n71 & n74 ;
  assign n76 = ~x2 & x3 ;
  assign n77 = ~x4 & x9 ;
  assign n78 = n76 & n77 ;
  assign n79 = ~n75 & ~n78 ;
  assign n80 = ~n73 & n79 ;
  assign n81 = n70 & ~n80 ;
  assign n82 = ~x1 & ~n81 ;
  assign n83 = x3 & x9 ;
  assign n84 = ~x4 & ~x5 ;
  assign n85 = x2 & n84 ;
  assign n88 = n85 ^ x4 ;
  assign n86 = x4 & ~x5 ;
  assign n87 = n86 ^ n85 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = n88 ^ x2 ;
  assign n91 = n90 ^ n88 ;
  assign n92 = ~n89 & n91 ;
  assign n93 = n92 ^ n88 ;
  assign n94 = x0 & ~n93 ;
  assign n95 = n94 ^ n85 ;
  assign n96 = n83 & n95 ;
  assign n97 = x4 & n57 ;
  assign n98 = n27 & n97 ;
  assign n99 = ~x0 & x4 ;
  assign n100 = x0 & ~n12 ;
  assign n101 = n22 & ~n100 ;
  assign n102 = ~n99 & n101 ;
  assign n103 = ~n98 & ~n102 ;
  assign n104 = ~n96 & n103 ;
  assign n105 = ~x8 & ~n104 ;
  assign n106 = x9 & n71 ;
  assign n107 = n106 ^ n41 ;
  assign n108 = ~n85 & ~n97 ;
  assign n109 = n108 ^ n107 ;
  assign n110 = n109 ^ n106 ;
  assign n111 = n110 ^ n109 ;
  assign n112 = x2 & ~x3 ;
  assign n113 = n77 & n112 ;
  assign n114 = x2 & x8 ;
  assign n115 = n72 & n114 ;
  assign n116 = ~n113 & ~n115 ;
  assign n117 = n116 ^ n109 ;
  assign n118 = n117 ^ n107 ;
  assign n119 = n111 & ~n118 ;
  assign n120 = n119 ^ n116 ;
  assign n121 = ~x4 & n116 ;
  assign n122 = n121 ^ n107 ;
  assign n123 = n120 & ~n122 ;
  assign n124 = n123 ^ n121 ;
  assign n125 = ~n107 & n124 ;
  assign n126 = n125 ^ n119 ;
  assign n127 = n126 ^ n41 ;
  assign n128 = n127 ^ n116 ;
  assign n129 = ~n105 & ~n128 ;
  assign n130 = n82 & n129 ;
  assign n131 = ~x0 & x5 ;
  assign n132 = x3 & x8 ;
  assign n133 = n74 & n132 ;
  assign n134 = n131 & n133 ;
  assign n135 = x1 & ~n134 ;
  assign n136 = n131 ^ x0 ;
  assign n137 = n136 ^ x8 ;
  assign n138 = n137 ^ x9 ;
  assign n146 = n138 ^ n136 ;
  assign n139 = ~x5 & x8 ;
  assign n140 = n139 ^ n138 ;
  assign n141 = n140 ^ n136 ;
  assign n142 = n138 ^ n131 ;
  assign n143 = n142 ^ n139 ;
  assign n144 = n143 ^ n141 ;
  assign n145 = ~n141 & ~n144 ;
  assign n147 = n146 ^ n145 ;
  assign n148 = n147 ^ n141 ;
  assign n149 = n136 ^ x9 ;
  assign n150 = n145 ^ n141 ;
  assign n151 = n149 & ~n150 ;
  assign n152 = n151 ^ n136 ;
  assign n153 = ~n148 & n152 ;
  assign n154 = n153 ^ n136 ;
  assign n155 = n154 ^ x0 ;
  assign n156 = n155 ^ n136 ;
  assign n157 = n112 & n156 ;
  assign n158 = x8 ^ x5 ;
  assign n159 = x9 ^ x0 ;
  assign n160 = x8 ^ x0 ;
  assign n161 = n160 ^ x0 ;
  assign n162 = n159 & n161 ;
  assign n163 = n162 ^ x0 ;
  assign n164 = n158 & ~n163 ;
  assign n165 = n76 & n164 ;
  assign n166 = ~n157 & ~n165 ;
  assign n167 = n166 ^ x4 ;
  assign n168 = n167 ^ n166 ;
  assign n169 = n168 ^ n135 ;
  assign n170 = ~x3 & ~x8 ;
  assign n171 = ~x0 & x2 ;
  assign n172 = n170 & n171 ;
  assign n173 = ~x9 & ~n172 ;
  assign n174 = x3 & n114 ;
  assign n177 = n174 ^ n132 ;
  assign n178 = n177 ^ n174 ;
  assign n175 = n174 ^ x0 ;
  assign n176 = n175 ^ n174 ;
  assign n179 = n178 ^ n176 ;
  assign n180 = n174 ^ x2 ;
  assign n181 = n180 ^ n174 ;
  assign n182 = n181 ^ n178 ;
  assign n183 = ~n178 & n182 ;
  assign n184 = n183 ^ n178 ;
  assign n185 = ~n179 & ~n184 ;
  assign n186 = n185 ^ n183 ;
  assign n187 = n186 ^ n174 ;
  assign n188 = n187 ^ n178 ;
  assign n189 = x5 & ~n188 ;
  assign n190 = n189 ^ n174 ;
  assign n191 = n173 & ~n190 ;
  assign n192 = n70 & n174 ;
  assign n193 = ~x0 & ~x5 ;
  assign n194 = x8 ^ x3 ;
  assign n195 = x3 ^ x2 ;
  assign n196 = n194 & n195 ;
  assign n197 = n193 & n196 ;
  assign n198 = x9 & ~n197 ;
  assign n199 = ~n192 & n198 ;
  assign n200 = n199 ^ n191 ;
  assign n201 = ~n191 & n200 ;
  assign n202 = n201 ^ n166 ;
  assign n203 = n202 ^ n191 ;
  assign n204 = n169 & n203 ;
  assign n205 = n204 ^ n201 ;
  assign n206 = n205 ^ n191 ;
  assign n207 = n135 & ~n206 ;
  assign n208 = n207 ^ n135 ;
  assign n209 = ~n130 & ~n208 ;
  assign n210 = n42 & n48 ;
  assign n211 = x2 & n210 ;
  assign n212 = ~n209 & ~n211 ;
  assign n213 = n212 ^ x7 ;
  assign n214 = n213 ^ n212 ;
  assign n215 = x9 ^ x4 ;
  assign n217 = n215 ^ x0 ;
  assign n216 = n215 ^ x1 ;
  assign n218 = n217 ^ n216 ;
  assign n219 = n218 ^ x9 ;
  assign n224 = n219 ^ n215 ;
  assign n225 = n224 ^ n217 ;
  assign n226 = n225 ^ n217 ;
  assign n227 = n215 ^ x9 ;
  assign n228 = n227 ^ n215 ;
  assign n229 = n228 ^ n217 ;
  assign n230 = n226 & n229 ;
  assign n220 = n215 ^ x5 ;
  assign n221 = n220 ^ n219 ;
  assign n222 = n221 ^ n217 ;
  assign n223 = n219 & n222 ;
  assign n231 = n230 ^ n223 ;
  assign n232 = n231 ^ n219 ;
  assign n233 = n223 ^ n217 ;
  assign n234 = n233 ^ n225 ;
  assign n235 = n217 & n234 ;
  assign n236 = n235 ^ n223 ;
  assign n237 = n232 & n236 ;
  assign n238 = n237 ^ n230 ;
  assign n239 = n238 ^ n235 ;
  assign n240 = n239 ^ n219 ;
  assign n241 = n240 ^ n217 ;
  assign n242 = n241 ^ n225 ;
  assign n243 = n76 & n242 ;
  assign n244 = ~n21 & ~n58 ;
  assign n245 = x4 & n28 ;
  assign n246 = ~n74 & n245 ;
  assign n247 = ~n244 & n246 ;
  assign n248 = x0 & x3 ;
  assign n249 = x9 & n86 ;
  assign n250 = ~n248 & n249 ;
  assign n251 = n64 & n250 ;
  assign n252 = ~n247 & ~n251 ;
  assign n253 = x1 & ~x4 ;
  assign n254 = ~x1 & x4 ;
  assign n255 = ~n253 & ~n254 ;
  assign n256 = n21 & ~n255 ;
  assign n257 = ~x4 & x5 ;
  assign n258 = ~x1 & n257 ;
  assign n259 = ~x9 & n258 ;
  assign n260 = ~n256 & ~n259 ;
  assign n261 = n171 & ~n260 ;
  assign n262 = x0 & x1 ;
  assign n263 = ~x5 & n262 ;
  assign n264 = n72 & n263 ;
  assign n265 = ~n261 & ~n264 ;
  assign n266 = x3 & ~n265 ;
  assign n267 = n252 & ~n266 ;
  assign n268 = ~n243 & n267 ;
  assign n269 = ~x8 & ~n268 ;
  assign n270 = n170 & n193 ;
  assign n271 = x1 & ~x2 ;
  assign n272 = x9 & n271 ;
  assign n273 = n270 & n272 ;
  assign n274 = ~x3 & ~x4 ;
  assign n275 = n26 & n59 ;
  assign n276 = n274 & n275 ;
  assign n277 = n65 & n84 ;
  assign n278 = n277 ^ x3 ;
  assign n279 = n278 ^ n277 ;
  assign n280 = n279 ^ x8 ;
  assign n281 = n59 & n249 ;
  assign n282 = ~n11 & ~n253 ;
  assign n283 = n57 & ~n282 ;
  assign n284 = n41 & ~n271 ;
  assign n285 = ~n255 & n284 ;
  assign n286 = ~n283 & ~n285 ;
  assign n287 = ~x9 & ~n286 ;
  assign n288 = n287 ^ n281 ;
  assign n289 = ~n281 & n288 ;
  assign n290 = n289 ^ n277 ;
  assign n291 = n290 ^ n281 ;
  assign n292 = n280 & n291 ;
  assign n293 = n292 ^ n289 ;
  assign n294 = n293 ^ n281 ;
  assign n295 = x8 & ~n294 ;
  assign n296 = n295 ^ x8 ;
  assign n297 = ~n276 & ~n296 ;
  assign n298 = ~n273 & n297 ;
  assign n299 = ~n269 & n298 ;
  assign n300 = n299 ^ n212 ;
  assign n301 = ~n214 & n300 ;
  assign n302 = n301 ^ n212 ;
  assign n303 = ~n69 & n302 ;
  assign n304 = ~n55 & n303 ;
  assign n305 = n304 ^ x6 ;
  assign n306 = n305 ^ n304 ;
  assign n307 = ~x4 & x7 ;
  assign n308 = n133 & n307 ;
  assign n309 = x7 & n73 ;
  assign n310 = ~x7 & ~x8 ;
  assign n311 = x3 & ~x4 ;
  assign n312 = n310 & n311 ;
  assign n313 = ~n309 & ~n312 ;
  assign n314 = n271 & ~n313 ;
  assign n315 = ~n308 & ~n314 ;
  assign n317 = ~n132 & ~n170 ;
  assign n318 = n74 & n254 ;
  assign n319 = ~n317 & n318 ;
  assign n316 = x8 ^ x7 ;
  assign n320 = n319 ^ n316 ;
  assign n321 = n319 ^ x8 ;
  assign n322 = n321 ^ x8 ;
  assign n323 = n322 ^ n320 ;
  assign n324 = ~x1 & ~x9 ;
  assign n325 = x2 & n324 ;
  assign n326 = n325 ^ n311 ;
  assign n327 = n325 & n326 ;
  assign n328 = n327 ^ x8 ;
  assign n329 = n328 ^ n325 ;
  assign n330 = ~n323 & n329 ;
  assign n331 = n330 ^ n327 ;
  assign n332 = n331 ^ n325 ;
  assign n333 = n320 & n332 ;
  assign n334 = n333 ^ n319 ;
  assign n335 = n315 & ~n334 ;
  assign n336 = n193 & ~n335 ;
  assign n337 = n59 & n131 ;
  assign n338 = x7 ^ x3 ;
  assign n339 = n338 ^ x8 ;
  assign n340 = n72 ^ x7 ;
  assign n341 = n340 ^ n72 ;
  assign n342 = x8 ^ x4 ;
  assign n343 = n342 ^ n72 ;
  assign n344 = n341 & ~n343 ;
  assign n345 = n344 ^ n72 ;
  assign n346 = n339 & n345 ;
  assign n347 = n337 & n346 ;
  assign n348 = x7 & x8 ;
  assign n349 = n86 & n348 ;
  assign n350 = n112 & n349 ;
  assign n374 = x5 & ~x8 ;
  assign n375 = ~n63 & ~n374 ;
  assign n376 = x2 & ~n375 ;
  assign n377 = n317 & n376 ;
  assign n378 = ~x5 & ~n63 ;
  assign n379 = ~n170 & ~n311 ;
  assign n380 = n379 ^ x2 ;
  assign n381 = n378 & n380 ;
  assign n382 = ~n377 & ~n381 ;
  assign n383 = x7 & ~n382 ;
  assign n351 = ~x7 & n132 ;
  assign n352 = x5 ^ x4 ;
  assign n353 = n351 & ~n352 ;
  assign n356 = n310 ^ x5 ;
  assign n357 = n356 ^ x2 ;
  assign n361 = n357 ^ n310 ;
  assign n354 = x4 ^ x2 ;
  assign n355 = n354 ^ x2 ;
  assign n358 = n357 ^ x2 ;
  assign n359 = n358 ^ n310 ;
  assign n360 = ~n355 & n359 ;
  assign n362 = n361 ^ n360 ;
  assign n363 = n362 ^ n15 ;
  assign n364 = n348 ^ n310 ;
  assign n365 = n361 ^ n15 ;
  assign n366 = n364 & ~n365 ;
  assign n367 = n366 ^ n360 ;
  assign n368 = n367 ^ n310 ;
  assign n369 = n368 ^ n364 ;
  assign n370 = n369 ^ n361 ;
  assign n371 = n15 & ~n370 ;
  assign n372 = ~n363 & n371 ;
  assign n373 = ~n353 & ~n372 ;
  assign n384 = n383 ^ n373 ;
  assign n385 = n384 ^ n373 ;
  assign n386 = ~x8 & n76 ;
  assign n387 = n257 & n386 ;
  assign n388 = n387 ^ n373 ;
  assign n389 = n388 ^ n373 ;
  assign n390 = ~n385 & ~n389 ;
  assign n391 = n390 ^ n373 ;
  assign n392 = x1 & n391 ;
  assign n393 = n392 ^ n373 ;
  assign n394 = ~n350 & n393 ;
  assign n395 = x0 & ~n394 ;
  assign n396 = ~n63 & ~n348 ;
  assign n397 = ~n76 & ~n396 ;
  assign n398 = x2 & ~n374 ;
  assign n399 = x3 & ~n139 ;
  assign n400 = ~n398 & n399 ;
  assign n401 = ~n397 & ~n400 ;
  assign n402 = ~x4 & n310 ;
  assign n403 = ~n84 & ~n112 ;
  assign n404 = ~n402 & n403 ;
  assign n405 = x1 & ~x7 ;
  assign n406 = n405 ^ x0 ;
  assign n407 = n405 ^ x5 ;
  assign n408 = n407 ^ x5 ;
  assign n409 = ~n356 & ~n408 ;
  assign n410 = n409 ^ x5 ;
  assign n411 = n406 & ~n410 ;
  assign n412 = n411 ^ x0 ;
  assign n413 = ~n64 & ~n412 ;
  assign n414 = n404 & n413 ;
  assign n415 = n401 & n414 ;
  assign n416 = ~n395 & ~n415 ;
  assign n417 = n416 ^ x9 ;
  assign n418 = n417 ^ n416 ;
  assign n419 = n97 & n405 ;
  assign n420 = ~x1 & ~x5 ;
  assign n421 = ~x7 & x8 ;
  assign n422 = n421 ^ x2 ;
  assign n423 = n422 ^ n421 ;
  assign n424 = n423 ^ n420 ;
  assign n425 = n307 ^ x8 ;
  assign n426 = ~x8 & n425 ;
  assign n427 = n426 ^ n421 ;
  assign n428 = n427 ^ x8 ;
  assign n429 = n424 & ~n428 ;
  assign n430 = n429 ^ n426 ;
  assign n431 = n430 ^ x8 ;
  assign n432 = n420 & ~n431 ;
  assign n433 = ~n419 & ~n432 ;
  assign n434 = n28 & ~n433 ;
  assign n435 = n112 ^ n76 ;
  assign n436 = n76 ^ x8 ;
  assign n437 = n436 ^ n76 ;
  assign n438 = n435 & ~n437 ;
  assign n439 = n438 ^ n76 ;
  assign n440 = n316 & n439 ;
  assign n441 = n258 & n440 ;
  assign n442 = ~n76 & ~n311 ;
  assign n443 = x5 & n348 ;
  assign n444 = n262 & n443 ;
  assign n445 = ~n442 & n444 ;
  assign n446 = ~n441 & ~n445 ;
  assign n447 = ~n434 & n446 ;
  assign n448 = n447 ^ n416 ;
  assign n449 = ~n418 & n448 ;
  assign n450 = n449 ^ n416 ;
  assign n451 = ~n347 & n450 ;
  assign n452 = ~n336 & n451 ;
  assign n453 = n452 ^ n304 ;
  assign n454 = n306 & n453 ;
  assign n455 = n454 ^ n304 ;
  assign n456 = ~n40 & n455 ;
  assign y0 = ~n456 ;
endmodule
