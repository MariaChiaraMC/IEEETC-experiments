module top( x0 , x1 , x2 , x3 , x4 , y0 );
  input x0 , x1 , x2 , x3 , x4 ;
  output y0 ;
  wire n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ;
  assign n6 = x3 ^ x1 ;
  assign n7 = n6 ^ x2 ;
  assign n8 = n7 ^ x4 ;
  assign n9 = n8 ^ n6 ;
  assign n10 = n6 ^ x3 ;
  assign n11 = n10 ^ x4 ;
  assign n12 = n11 ^ n9 ;
  assign n13 = n12 ^ x0 ;
  assign n14 = n13 ^ n7 ;
  assign n15 = n14 ^ n6 ;
  assign n16 = n15 ^ x0 ;
  assign n22 = n16 ^ x0 ;
  assign n23 = n22 ^ n9 ;
  assign n24 = n23 ^ n13 ;
  assign n25 = n9 & ~n24 ;
  assign n17 = n16 ^ n9 ;
  assign n18 = n9 ^ n6 ;
  assign n19 = n18 ^ n9 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = ~n17 & ~n20 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = n26 ^ n9 ;
  assign n28 = n27 ^ n16 ;
  assign n29 = n22 ^ n16 ;
  assign n30 = n21 ^ n18 ;
  assign n31 = n30 ^ n16 ;
  assign n32 = ~n29 & ~n31 ;
  assign n33 = n32 ^ n21 ;
  assign n34 = n33 ^ n9 ;
  assign n35 = n34 ^ n22 ;
  assign n36 = n35 ^ n13 ;
  assign n37 = ~n28 & ~n36 ;
  assign n38 = n37 ^ n32 ;
  assign n39 = n38 ^ x1 ;
  assign y0 = ~n39 ;
endmodule
