module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;
  assign n15 = x2 & x5 ;
  assign n16 = x1 & ~x12 ;
  assign n17 = ~x8 & n16 ;
  assign n18 = ~x7 & ~x9 ;
  assign n19 = x3 & ~n18 ;
  assign n20 = x4 & n19 ;
  assign n21 = ~x11 & n20 ;
  assign n22 = ~x10 & ~x13 ;
  assign n23 = n21 & n22 ;
  assign n24 = n17 & n23 ;
  assign n25 = n15 & ~n24 ;
  assign n30 = x5 ^ x2 ;
  assign n31 = ~x3 & ~x4 ;
  assign n32 = n31 ^ x2 ;
  assign n33 = n30 & n32 ;
  assign n26 = x6 ^ x2 ;
  assign n27 = n26 ^ x2 ;
  assign n28 = x2 ^ x1 ;
  assign n29 = ~n27 & ~n28 ;
  assign n34 = n33 ^ n29 ;
  assign n35 = n29 ^ x2 ;
  assign n36 = x0 & n35 ;
  assign n37 = n36 ^ n29 ;
  assign n38 = n37 ^ x2 ;
  assign n39 = n34 & n38 ;
  assign n40 = n39 ^ n29 ;
  assign n41 = n40 ^ n36 ;
  assign n42 = n41 ^ x2 ;
  assign n43 = ~n25 & n42 ;
  assign y0 = n43 ;
endmodule
