module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 ;
  assign n17 = ~x3 & ~x7 ;
  assign n18 = ~x5 & ~n17 ;
  assign n19 = x5 & x7 ;
  assign n20 = ~x3 & ~n19 ;
  assign n21 = x10 ^ x9 ;
  assign n22 = ~n20 & ~n21 ;
  assign n23 = ~x8 & ~n22 ;
  assign n24 = ~x9 & ~x10 ;
  assign n25 = x15 ^ x14 ;
  assign n26 = n25 ^ x13 ;
  assign n27 = x15 ^ x13 ;
  assign n28 = ~x11 & ~x12 ;
  assign n29 = n28 ^ x13 ;
  assign n30 = x13 & n29 ;
  assign n31 = n30 ^ x13 ;
  assign n32 = n27 & n31 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ x13 ;
  assign n35 = n34 ^ n28 ;
  assign n36 = n26 & n35 ;
  assign n37 = ~n24 & ~n36 ;
  assign n38 = n23 & ~n37 ;
  assign n39 = ~n18 & ~n38 ;
  assign n40 = ~x6 & ~x7 ;
  assign n41 = n24 ^ n22 ;
  assign n42 = ~x8 & ~n41 ;
  assign n43 = n42 ^ n24 ;
  assign n44 = n40 & n43 ;
  assign n45 = x3 & ~n44 ;
  assign n46 = ~x0 & x1 ;
  assign n47 = x5 & ~x6 ;
  assign n48 = ~x2 & ~n47 ;
  assign n49 = n46 & n48 ;
  assign n50 = ~n45 & n49 ;
  assign n51 = ~n39 & n50 ;
  assign n52 = x0 & ~x3 ;
  assign n53 = ~x1 & n52 ;
  assign n54 = ~n51 & ~n53 ;
  assign n55 = ~x4 & ~n54 ;
  assign y0 = n55 ;
endmodule
