module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 ;
  assign n30 = x4 & ~x5 ;
  assign n31 = x1 & ~n30 ;
  assign n32 = x6 & x8 ;
  assign n33 = x7 & n32 ;
  assign n17 = ~x4 & x5 ;
  assign n34 = ~n17 & ~n30 ;
  assign n35 = n33 & ~n34 ;
  assign n36 = ~n31 & n35 ;
  assign n37 = x5 & x6 ;
  assign n38 = ~x2 & x4 ;
  assign n39 = n37 & n38 ;
  assign n40 = x2 & ~x6 ;
  assign n41 = n34 & n40 ;
  assign n42 = ~n39 & ~n41 ;
  assign n43 = ~x8 & ~n42 ;
  assign n44 = ~n36 & ~n43 ;
  assign n12 = ~x7 & x8 ;
  assign n101 = ~x2 & ~n12 ;
  assign n45 = x4 & x6 ;
  assign n92 = ~x5 & ~x8 ;
  assign n102 = x2 & ~n92 ;
  assign n103 = n45 & ~n102 ;
  assign n104 = ~n101 & n103 ;
  assign n74 = ~x5 & x7 ;
  assign n105 = x2 & ~n74 ;
  assign n88 = ~x4 & ~x6 ;
  assign n106 = n88 ^ x5 ;
  assign n107 = n88 ^ x7 ;
  assign n108 = n107 ^ x7 ;
  assign n109 = x1 & ~x2 ;
  assign n110 = n109 ^ x7 ;
  assign n111 = ~n108 & ~n110 ;
  assign n112 = n111 ^ x7 ;
  assign n113 = ~n106 & n112 ;
  assign n114 = n113 ^ x5 ;
  assign n115 = x8 & ~n114 ;
  assign n116 = ~n105 & n115 ;
  assign n117 = ~n104 & ~n116 ;
  assign n68 = x4 & x7 ;
  assign n22 = ~x6 & x8 ;
  assign n118 = x2 & ~x4 ;
  assign n119 = ~n22 & ~n118 ;
  assign n120 = ~n68 & ~n119 ;
  assign n121 = ~n33 & ~n120 ;
  assign n122 = n121 ^ x1 ;
  assign n123 = n122 ^ n121 ;
  assign n124 = n123 ^ x5 ;
  assign n65 = x4 & ~x7 ;
  assign n125 = x8 & n65 ;
  assign n126 = x8 ^ x2 ;
  assign n127 = x8 ^ x7 ;
  assign n128 = x8 ^ x6 ;
  assign n129 = n128 ^ x8 ;
  assign n130 = x8 & ~n129 ;
  assign n131 = n130 ^ x8 ;
  assign n132 = ~n127 & n131 ;
  assign n133 = n132 ^ n130 ;
  assign n134 = n133 ^ x8 ;
  assign n135 = n134 ^ n128 ;
  assign n136 = n126 & ~n135 ;
  assign n137 = n136 ^ n128 ;
  assign n138 = n137 ^ n125 ;
  assign n139 = ~n125 & ~n138 ;
  assign n140 = n139 ^ n121 ;
  assign n141 = n140 ^ n125 ;
  assign n142 = ~n124 & n141 ;
  assign n143 = n142 ^ n139 ;
  assign n144 = n143 ^ n125 ;
  assign n145 = x5 & ~n144 ;
  assign n146 = n145 ^ x5 ;
  assign n147 = n117 & ~n146 ;
  assign n66 = ~n30 & ~n37 ;
  assign n67 = ~n65 & ~n66 ;
  assign n19 = ~x6 & ~x7 ;
  assign n69 = x5 & n19 ;
  assign n70 = ~n68 & ~n69 ;
  assign n71 = n70 ^ x2 ;
  assign n72 = n71 ^ n70 ;
  assign n73 = n72 ^ n67 ;
  assign n75 = x7 ^ x4 ;
  assign n76 = n75 ^ n74 ;
  assign n77 = ~n74 & ~n76 ;
  assign n78 = n77 ^ n70 ;
  assign n79 = n78 ^ n74 ;
  assign n80 = ~n73 & n79 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n81 ^ n74 ;
  assign n83 = ~n67 & ~n82 ;
  assign n84 = n83 ^ n67 ;
  assign n85 = x8 & n84 ;
  assign n46 = ~x8 & n45 ;
  assign n47 = x5 & n46 ;
  assign n48 = x4 ^ x2 ;
  assign n49 = n48 ^ x4 ;
  assign n50 = n48 ^ x6 ;
  assign n51 = n49 & n50 ;
  assign n52 = n51 ^ n48 ;
  assign n53 = n48 ^ x5 ;
  assign n54 = n53 ^ x4 ;
  assign n55 = n54 ^ x7 ;
  assign n56 = n55 ^ n52 ;
  assign n57 = n48 ^ x8 ;
  assign n58 = n55 ^ x7 ;
  assign n59 = ~n57 & n58 ;
  assign n60 = n59 ^ n48 ;
  assign n61 = n56 & ~n60 ;
  assign n62 = n61 ^ n58 ;
  assign n63 = ~n52 & n62 ;
  assign n64 = ~n47 & ~n63 ;
  assign n86 = n85 ^ n64 ;
  assign n87 = n86 ^ n64 ;
  assign n89 = ~x5 & ~x7 ;
  assign n90 = x8 & ~n89 ;
  assign n91 = n88 & ~n90 ;
  assign n93 = n38 & n92 ;
  assign n94 = ~n91 & ~n93 ;
  assign n95 = n94 ^ n64 ;
  assign n96 = n95 ^ n64 ;
  assign n97 = ~n87 & n96 ;
  assign n98 = n97 ^ n64 ;
  assign n99 = x1 & n98 ;
  assign n100 = n99 ^ n64 ;
  assign n148 = n147 ^ n100 ;
  assign n149 = n148 ^ n147 ;
  assign n150 = n92 & n118 ;
  assign n151 = n46 ^ x2 ;
  assign n152 = n151 ^ n46 ;
  assign n153 = x6 & n12 ;
  assign n154 = n153 ^ n46 ;
  assign n155 = n152 & n154 ;
  assign n156 = n155 ^ n46 ;
  assign n157 = ~n150 & ~n156 ;
  assign n158 = n157 ^ n147 ;
  assign n159 = n158 ^ n147 ;
  assign n160 = n149 & n159 ;
  assign n161 = n160 ^ n147 ;
  assign n162 = ~x3 & n161 ;
  assign n163 = n162 ^ n147 ;
  assign n164 = n44 & n163 ;
  assign n10 = ~x1 & ~x3 ;
  assign n11 = ~x2 & n10 ;
  assign n13 = n12 ^ x6 ;
  assign n14 = ~x4 & n13 ;
  assign n15 = n14 ^ x6 ;
  assign n16 = ~x5 & n15 ;
  assign n18 = n17 ^ x0 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n20 ^ n19 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n21 & n23 ;
  assign n25 = n24 ^ n19 ;
  assign n26 = ~n18 & ~n25 ;
  assign n27 = n26 ^ x0 ;
  assign n28 = ~n16 & n27 ;
  assign n29 = n11 & n28 ;
  assign n165 = n164 ^ n29 ;
  assign n166 = n165 ^ x0 ;
  assign n173 = n166 ^ n165 ;
  assign n167 = n166 ^ n68 ;
  assign n168 = n167 ^ n165 ;
  assign n169 = n68 ^ n29 ;
  assign n170 = n169 ^ n68 ;
  assign n171 = n170 ^ n168 ;
  assign n172 = ~n168 & ~n171 ;
  assign n174 = n173 ^ n172 ;
  assign n175 = n174 ^ n168 ;
  assign n176 = n165 ^ x8 ;
  assign n177 = n172 ^ n168 ;
  assign n178 = ~n176 & ~n177 ;
  assign n179 = n178 ^ n165 ;
  assign n180 = n175 & ~n179 ;
  assign n181 = n180 ^ n165 ;
  assign n182 = n181 ^ n29 ;
  assign n183 = n182 ^ n165 ;
  assign y0 = n183 ;
endmodule
