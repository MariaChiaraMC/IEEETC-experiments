module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ;
  assign n8 = x5 & x6 ;
  assign n9 = ~x0 & n8 ;
  assign n10 = x3 ^ x2 ;
  assign n11 = n8 ^ x3 ;
  assign n12 = n11 ^ n8 ;
  assign n13 = n12 ^ n10 ;
  assign n14 = x5 ^ x0 ;
  assign n15 = ~x5 & ~n14 ;
  assign n16 = n15 ^ n8 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = ~n13 & ~n17 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n19 ^ x5 ;
  assign n21 = n10 & ~n20 ;
  assign n22 = n21 ^ x1 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = x2 & ~x3 ;
  assign n25 = n24 ^ x3 ;
  assign n26 = n25 ^ x3 ;
  assign n27 = x6 ^ x3 ;
  assign n28 = n27 ^ x3 ;
  assign n29 = n26 & n28 ;
  assign n30 = n29 ^ x3 ;
  assign n31 = x5 & n30 ;
  assign n32 = n31 ^ x3 ;
  assign n33 = n32 ^ n21 ;
  assign n34 = n23 & n33 ;
  assign n35 = n34 ^ n21 ;
  assign n36 = ~n9 & ~n35 ;
  assign n37 = ~x4 & ~n36 ;
  assign n38 = ~x5 & ~x6 ;
  assign n39 = ~n37 & ~n38 ;
  assign y0 = ~n39 ;
endmodule
