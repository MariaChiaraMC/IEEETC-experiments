module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 ;
  assign n11 = ~x1 & x9 ;
  assign n12 = ~x8 & ~n11 ;
  assign n13 = ~x4 & ~x5 ;
  assign n14 = n13 ^ x3 ;
  assign n15 = x9 & ~n14 ;
  assign n16 = n15 ^ x3 ;
  assign n17 = ~n12 & ~n16 ;
  assign n18 = x7 & ~n17 ;
  assign n19 = ~x1 & ~x3 ;
  assign n20 = n19 ^ x7 ;
  assign n21 = n20 ^ x7 ;
  assign n22 = x9 ^ x7 ;
  assign n23 = n21 & ~n22 ;
  assign n24 = n23 ^ x7 ;
  assign n25 = x8 & ~n24 ;
  assign n26 = ~n18 & ~n25 ;
  assign y0 = ~n26 ;
endmodule
