module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
  assign n9 = x2 & x3 ;
  assign n10 = x1 & n9 ;
  assign n11 = x0 & ~n10 ;
  assign n12 = x4 & ~n11 ;
  assign n18 = x6 ^ x3 ;
  assign n19 = x6 ^ x2 ;
  assign n20 = n19 ^ x6 ;
  assign n21 = n18 & n20 ;
  assign n13 = x6 ^ x5 ;
  assign n23 = n21 ^ n13 ;
  assign n14 = n13 ^ x6 ;
  assign n15 = x6 ^ x1 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n14 & ~n16 ;
  assign n24 = n17 ^ n13 ;
  assign n25 = n24 ^ n14 ;
  assign n26 = n25 ^ x7 ;
  assign n27 = ~n23 & ~n26 ;
  assign n22 = n21 ^ n17 ;
  assign n28 = n27 ^ n22 ;
  assign n29 = x7 & n28 ;
  assign n30 = n29 ^ n17 ;
  assign n31 = n30 ^ n21 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = n32 ^ x7 ;
  assign n34 = n33 ^ x7 ;
  assign n35 = ~n12 & n34 ;
  assign y0 = n35 ;
endmodule
