module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 ;
  assign n9 = x0 & ~x6 ;
  assign n10 = ~x1 & ~x4 ;
  assign n11 = x2 & n10 ;
  assign n12 = n9 & n11 ;
  assign n13 = x3 & n12 ;
  assign n22 = x4 & x6 ;
  assign n18 = ~x0 & ~x7 ;
  assign n81 = ~x1 & ~x3 ;
  assign n82 = n18 & n81 ;
  assign n83 = n22 & n82 ;
  assign n88 = x7 ^ x4 ;
  assign n84 = x4 ^ x3 ;
  assign n85 = n84 ^ x0 ;
  assign n86 = n85 ^ x1 ;
  assign n87 = n86 ^ x7 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = n84 ^ x6 ;
  assign n91 = n90 ^ n87 ;
  assign n92 = n91 ^ n87 ;
  assign n93 = n92 ^ n88 ;
  assign n94 = n93 ^ n84 ;
  assign n95 = n94 ^ n88 ;
  assign n96 = n95 ^ n84 ;
  assign n97 = ~n89 & n96 ;
  assign n98 = n97 ^ n84 ;
  assign n99 = n98 ^ n94 ;
  assign n100 = n88 ^ x7 ;
  assign n101 = n88 ^ x1 ;
  assign n102 = ~n100 & n101 ;
  assign n103 = n102 ^ n84 ;
  assign n104 = n103 ^ n94 ;
  assign n105 = ~n98 & n104 ;
  assign n106 = n105 ^ n84 ;
  assign n107 = n99 & ~n106 ;
  assign n108 = n107 ^ x2 ;
  assign n109 = n108 ^ n107 ;
  assign n58 = x4 & ~x7 ;
  assign n59 = ~x1 & n58 ;
  assign n110 = ~x3 & n59 ;
  assign n45 = x0 & ~x7 ;
  assign n111 = x3 & ~x4 ;
  assign n112 = n45 & n111 ;
  assign n113 = x3 & x7 ;
  assign n114 = ~x3 & x4 ;
  assign n115 = ~n111 & ~n114 ;
  assign n30 = ~x0 & x4 ;
  assign n116 = n115 ^ n30 ;
  assign n117 = n116 ^ n30 ;
  assign n118 = n30 ^ x1 ;
  assign n119 = n118 ^ n30 ;
  assign n120 = ~n117 & ~n119 ;
  assign n121 = n120 ^ n30 ;
  assign n122 = ~n113 & n121 ;
  assign n123 = n122 ^ n30 ;
  assign n124 = ~n112 & ~n123 ;
  assign n125 = n124 ^ x6 ;
  assign n126 = n125 ^ n124 ;
  assign n127 = n126 ^ n110 ;
  assign n61 = x1 & x7 ;
  assign n128 = n61 & ~n114 ;
  assign n129 = ~n58 & ~n128 ;
  assign n130 = n129 ^ x0 ;
  assign n131 = x0 & ~n130 ;
  assign n132 = n131 ^ n124 ;
  assign n133 = n132 ^ x0 ;
  assign n134 = n127 & ~n133 ;
  assign n135 = n134 ^ n131 ;
  assign n136 = n135 ^ x0 ;
  assign n137 = ~n110 & n136 ;
  assign n138 = n137 ^ n110 ;
  assign n139 = n138 ^ n107 ;
  assign n140 = n109 & n139 ;
  assign n141 = n140 ^ n107 ;
  assign n142 = ~n83 & ~n141 ;
  assign n14 = x1 & x2 ;
  assign n15 = ~x4 & ~x6 ;
  assign n16 = n15 ^ x7 ;
  assign n17 = n16 ^ x7 ;
  assign n19 = n18 ^ x7 ;
  assign n20 = ~n17 & n19 ;
  assign n21 = n20 ^ x7 ;
  assign n23 = ~x7 & n22 ;
  assign n24 = n23 ^ n14 ;
  assign n25 = ~n21 & n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n14 & n26 ;
  assign n28 = n27 ^ n14 ;
  assign n29 = x6 & ~x7 ;
  assign n31 = ~x2 & ~x4 ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = n29 & ~n32 ;
  assign n34 = x0 & x6 ;
  assign n35 = n31 & n34 ;
  assign n36 = x2 & x7 ;
  assign n37 = n9 & n36 ;
  assign n38 = ~n35 & ~n37 ;
  assign n39 = ~n33 & n38 ;
  assign n40 = n39 ^ x1 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = n41 ^ n28 ;
  assign n43 = x6 & x7 ;
  assign n44 = ~x0 & n43 ;
  assign n46 = ~x2 & n45 ;
  assign n47 = ~n44 & ~n46 ;
  assign n48 = n47 ^ x4 ;
  assign n49 = ~n47 & ~n48 ;
  assign n50 = n49 ^ n39 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = ~n42 & n51 ;
  assign n53 = n52 ^ n49 ;
  assign n54 = n53 ^ n47 ;
  assign n55 = ~n28 & ~n54 ;
  assign n56 = n55 ^ n28 ;
  assign n57 = x3 & n56 ;
  assign n60 = x3 & ~n59 ;
  assign n62 = n15 & n61 ;
  assign n63 = ~n58 & ~n62 ;
  assign n64 = ~x0 & ~n63 ;
  assign n65 = x1 & x4 ;
  assign n66 = n29 & n65 ;
  assign n67 = ~n64 & ~n66 ;
  assign n68 = ~n60 & ~n67 ;
  assign n69 = n68 ^ x2 ;
  assign n70 = n69 ^ n68 ;
  assign n71 = n70 ^ n57 ;
  assign n72 = n44 ^ n10 ;
  assign n73 = n44 & n72 ;
  assign n74 = n73 ^ n68 ;
  assign n75 = n74 ^ n44 ;
  assign n76 = ~n71 & n75 ;
  assign n77 = n76 ^ n73 ;
  assign n78 = n77 ^ n44 ;
  assign n79 = ~n57 & n78 ;
  assign n80 = n79 ^ n57 ;
  assign n143 = n142 ^ n80 ;
  assign n144 = x5 & ~n143 ;
  assign n145 = n144 ^ n142 ;
  assign n146 = ~n13 & n145 ;
  assign y0 = ~n146 ;
endmodule
