module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 ;
  assign n8 = ~x5 & ~x6 ;
  assign n9 = ~x4 & n8 ;
  assign n10 = x3 & ~n9 ;
  assign n11 = x5 ^ x4 ;
  assign n12 = x6 ^ x5 ;
  assign n13 = n11 & ~n12 ;
  assign n14 = n13 ^ x4 ;
  assign n15 = ~n10 & ~n14 ;
  assign n16 = x5 & x6 ;
  assign n17 = x4 & n16 ;
  assign n18 = x3 & n14 ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = ~x2 & n19 ;
  assign n21 = ~n15 & ~n20 ;
  assign n22 = n21 ^ x1 ;
  assign n23 = n17 ^ x2 ;
  assign n24 = n23 ^ x0 ;
  assign n25 = n18 ^ x3 ;
  assign n26 = ~x2 & ~n25 ;
  assign n27 = n26 ^ n18 ;
  assign n28 = ~n24 & ~n27 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = n29 ^ n18 ;
  assign n31 = n30 ^ x2 ;
  assign n32 = ~x0 & n31 ;
  assign n33 = n32 ^ n21 ;
  assign n34 = n33 ^ n32 ;
  assign n35 = n9 ^ x3 ;
  assign n36 = n9 ^ x2 ;
  assign n37 = n36 ^ n9 ;
  assign n38 = n14 ^ n9 ;
  assign n39 = n38 ^ n9 ;
  assign n40 = ~n37 & ~n39 ;
  assign n41 = n40 ^ n9 ;
  assign n42 = ~n35 & ~n41 ;
  assign n43 = n42 ^ x3 ;
  assign n44 = ~n32 & n43 ;
  assign n45 = n44 ^ n32 ;
  assign n46 = ~n34 & n45 ;
  assign n47 = n46 ^ n32 ;
  assign n48 = n22 & ~n47 ;
  assign n49 = n48 ^ x1 ;
  assign y0 = n49 ;
endmodule
