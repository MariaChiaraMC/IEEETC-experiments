module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 ;
  assign n12 = x3 ^ x2 ;
  assign n13 = n12 ^ x5 ;
  assign n14 = n13 ^ x2 ;
  assign n9 = x5 ^ x4 ;
  assign n10 = n9 ^ x2 ;
  assign n11 = n10 ^ x2 ;
  assign n15 = n14 ^ n11 ;
  assign n23 = n13 ^ x6 ;
  assign n24 = n23 ^ n9 ;
  assign n17 = x5 ^ x2 ;
  assign n18 = n17 ^ n13 ;
  assign n25 = n24 ^ n18 ;
  assign n19 = n18 ^ n9 ;
  assign n20 = n19 ^ n13 ;
  assign n21 = n20 ^ x2 ;
  assign n16 = n11 ^ n10 ;
  assign n22 = n21 ^ n16 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = ~n15 & n26 ;
  assign n28 = n27 ^ n10 ;
  assign n29 = n28 ^ n14 ;
  assign n30 = n21 ^ n14 ;
  assign n31 = n25 & n30 ;
  assign n32 = n31 ^ n14 ;
  assign n33 = n32 ^ n11 ;
  assign n34 = n13 ^ x7 ;
  assign n35 = n34 ^ n18 ;
  assign n36 = n35 ^ n14 ;
  assign n37 = n36 ^ n11 ;
  assign n38 = ~n21 & n37 ;
  assign n39 = n38 ^ n10 ;
  assign n40 = n39 ^ n14 ;
  assign n41 = n40 ^ n11 ;
  assign n42 = ~n33 & n41 ;
  assign n43 = n42 ^ n10 ;
  assign n44 = n43 ^ n14 ;
  assign n45 = n44 ^ n11 ;
  assign n46 = n29 & n45 ;
  assign n47 = n46 ^ x2 ;
  assign y0 = ~n47 ;
endmodule
