module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 ;
  assign n25 = x2 & ~x6 ;
  assign n26 = ~x3 & n25 ;
  assign n76 = x1 & ~x4 ;
  assign n77 = n26 & n76 ;
  assign n22 = x2 & x4 ;
  assign n23 = x6 & n22 ;
  assign n24 = x3 & n23 ;
  assign n27 = ~x2 & x6 ;
  assign n78 = x3 & n27 ;
  assign n79 = x1 & x3 ;
  assign n80 = x6 & n79 ;
  assign n81 = ~n78 & ~n80 ;
  assign n82 = ~x4 & ~n81 ;
  assign n83 = ~n24 & ~n82 ;
  assign n84 = ~n77 & n83 ;
  assign n85 = x7 & ~n84 ;
  assign n9 = x3 & ~x4 ;
  assign n86 = x1 & ~x7 ;
  assign n87 = ~n9 & ~n86 ;
  assign n88 = ~x2 & ~x6 ;
  assign n89 = ~n79 & n88 ;
  assign n90 = ~n87 & n89 ;
  assign n91 = ~x0 & ~n90 ;
  assign n92 = ~n85 & n91 ;
  assign n94 = x6 ^ x4 ;
  assign n10 = x3 ^ x2 ;
  assign n99 = n94 ^ n10 ;
  assign n100 = n99 ^ n94 ;
  assign n93 = x4 ^ x1 ;
  assign n95 = n94 ^ n93 ;
  assign n96 = n95 ^ x4 ;
  assign n97 = n96 ^ x3 ;
  assign n98 = n97 ^ n94 ;
  assign n101 = n100 ^ n98 ;
  assign n104 = n97 ^ x3 ;
  assign n102 = x4 ^ x3 ;
  assign n103 = n102 ^ n98 ;
  assign n105 = n104 ^ n103 ;
  assign n106 = n101 & ~n105 ;
  assign n107 = n106 ^ n97 ;
  assign n108 = n107 ^ n102 ;
  assign n109 = n108 ^ n104 ;
  assign n110 = n103 ^ n100 ;
  assign n111 = n107 & ~n110 ;
  assign n112 = n111 ^ n97 ;
  assign n113 = n112 ^ n98 ;
  assign n114 = n113 ^ n100 ;
  assign n115 = n109 & n114 ;
  assign n116 = n115 ^ x7 ;
  assign n117 = n116 ^ n115 ;
  assign n118 = ~n25 & ~n78 ;
  assign n119 = ~x1 & x4 ;
  assign n120 = ~n118 & n119 ;
  assign n121 = ~n10 & n76 ;
  assign n122 = n121 ^ x6 ;
  assign n123 = n122 ^ n121 ;
  assign n124 = n123 ^ n120 ;
  assign n125 = n79 ^ x4 ;
  assign n126 = n79 & n125 ;
  assign n127 = n126 ^ n121 ;
  assign n128 = n127 ^ n79 ;
  assign n129 = n124 & n128 ;
  assign n130 = n129 ^ n126 ;
  assign n131 = n130 ^ n79 ;
  assign n132 = ~n120 & n131 ;
  assign n133 = n132 ^ n120 ;
  assign n134 = n133 ^ n115 ;
  assign n135 = ~n117 & n134 ;
  assign n136 = n135 ^ n115 ;
  assign n137 = x0 & ~n136 ;
  assign n138 = ~n92 & ~n137 ;
  assign n11 = ~n9 & ~n10 ;
  assign n12 = ~x6 & n11 ;
  assign n13 = n12 ^ x1 ;
  assign n14 = n13 ^ x0 ;
  assign n20 = n14 ^ n13 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n15 ^ x7 ;
  assign n17 = n14 ^ x7 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = n16 & n18 ;
  assign n21 = n20 ^ n19 ;
  assign n28 = ~x4 & n27 ;
  assign n29 = ~n26 & ~n28 ;
  assign n30 = ~n24 & n29 ;
  assign n31 = n30 ^ n14 ;
  assign n32 = ~n20 & ~n31 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = ~n21 & n33 ;
  assign n35 = n34 ^ n19 ;
  assign n36 = n35 ^ n14 ;
  assign n37 = n36 ^ x1 ;
  assign n38 = n37 ^ n13 ;
  assign n39 = n38 ^ x1 ;
  assign n40 = x2 & x3 ;
  assign n41 = x0 & ~n40 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = n42 ^ n39 ;
  assign n47 = x4 & ~x6 ;
  assign n48 = x7 & n47 ;
  assign n64 = x2 & ~x3 ;
  assign n65 = ~x0 & ~n64 ;
  assign n66 = n48 & ~n65 ;
  assign n44 = x7 ^ x3 ;
  assign n45 = n44 ^ x7 ;
  assign n46 = n45 ^ n9 ;
  assign n49 = x6 & ~x7 ;
  assign n50 = ~x4 & n49 ;
  assign n51 = ~n48 & ~n50 ;
  assign n52 = x2 & ~n51 ;
  assign n53 = ~x2 & ~x4 ;
  assign n54 = ~n49 & n53 ;
  assign n55 = n54 ^ n52 ;
  assign n56 = ~n52 & n55 ;
  assign n57 = n56 ^ x7 ;
  assign n58 = n57 ^ n52 ;
  assign n59 = n46 & n58 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = n60 ^ n52 ;
  assign n62 = ~n9 & ~n61 ;
  assign n63 = n62 ^ n9 ;
  assign n67 = n66 ^ n63 ;
  assign n68 = n38 & ~n67 ;
  assign n69 = n68 ^ n63 ;
  assign n70 = n43 & ~n69 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = n71 ^ n63 ;
  assign n73 = n72 ^ n38 ;
  assign n74 = n39 & ~n73 ;
  assign n75 = n74 ^ x1 ;
  assign n139 = n138 ^ n75 ;
  assign n140 = n139 ^ n75 ;
  assign n141 = n47 & n86 ;
  assign n142 = n40 & n141 ;
  assign n143 = n142 ^ n75 ;
  assign n144 = n143 ^ n75 ;
  assign n145 = ~n140 & ~n144 ;
  assign n146 = n145 ^ n75 ;
  assign n147 = x5 & n146 ;
  assign n148 = n147 ^ n75 ;
  assign y0 = ~n148 ;
endmodule
