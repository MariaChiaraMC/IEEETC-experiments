module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 ;
  assign n17 = x4 & x8 ;
  assign n40 = ~x7 & ~n17 ;
  assign n42 = x6 ^ x3 ;
  assign n41 = x7 ^ x3 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = n43 ^ x8 ;
  assign n45 = n44 ^ n43 ;
  assign n46 = n45 ^ x3 ;
  assign n47 = n43 ^ n42 ;
  assign n48 = n47 ^ x3 ;
  assign n49 = n48 ^ n42 ;
  assign n50 = n49 ^ x3 ;
  assign n51 = n50 ^ n48 ;
  assign n52 = ~n46 & ~n51 ;
  assign n53 = n52 ^ n45 ;
  assign n54 = n43 ^ x2 ;
  assign n55 = n54 ^ n44 ;
  assign n56 = n43 ^ x4 ;
  assign n57 = n56 ^ n44 ;
  assign n58 = n55 & n57 ;
  assign n59 = n58 ^ n45 ;
  assign n60 = n53 ^ n48 ;
  assign n61 = n59 & ~n60 ;
  assign n62 = n61 ^ n50 ;
  assign n63 = n62 ^ n48 ;
  assign n64 = n53 & ~n63 ;
  assign n65 = n64 ^ n45 ;
  assign n66 = n65 ^ n46 ;
  assign n67 = n66 ^ x6 ;
  assign n68 = n67 ^ x3 ;
  assign n69 = ~n40 & n68 ;
  assign n70 = x0 & ~n69 ;
  assign n71 = x6 & x8 ;
  assign n72 = ~x1 & ~n71 ;
  assign n73 = ~n70 & ~n72 ;
  assign n10 = x2 & x6 ;
  assign n11 = x1 & ~n10 ;
  assign n12 = x6 ^ x4 ;
  assign n13 = x8 ^ x6 ;
  assign n14 = n12 & ~n13 ;
  assign n15 = n14 ^ x4 ;
  assign n16 = n11 & ~n15 ;
  assign n18 = ~x1 & x2 ;
  assign n19 = n17 & n18 ;
  assign n20 = ~n16 & ~n19 ;
  assign n21 = ~x7 & ~n20 ;
  assign n22 = x4 & x6 ;
  assign n23 = x8 & n22 ;
  assign n24 = n23 ^ x0 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = ~x6 & ~x7 ;
  assign n28 = ~x2 & ~n17 ;
  assign n29 = ~n22 & n28 ;
  assign n30 = ~n27 & ~n29 ;
  assign n31 = n30 ^ x1 ;
  assign n32 = ~x1 & n31 ;
  assign n33 = n32 ^ n23 ;
  assign n34 = n33 ^ x1 ;
  assign n35 = ~n26 & ~n34 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ x1 ;
  assign n38 = ~n21 & ~n37 ;
  assign n39 = n38 ^ n21 ;
  assign n74 = n73 ^ n39 ;
  assign n75 = n74 ^ x3 ;
  assign n85 = n75 ^ n74 ;
  assign n76 = x4 & x7 ;
  assign n77 = ~x0 & x1 ;
  assign n78 = ~n76 & ~n77 ;
  assign n79 = n78 ^ n75 ;
  assign n80 = n79 ^ n74 ;
  assign n81 = n78 ^ n73 ;
  assign n82 = n81 ^ n78 ;
  assign n83 = n82 ^ n80 ;
  assign n84 = n80 & n83 ;
  assign n86 = n85 ^ n84 ;
  assign n87 = n86 ^ n80 ;
  assign n88 = n74 ^ n11 ;
  assign n89 = n84 ^ n80 ;
  assign n90 = ~n88 & n89 ;
  assign n91 = n90 ^ n74 ;
  assign n92 = n87 & n91 ;
  assign n93 = n92 ^ n74 ;
  assign n94 = n93 ^ n73 ;
  assign n95 = n94 ^ n74 ;
  assign n96 = x5 & n95 ;
  assign n97 = ~x4 & x5 ;
  assign n98 = x2 & n97 ;
  assign n101 = x4 ^ x0 ;
  assign n105 = n101 ^ x4 ;
  assign n99 = x6 ^ x2 ;
  assign n100 = n99 ^ x6 ;
  assign n102 = n101 ^ x6 ;
  assign n103 = n102 ^ x4 ;
  assign n104 = ~n100 & ~n103 ;
  assign n106 = n105 ^ n104 ;
  assign n107 = ~x5 & ~x7 ;
  assign n108 = n107 ^ x4 ;
  assign n109 = ~n105 & n108 ;
  assign n110 = n109 ^ n107 ;
  assign n111 = ~n106 & n110 ;
  assign n112 = n111 ^ x4 ;
  assign n113 = n112 ^ x4 ;
  assign n114 = ~n98 & ~n113 ;
  assign n115 = n114 ^ x5 ;
  assign n116 = n115 ^ n114 ;
  assign n117 = n114 ^ n10 ;
  assign n118 = n117 ^ n114 ;
  assign n119 = ~n116 & n118 ;
  assign n120 = n119 ^ n114 ;
  assign n121 = ~x8 & ~n120 ;
  assign n122 = n121 ^ n114 ;
  assign n123 = x1 & ~n122 ;
  assign n124 = ~x2 & ~x6 ;
  assign n125 = ~x1 & ~x5 ;
  assign n126 = ~x0 & ~n125 ;
  assign n127 = ~n124 & n126 ;
  assign n128 = n13 ^ x6 ;
  assign n129 = n128 ^ n97 ;
  assign n130 = n18 ^ x6 ;
  assign n131 = ~n129 & n130 ;
  assign n132 = n131 ^ n18 ;
  assign n133 = n97 & n132 ;
  assign n134 = ~n127 & ~n133 ;
  assign n135 = x2 & ~x8 ;
  assign n136 = n22 & ~n135 ;
  assign n137 = n125 & n136 ;
  assign n138 = x0 & n137 ;
  assign n139 = ~x4 & x8 ;
  assign n140 = x1 & ~n139 ;
  assign n141 = x0 & ~x5 ;
  assign n142 = n141 ^ x4 ;
  assign n143 = n142 ^ n141 ;
  assign n144 = n143 ^ n140 ;
  assign n145 = x5 & x8 ;
  assign n146 = n124 & n145 ;
  assign n147 = n146 ^ n135 ;
  assign n148 = ~n146 & n147 ;
  assign n149 = n148 ^ n141 ;
  assign n150 = n149 ^ n146 ;
  assign n151 = n144 & n150 ;
  assign n152 = n151 ^ n148 ;
  assign n153 = n152 ^ n146 ;
  assign n154 = n140 & ~n153 ;
  assign n155 = n154 ^ n140 ;
  assign n156 = ~n138 & ~n155 ;
  assign n157 = x8 & n18 ;
  assign n158 = n141 & n157 ;
  assign n159 = ~x6 & n158 ;
  assign n160 = n156 & ~n159 ;
  assign n161 = n134 & n160 ;
  assign n162 = x7 & ~n161 ;
  assign n163 = ~n123 & ~n162 ;
  assign n164 = x3 & ~n163 ;
  assign n165 = x1 & ~x5 ;
  assign n176 = ~x6 & ~x8 ;
  assign n166 = x3 ^ x0 ;
  assign n167 = n166 ^ n23 ;
  assign n168 = n167 ^ x3 ;
  assign n177 = n176 ^ n168 ;
  assign n181 = n177 ^ n167 ;
  assign n182 = n181 ^ n166 ;
  assign n169 = n168 ^ n167 ;
  assign n170 = n169 ^ n166 ;
  assign n171 = n170 ^ n166 ;
  assign n172 = ~x4 & ~x6 ;
  assign n173 = n172 ^ n167 ;
  assign n174 = n173 ^ n166 ;
  assign n175 = n171 & n174 ;
  assign n178 = n177 ^ n175 ;
  assign n179 = n178 ^ n166 ;
  assign n180 = ~n170 & ~n179 ;
  assign n183 = n182 ^ n180 ;
  assign n184 = n183 ^ n170 ;
  assign n185 = n166 ^ x2 ;
  assign n186 = n182 ^ n179 ;
  assign n187 = n186 ^ n170 ;
  assign n188 = ~n185 & ~n187 ;
  assign n189 = n188 ^ n166 ;
  assign n190 = n184 & ~n189 ;
  assign n191 = n190 ^ n188 ;
  assign n192 = n191 ^ n166 ;
  assign n193 = n192 ^ x0 ;
  assign n194 = n165 & ~n193 ;
  assign n219 = n194 ^ x7 ;
  assign n228 = n219 ^ n194 ;
  assign n195 = n126 & ~n176 ;
  assign n196 = ~x5 & ~x6 ;
  assign n197 = x0 & ~n196 ;
  assign n198 = ~x5 & ~x8 ;
  assign n199 = x7 & ~n198 ;
  assign n200 = ~n145 & ~n199 ;
  assign n201 = n22 & ~n200 ;
  assign n202 = n197 & ~n201 ;
  assign n203 = n40 ^ x3 ;
  assign n204 = n140 ^ n40 ;
  assign n205 = n204 ^ n140 ;
  assign n206 = n205 ^ n203 ;
  assign n207 = n125 ^ x4 ;
  assign n208 = ~n125 & n207 ;
  assign n209 = n208 ^ n140 ;
  assign n210 = n209 ^ n125 ;
  assign n211 = ~n206 & n210 ;
  assign n212 = n211 ^ n208 ;
  assign n213 = n212 ^ n125 ;
  assign n214 = ~n203 & ~n213 ;
  assign n215 = n214 ^ n40 ;
  assign n216 = n202 & n215 ;
  assign n217 = ~n195 & ~n216 ;
  assign n218 = n217 ^ n194 ;
  assign n220 = n219 ^ n218 ;
  assign n221 = n220 ^ n219 ;
  assign n222 = n221 ^ n194 ;
  assign n223 = x2 & ~n172 ;
  assign n224 = n223 ^ n220 ;
  assign n225 = n224 ^ n220 ;
  assign n226 = n225 ^ n222 ;
  assign n227 = ~n222 & ~n226 ;
  assign n229 = n228 ^ n227 ;
  assign n230 = n229 ^ n222 ;
  assign n231 = n194 ^ x6 ;
  assign n232 = n227 ^ n222 ;
  assign n233 = ~n231 & ~n232 ;
  assign n234 = n233 ^ n194 ;
  assign n235 = ~n230 & ~n234 ;
  assign n236 = n235 ^ n194 ;
  assign n237 = n236 ^ x7 ;
  assign n238 = n237 ^ n194 ;
  assign n239 = ~n164 & ~n238 ;
  assign n240 = ~n96 & n239 ;
  assign y0 = ~n240 ;
endmodule
