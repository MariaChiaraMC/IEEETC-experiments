module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 ;
  assign n7 = x1 ^ x0 ;
  assign n8 = n7 ^ x2 ;
  assign n10 = n8 ^ x1 ;
  assign n17 = n10 ^ x4 ;
  assign n12 = n10 ^ x2 ;
  assign n13 = n12 ^ x3 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = n18 ^ n8 ;
  assign n9 = n8 ^ x3 ;
  assign n11 = n10 ^ n9 ;
  assign n14 = n13 ^ n11 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = n15 ^ n8 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = n15 ^ n13 ;
  assign n22 = n21 ^ n10 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = ~n20 & ~n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n22 ^ n15 ;
  assign n27 = n26 ^ n21 ;
  assign n28 = n23 ^ n21 ;
  assign n29 = ~n27 & n28 ;
  assign n30 = n29 ^ n22 ;
  assign n31 = n30 ^ n19 ;
  assign n32 = n21 ^ n19 ;
  assign n33 = n13 ^ x5 ;
  assign n34 = n33 ^ n8 ;
  assign n35 = n34 ^ n8 ;
  assign n36 = n35 ^ n22 ;
  assign n37 = ~n32 & n36 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = n38 ^ n15 ;
  assign n40 = n31 & ~n39 ;
  assign n41 = n40 ^ n15 ;
  assign n42 = n25 & n41 ;
  assign n43 = n42 ^ n29 ;
  assign n44 = n43 ^ n24 ;
  assign n45 = n44 ^ n40 ;
  assign n46 = n45 ^ n15 ;
  assign n47 = n46 ^ n22 ;
  assign n48 = n47 ^ n7 ;
  assign n49 = n48 ^ n8 ;
  assign y0 = n49 ;
endmodule
