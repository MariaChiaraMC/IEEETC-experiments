module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n15 = x2 & x5 ;
  assign n16 = ~x0 & n15 ;
  assign n17 = ~x11 & ~x13 ;
  assign n18 = x8 & n17 ;
  assign n19 = x4 & ~x7 ;
  assign n20 = x1 & ~x9 ;
  assign n21 = n19 & n20 ;
  assign n22 = x6 & ~x12 ;
  assign n23 = ~x10 & n22 ;
  assign n24 = n21 & n23 ;
  assign n25 = n18 & n24 ;
  assign n26 = n25 ^ x3 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = ~x4 & ~x6 ;
  assign n29 = n28 ^ n25 ;
  assign n30 = ~n27 & n29 ;
  assign n31 = n30 ^ n25 ;
  assign n32 = n16 & n31 ;
  assign y0 = n32 ;
endmodule
