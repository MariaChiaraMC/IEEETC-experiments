// Benchmark "./pla/mish.pla_dbb_orig_7NonExact" written by ABC on Fri Nov 20 10:25:32 2020

module \./pla/mish.pla_dbb_orig_7NonExact  ( 
    x0, x1,
    z0  );
  input  x0, x1;
  output z0;
  assign z0 = x0 | ~x1;
endmodule


