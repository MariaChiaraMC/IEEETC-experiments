module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 ;
  assign n12 = x1 & x2 ;
  assign n13 = ~x7 & ~n12 ;
  assign n14 = ~x6 & ~n13 ;
  assign n15 = ~x3 & ~n14 ;
  assign n16 = x3 & x7 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = ~x8 & x9 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = ~x2 & x6 ;
  assign n23 = x3 & ~n22 ;
  assign n24 = n23 ^ x10 ;
  assign n25 = n16 & ~n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n21 & ~n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n28 ^ n23 ;
  assign n30 = n29 ^ n16 ;
  assign n31 = n17 & ~n30 ;
  assign n32 = x10 ^ x4 ;
  assign n33 = n32 ^ x4 ;
  assign n34 = n33 ^ x0 ;
  assign n35 = x6 ^ x4 ;
  assign n36 = n35 ^ x5 ;
  assign n37 = ~x5 & n36 ;
  assign n38 = n37 ^ x4 ;
  assign n39 = n38 ^ x5 ;
  assign n40 = n34 & n39 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n41 ^ x5 ;
  assign n43 = ~x0 & ~n42 ;
  assign n44 = n31 & n43 ;
  assign n45 = ~n15 & n44 ;
  assign y0 = n45 ;
endmodule
