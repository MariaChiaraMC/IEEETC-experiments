module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 ;
  assign n8 = ~x3 & ~x4 ;
  assign n9 = x1 & ~n8 ;
  assign n10 = ~x5 & ~x6 ;
  assign n11 = ~n9 & ~n10 ;
  assign n12 = x4 ^ x3 ;
  assign n13 = x3 ^ x2 ;
  assign n14 = n13 ^ x4 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = n13 ^ x0 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = ~n15 & ~n17 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = ~n12 & n19 ;
  assign n21 = n20 ^ n13 ;
  assign n22 = n11 & n21 ;
  assign y0 = n22 ;
endmodule
