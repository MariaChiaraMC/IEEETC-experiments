module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 ;
  assign n12 = x4 & x5 ;
  assign n13 = x8 & ~n12 ;
  assign n14 = ~x5 & x9 ;
  assign n15 = ~x4 & ~x5 ;
  assign n16 = ~n14 & ~n15 ;
  assign n17 = n13 & n16 ;
  assign n18 = x2 ^ x1 ;
  assign n19 = ~x4 & n18 ;
  assign n20 = ~x4 & x8 ;
  assign n21 = x5 & x9 ;
  assign n22 = ~n20 & n21 ;
  assign n23 = ~n19 & n22 ;
  assign n24 = x4 & x8 ;
  assign n25 = x5 & n18 ;
  assign n26 = ~n24 & n25 ;
  assign n27 = ~n23 & ~n26 ;
  assign n28 = ~n17 & n27 ;
  assign n29 = x1 & x4 ;
  assign n30 = n29 ^ x0 ;
  assign n31 = n20 ^ x0 ;
  assign n32 = ~x5 & ~x9 ;
  assign n33 = n32 ^ x0 ;
  assign n34 = x0 & n33 ;
  assign n35 = n34 ^ x0 ;
  assign n36 = n31 & n35 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = n37 ^ x0 ;
  assign n39 = n38 ^ n32 ;
  assign n40 = n30 & n39 ;
  assign n41 = n28 & ~n40 ;
  assign n42 = ~x10 & ~n41 ;
  assign n43 = ~x6 & ~n42 ;
  assign n44 = x5 & ~x9 ;
  assign n45 = ~x4 & ~n44 ;
  assign n46 = n13 & ~n45 ;
  assign n47 = ~x2 & ~x3 ;
  assign n48 = x5 & ~n47 ;
  assign n49 = x8 & x9 ;
  assign n50 = ~x4 & n49 ;
  assign n51 = ~n48 & n50 ;
  assign n52 = x10 & ~n51 ;
  assign n53 = ~n46 & ~n52 ;
  assign n54 = x5 & x10 ;
  assign n55 = x3 ^ x2 ;
  assign n56 = ~n54 & ~n55 ;
  assign n57 = n51 & ~n56 ;
  assign n58 = x6 & ~n57 ;
  assign n59 = x2 & x3 ;
  assign n60 = ~n47 & ~n59 ;
  assign n61 = ~x8 & ~n21 ;
  assign n62 = n61 ^ n14 ;
  assign n63 = n60 & n62 ;
  assign n64 = n63 ^ n14 ;
  assign n65 = n58 & ~n64 ;
  assign n66 = n53 & n65 ;
  assign n67 = ~x7 & ~n66 ;
  assign n68 = ~n43 & n67 ;
  assign n69 = ~x3 & ~x4 ;
  assign n70 = x3 & x4 ;
  assign n71 = ~x8 & ~x9 ;
  assign n72 = ~n70 & n71 ;
  assign n73 = ~n69 & n72 ;
  assign n74 = ~n14 & ~n46 ;
  assign n75 = ~n73 & n74 ;
  assign n76 = ~x10 & ~n75 ;
  assign n77 = n58 & ~n76 ;
  assign n78 = n77 ^ x10 ;
  assign n79 = n78 ^ x7 ;
  assign n80 = x5 ^ x4 ;
  assign n81 = n80 ^ x3 ;
  assign n82 = n81 ^ x4 ;
  assign n83 = x8 ^ x4 ;
  assign n84 = n83 ^ x4 ;
  assign n85 = n82 & ~n84 ;
  assign n86 = n85 ^ x4 ;
  assign n87 = ~x9 & n86 ;
  assign n88 = n87 ^ x5 ;
  assign n89 = ~x6 & ~n88 ;
  assign n90 = n89 ^ n49 ;
  assign n91 = x10 & n90 ;
  assign n92 = n91 ^ n89 ;
  assign n93 = ~n79 & ~n92 ;
  assign n94 = n93 ^ n91 ;
  assign n95 = n94 ^ n89 ;
  assign n96 = n95 ^ x10 ;
  assign n97 = x7 & ~n96 ;
  assign n98 = ~n68 & ~n97 ;
  assign y0 = ~n98 ;
endmodule
