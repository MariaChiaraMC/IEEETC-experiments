module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 ;
  assign n9 = ~x0 & ~x2 ;
  assign n10 = x1 & n9 ;
  assign n11 = x5 ^ x4 ;
  assign n12 = n11 ^ x3 ;
  assign n13 = x7 ^ x6 ;
  assign n14 = x6 & n13 ;
  assign n15 = n14 ^ x4 ;
  assign n16 = n15 ^ x6 ;
  assign n17 = n12 & n16 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = n18 ^ x6 ;
  assign n20 = x3 & n19 ;
  assign n21 = n20 ^ x3 ;
  assign n22 = n10 & ~n21 ;
  assign y0 = ~n22 ;
endmodule
