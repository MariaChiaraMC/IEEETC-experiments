module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 ;
  assign n11 = x2 & ~x6 ;
  assign n12 = ~x5 & x7 ;
  assign n13 = ~x1 & x4 ;
  assign n14 = ~x3 & x8 ;
  assign n15 = n13 & n14 ;
  assign n16 = n12 & n15 ;
  assign n17 = n11 & n16 ;
  assign n18 = x5 & x6 ;
  assign n19 = x3 & x4 ;
  assign n20 = n18 & n19 ;
  assign n21 = x2 & ~x7 ;
  assign n22 = ~x1 & ~x8 ;
  assign n23 = n21 & n22 ;
  assign n24 = n20 & n23 ;
  assign n25 = n24 ^ n17 ;
  assign n26 = ~x2 & x7 ;
  assign n30 = ~x6 & ~x8 ;
  assign n27 = ~x1 & x6 ;
  assign n28 = ~n14 & ~n19 ;
  assign n29 = n27 & ~n28 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = ~x3 & x4 ;
  assign n34 = x1 & n33 ;
  assign n35 = n34 ^ n29 ;
  assign n36 = n35 ^ n29 ;
  assign n37 = n32 & n36 ;
  assign n38 = n37 ^ n29 ;
  assign n39 = x5 & n38 ;
  assign n40 = n39 ^ n29 ;
  assign n41 = n26 & n40 ;
  assign n42 = ~x1 & ~x3 ;
  assign n43 = ~x5 & ~x8 ;
  assign n44 = n11 & n43 ;
  assign n45 = n42 & n44 ;
  assign n46 = x4 & n45 ;
  assign n67 = ~x3 & ~x5 ;
  assign n68 = x3 & x5 ;
  assign n69 = ~n67 & ~n68 ;
  assign n47 = x1 & ~x2 ;
  assign n48 = ~x3 & ~x6 ;
  assign n49 = x5 & x8 ;
  assign n50 = n48 & n49 ;
  assign n51 = x3 & ~x6 ;
  assign n52 = ~x3 & x6 ;
  assign n53 = ~n51 & ~n52 ;
  assign n54 = x6 & ~x8 ;
  assign n55 = x1 & ~x5 ;
  assign n56 = ~n54 & n55 ;
  assign n57 = ~n53 & n56 ;
  assign n58 = ~n50 & ~n57 ;
  assign n59 = ~n47 & ~n58 ;
  assign n60 = x1 & x5 ;
  assign n61 = ~x2 & x3 ;
  assign n62 = n54 & n61 ;
  assign n63 = ~n60 & n62 ;
  assign n64 = ~n59 & ~n63 ;
  assign n70 = n69 ^ n64 ;
  assign n71 = n70 ^ n64 ;
  assign n65 = n64 ^ n47 ;
  assign n66 = n65 ^ n64 ;
  assign n72 = n71 ^ n66 ;
  assign n73 = n52 ^ x6 ;
  assign n74 = ~x8 & ~n73 ;
  assign n75 = n74 ^ x6 ;
  assign n76 = n75 ^ n64 ;
  assign n77 = n76 ^ n64 ;
  assign n78 = n77 ^ n71 ;
  assign n79 = n71 & ~n78 ;
  assign n80 = n79 ^ n71 ;
  assign n81 = n72 & n80 ;
  assign n82 = n81 ^ n79 ;
  assign n83 = n82 ^ n64 ;
  assign n84 = n83 ^ n71 ;
  assign n85 = x4 & ~n84 ;
  assign n86 = n85 ^ n64 ;
  assign n87 = n86 ^ x7 ;
  assign n88 = n87 ^ n86 ;
  assign n89 = n88 ^ n46 ;
  assign n90 = ~x4 & ~x5 ;
  assign n91 = n22 & n90 ;
  assign n92 = ~x4 & ~x8 ;
  assign n93 = x1 & x3 ;
  assign n94 = x5 ^ x4 ;
  assign n95 = n93 & n94 ;
  assign n96 = ~n92 & n95 ;
  assign n97 = ~n91 & ~n96 ;
  assign n98 = n97 ^ n11 ;
  assign n99 = ~n97 & ~n98 ;
  assign n100 = n99 ^ n86 ;
  assign n101 = n100 ^ n97 ;
  assign n102 = ~n89 & n101 ;
  assign n103 = n102 ^ n99 ;
  assign n104 = n103 ^ n97 ;
  assign n105 = ~n46 & ~n104 ;
  assign n106 = n105 ^ n46 ;
  assign n107 = ~n41 & ~n106 ;
  assign n108 = n107 ^ x0 ;
  assign n109 = n108 ^ n107 ;
  assign n110 = ~x5 & ~x7 ;
  assign n111 = n53 & n110 ;
  assign n112 = ~x1 & n111 ;
  assign n113 = x6 ^ x1 ;
  assign n114 = n69 ^ x1 ;
  assign n115 = n113 & ~n114 ;
  assign n116 = x7 & n115 ;
  assign n117 = ~n112 & ~n116 ;
  assign n118 = ~x4 & ~n117 ;
  assign n119 = x7 ^ x5 ;
  assign n120 = n119 ^ x3 ;
  assign n121 = n120 ^ n13 ;
  assign n122 = x6 ^ x3 ;
  assign n123 = n122 ^ x3 ;
  assign n124 = x7 ^ x3 ;
  assign n125 = n124 ^ x3 ;
  assign n126 = ~n123 & n125 ;
  assign n127 = n126 ^ x3 ;
  assign n128 = n127 ^ n120 ;
  assign n129 = ~n121 & ~n128 ;
  assign n130 = n129 ^ n126 ;
  assign n131 = n130 ^ x3 ;
  assign n132 = n131 ^ n13 ;
  assign n133 = ~n120 & n132 ;
  assign n134 = n133 ^ n120 ;
  assign n135 = ~n118 & n134 ;
  assign n136 = x2 & ~n135 ;
  assign n137 = x6 & x7 ;
  assign n138 = x4 & ~n137 ;
  assign n139 = x1 & ~x6 ;
  assign n140 = ~x2 & ~x3 ;
  assign n141 = ~n139 & n140 ;
  assign n142 = x1 & ~x7 ;
  assign n143 = n142 ^ n13 ;
  assign n144 = n143 ^ n13 ;
  assign n145 = n13 ^ x6 ;
  assign n146 = n145 ^ n13 ;
  assign n147 = ~n144 & n146 ;
  assign n148 = n147 ^ n13 ;
  assign n149 = x5 & ~n148 ;
  assign n150 = n149 ^ n13 ;
  assign n151 = n141 & n150 ;
  assign n152 = ~n138 & n151 ;
  assign n153 = ~n136 & ~n152 ;
  assign n154 = ~x8 & ~n153 ;
  assign n155 = x2 & ~n49 ;
  assign n156 = ~x1 & ~n155 ;
  assign n157 = x7 & ~n94 ;
  assign n158 = n156 & n157 ;
  assign n159 = ~x2 & ~x7 ;
  assign n160 = x8 & n159 ;
  assign n161 = n90 & n160 ;
  assign n162 = ~n158 & ~n161 ;
  assign n163 = x6 & ~n162 ;
  assign n164 = x3 & n163 ;
  assign n165 = n33 & n159 ;
  assign n166 = x6 & x8 ;
  assign n167 = ~n60 & n166 ;
  assign n168 = n165 & n167 ;
  assign n169 = x5 & ~x7 ;
  assign n170 = n11 & n169 ;
  assign n171 = n170 ^ x7 ;
  assign n172 = n171 ^ n170 ;
  assign n173 = ~x5 & n166 ;
  assign n174 = n173 ^ n170 ;
  assign n175 = n174 ^ n170 ;
  assign n176 = n172 & n175 ;
  assign n177 = n176 ^ n170 ;
  assign n178 = x4 & n177 ;
  assign n179 = n178 ^ n170 ;
  assign n180 = n93 & n179 ;
  assign n181 = ~n168 & ~n180 ;
  assign n182 = ~n164 & n181 ;
  assign n183 = ~n154 & n182 ;
  assign n184 = n183 ^ n107 ;
  assign n185 = n109 & n184 ;
  assign n186 = n185 ^ n107 ;
  assign n187 = n186 ^ n17 ;
  assign n188 = n25 & ~n187 ;
  assign n189 = n188 ^ n185 ;
  assign n190 = n189 ^ n107 ;
  assign n191 = n190 ^ n24 ;
  assign n192 = ~n17 & ~n191 ;
  assign n193 = n192 ^ n17 ;
  assign n194 = ~x9 & n193 ;
  assign n195 = x3 & x9 ;
  assign n196 = x1 ^ x0 ;
  assign n197 = n26 ^ n21 ;
  assign n198 = n21 ^ x1 ;
  assign n199 = n198 ^ n21 ;
  assign n200 = n197 & n199 ;
  assign n201 = n200 ^ n21 ;
  assign n202 = n196 & n201 ;
  assign n203 = n195 & n202 ;
  assign n204 = n173 & n203 ;
  assign n217 = x5 & n197 ;
  assign n218 = n217 ^ n21 ;
  assign n219 = n22 & n218 ;
  assign n220 = n47 & n110 ;
  assign n221 = x8 & n220 ;
  assign n222 = ~n219 & ~n221 ;
  assign n205 = n11 & n49 ;
  assign n206 = n205 ^ n54 ;
  assign n207 = n206 ^ n205 ;
  assign n208 = x5 ^ x2 ;
  assign n209 = ~n119 & ~n208 ;
  assign n210 = n209 ^ x2 ;
  assign n211 = n210 ^ n205 ;
  assign n212 = n211 ^ n205 ;
  assign n213 = n207 & n212 ;
  assign n214 = n213 ^ n205 ;
  assign n215 = x1 & n214 ;
  assign n216 = n215 ^ n205 ;
  assign n223 = n222 ^ n216 ;
  assign n224 = n223 ^ n216 ;
  assign n225 = n216 ^ x6 ;
  assign n226 = n225 ^ n216 ;
  assign n227 = ~n224 & ~n226 ;
  assign n228 = n227 ^ n216 ;
  assign n229 = x3 & n228 ;
  assign n230 = n229 ^ n216 ;
  assign n231 = x0 & n230 ;
  assign n232 = x2 & x5 ;
  assign n233 = x7 & ~n49 ;
  assign n234 = ~n232 & n233 ;
  assign n235 = ~n166 & ~n234 ;
  assign n236 = x2 & ~x3 ;
  assign n237 = ~n21 & ~n236 ;
  assign n238 = ~n18 & n237 ;
  assign n239 = n47 & ~n67 ;
  assign n240 = ~x0 & ~n239 ;
  assign n241 = n238 & n240 ;
  assign n242 = n69 ^ x8 ;
  assign n243 = n242 ^ n69 ;
  assign n244 = n69 ^ n61 ;
  assign n245 = ~n243 & n244 ;
  assign n246 = n245 ^ n69 ;
  assign n247 = ~x1 & ~n246 ;
  assign n248 = n247 ^ x8 ;
  assign n249 = n241 & n248 ;
  assign n250 = n235 & n249 ;
  assign n251 = x0 & x3 ;
  assign n252 = n166 & n251 ;
  assign n253 = n232 & n252 ;
  assign n254 = n253 ^ x1 ;
  assign n255 = n254 ^ n253 ;
  assign n256 = ~x2 & x6 ;
  assign n257 = x3 & n256 ;
  assign n258 = n49 & n257 ;
  assign n259 = n258 ^ n253 ;
  assign n260 = n259 ^ n253 ;
  assign n261 = n255 & n260 ;
  assign n262 = n261 ^ n253 ;
  assign n263 = ~x7 & n262 ;
  assign n264 = n263 ^ n253 ;
  assign n265 = ~n250 & ~n264 ;
  assign n266 = ~n231 & n265 ;
  assign n267 = x9 & ~n266 ;
  assign n268 = x0 & ~x1 ;
  assign n269 = n140 & n268 ;
  assign n270 = ~x0 & x2 ;
  assign n271 = n93 & n270 ;
  assign n272 = ~n269 & ~n271 ;
  assign n273 = n173 & ~n272 ;
  assign n274 = ~x7 & n273 ;
  assign n275 = ~n267 & ~n274 ;
  assign n276 = n275 ^ x4 ;
  assign n277 = n276 ^ n275 ;
  assign n278 = n68 & n270 ;
  assign n279 = ~x7 & x9 ;
  assign n280 = n278 & n279 ;
  assign n281 = n54 & n280 ;
  assign n322 = x6 ^ x2 ;
  assign n339 = n48 ^ x0 ;
  assign n340 = ~n322 & ~n339 ;
  assign n341 = n169 & n340 ;
  assign n342 = n11 & n67 ;
  assign n343 = ~n257 & ~n342 ;
  assign n344 = x0 & ~n343 ;
  assign n345 = n344 ^ x7 ;
  assign n346 = n345 ^ n344 ;
  assign n347 = n344 ^ n278 ;
  assign n348 = n346 & n347 ;
  assign n349 = n348 ^ n344 ;
  assign n350 = ~n341 & ~n349 ;
  assign n351 = ~x8 & ~n350 ;
  assign n352 = ~n14 & ~n256 ;
  assign n353 = n12 & ~n140 ;
  assign n354 = ~n352 & n353 ;
  assign n355 = ~x0 & n354 ;
  assign n356 = ~n351 & ~n355 ;
  assign n357 = x9 & ~n356 ;
  assign n287 = x8 & n52 ;
  assign n288 = x3 & ~n18 ;
  assign n289 = ~n287 & ~n288 ;
  assign n282 = ~x0 & n48 ;
  assign n283 = n43 & n282 ;
  assign n284 = ~n252 & ~n283 ;
  assign n290 = n289 ^ n284 ;
  assign n291 = n290 ^ n284 ;
  assign n285 = n284 ^ x0 ;
  assign n286 = n285 ^ n284 ;
  assign n292 = n291 ^ n286 ;
  assign n293 = ~n43 & ~n49 ;
  assign n294 = n293 ^ n284 ;
  assign n295 = n294 ^ n284 ;
  assign n296 = n295 ^ n291 ;
  assign n297 = ~n291 & n296 ;
  assign n298 = n297 ^ n291 ;
  assign n299 = n292 & ~n298 ;
  assign n300 = n299 ^ n297 ;
  assign n301 = n300 ^ n284 ;
  assign n302 = n301 ^ n291 ;
  assign n303 = ~x2 & n302 ;
  assign n304 = n303 ^ n284 ;
  assign n305 = n279 & ~n304 ;
  assign n306 = n232 & n287 ;
  assign n307 = n173 ^ n61 ;
  assign n308 = n307 ^ n173 ;
  assign n309 = n308 ^ x0 ;
  assign n310 = x5 & n30 ;
  assign n311 = x2 & ~n195 ;
  assign n312 = n311 ^ n310 ;
  assign n313 = n310 & ~n312 ;
  assign n314 = n313 ^ n173 ;
  assign n315 = n314 ^ n310 ;
  assign n316 = ~n309 & n315 ;
  assign n317 = n316 ^ n313 ;
  assign n318 = n317 ^ n310 ;
  assign n319 = x0 & n318 ;
  assign n320 = n319 ^ x0 ;
  assign n321 = ~n306 & n320 ;
  assign n323 = n322 ^ x6 ;
  assign n327 = ~x6 & x8 ;
  assign n328 = ~x5 & n327 ;
  assign n329 = n328 ^ n293 ;
  assign n324 = n323 ^ x6 ;
  assign n325 = n323 ^ n293 ;
  assign n326 = n324 & n325 ;
  assign n330 = n329 ^ n326 ;
  assign n331 = n323 & n330 ;
  assign n332 = n331 ^ n328 ;
  assign n333 = n332 ^ n323 ;
  assign n334 = n195 & n333 ;
  assign n335 = ~x0 & ~n334 ;
  assign n336 = x7 & ~n335 ;
  assign n337 = ~n321 & n336 ;
  assign n338 = ~n305 & ~n337 ;
  assign n358 = n357 ^ n338 ;
  assign n359 = n358 ^ x1 ;
  assign n366 = n359 ^ n358 ;
  assign n360 = n359 ^ n47 ;
  assign n361 = n360 ^ n358 ;
  assign n362 = n359 ^ n338 ;
  assign n363 = n362 ^ n47 ;
  assign n364 = n363 ^ n361 ;
  assign n365 = n361 & n364 ;
  assign n367 = n366 ^ n365 ;
  assign n368 = n367 ^ n361 ;
  assign n369 = x3 ^ x0 ;
  assign n370 = n169 ^ x3 ;
  assign n371 = n370 ^ n169 ;
  assign n372 = n169 ^ n12 ;
  assign n373 = ~n371 & n372 ;
  assign n374 = n373 ^ n169 ;
  assign n375 = ~n369 & n374 ;
  assign n376 = n327 & n375 ;
  assign n377 = n376 ^ n358 ;
  assign n378 = n365 ^ n361 ;
  assign n379 = ~n377 & n378 ;
  assign n380 = n379 ^ n358 ;
  assign n381 = ~n368 & ~n380 ;
  assign n382 = n381 ^ n358 ;
  assign n383 = n382 ^ n357 ;
  assign n384 = n383 ^ n358 ;
  assign n385 = ~n281 & ~n384 ;
  assign n386 = n385 ^ n275 ;
  assign n387 = ~n277 & n386 ;
  assign n388 = n387 ^ n275 ;
  assign n389 = ~n204 & n388 ;
  assign n390 = ~n194 & n389 ;
  assign y0 = ~n390 ;
endmodule
