module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 ;
  assign n15 = ~x5 & x6 ;
  assign n16 = x0 & ~x11 ;
  assign n17 = x9 & ~x13 ;
  assign n18 = n16 & n17 ;
  assign n25 = n18 ^ x10 ;
  assign n36 = n25 ^ n18 ;
  assign n19 = ~x0 & x10 ;
  assign n20 = ~x11 & ~x12 ;
  assign n21 = ~x13 & n20 ;
  assign n22 = ~n19 & n21 ;
  assign n23 = ~x9 & ~n22 ;
  assign n24 = n23 ^ n18 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = n27 ^ n18 ;
  assign n29 = ~x0 & x12 ;
  assign n30 = x13 & n29 ;
  assign n31 = x11 & n30 ;
  assign n32 = n31 ^ n26 ;
  assign n33 = n32 ^ n26 ;
  assign n34 = n33 ^ n28 ;
  assign n35 = n28 & ~n34 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = n37 ^ n28 ;
  assign n39 = n20 ^ n18 ;
  assign n40 = n35 ^ n28 ;
  assign n41 = ~n39 & n40 ;
  assign n42 = n41 ^ n18 ;
  assign n43 = ~n38 & ~n42 ;
  assign n44 = n43 ^ n18 ;
  assign n45 = n44 ^ x10 ;
  assign n46 = n45 ^ n18 ;
  assign n47 = n15 & ~n46 ;
  assign y0 = n47 ;
endmodule
