module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 ;
  assign n16 = x3 & x4 ;
  assign n17 = x1 & n16 ;
  assign n18 = x9 & x13 ;
  assign n19 = ~x8 & n18 ;
  assign n20 = x5 & x7 ;
  assign n21 = x2 & ~n20 ;
  assign n22 = n19 & n21 ;
  assign n23 = x10 ^ x7 ;
  assign n24 = x6 & n23 ;
  assign n25 = n22 & ~n24 ;
  assign n26 = n25 ^ x0 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = ~x5 & x14 ;
  assign n29 = x6 & x7 ;
  assign n30 = ~x2 & n29 ;
  assign n31 = n28 & n30 ;
  assign n32 = n31 ^ n25 ;
  assign n33 = n27 & n32 ;
  assign n34 = n33 ^ n25 ;
  assign n35 = n17 & n34 ;
  assign n36 = x2 & x7 ;
  assign n37 = x10 & n36 ;
  assign n38 = ~x4 & ~x6 ;
  assign n39 = ~x0 & ~x1 ;
  assign n40 = n38 & n39 ;
  assign n41 = n37 & n40 ;
  assign n42 = x3 & n41 ;
  assign n54 = ~x2 & ~x10 ;
  assign n55 = n17 & n29 ;
  assign n56 = n54 & n55 ;
  assign n43 = ~x7 & ~x10 ;
  assign n44 = ~x3 & ~x4 ;
  assign n45 = n43 & n44 ;
  assign n46 = n45 ^ x6 ;
  assign n47 = n46 ^ n45 ;
  assign n48 = x7 & x10 ;
  assign n49 = n16 & n48 ;
  assign n50 = n49 ^ n45 ;
  assign n51 = n47 & n50 ;
  assign n52 = n51 ^ n45 ;
  assign n53 = n39 & n52 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n56 ^ x2 ;
  assign n59 = n56 ^ x9 ;
  assign n60 = ~n56 & n59 ;
  assign n61 = n60 ^ n56 ;
  assign n62 = ~n58 & ~n61 ;
  assign n63 = n62 ^ n60 ;
  assign n64 = n63 ^ n56 ;
  assign n65 = n64 ^ x9 ;
  assign n66 = n57 & n65 ;
  assign n67 = n66 ^ n56 ;
  assign n68 = ~n42 & ~n67 ;
  assign n69 = ~x5 & ~x8 ;
  assign n70 = ~n68 & n69 ;
  assign n71 = n70 ^ x14 ;
  assign n72 = n71 ^ n70 ;
  assign n73 = n72 ^ x13 ;
  assign n74 = ~x2 & ~x8 ;
  assign n75 = ~x1 & ~n74 ;
  assign n76 = x0 & x6 ;
  assign n77 = n44 & n76 ;
  assign n78 = ~x8 & x9 ;
  assign n79 = ~x10 & ~n78 ;
  assign n80 = n77 & n79 ;
  assign n81 = x9 ^ x7 ;
  assign n82 = x5 ^ x2 ;
  assign n83 = x9 ^ x5 ;
  assign n84 = n83 ^ x5 ;
  assign n85 = ~n82 & n84 ;
  assign n86 = n85 ^ x5 ;
  assign n87 = ~n81 & ~n86 ;
  assign n88 = n87 ^ x5 ;
  assign n89 = n80 & ~n88 ;
  assign n90 = ~n75 & n89 ;
  assign n99 = ~x7 & x9 ;
  assign n91 = x8 & ~x10 ;
  assign n92 = x2 & x4 ;
  assign n93 = ~n91 & ~n92 ;
  assign n94 = x7 & ~x9 ;
  assign n95 = x4 & x8 ;
  assign n96 = n94 & ~n95 ;
  assign n97 = n76 & n96 ;
  assign n98 = ~n93 & n97 ;
  assign n100 = n99 ^ n98 ;
  assign n101 = n100 ^ x5 ;
  assign n111 = n101 ^ n100 ;
  assign n102 = ~x4 & n76 ;
  assign n103 = ~x5 & n102 ;
  assign n104 = n91 & n103 ;
  assign n105 = n104 ^ n101 ;
  assign n106 = n105 ^ n100 ;
  assign n107 = n101 ^ n98 ;
  assign n108 = n107 ^ n104 ;
  assign n109 = n108 ^ n106 ;
  assign n110 = n106 & ~n109 ;
  assign n112 = n111 ^ n110 ;
  assign n113 = n112 ^ n106 ;
  assign n114 = ~x0 & ~x8 ;
  assign n115 = x4 ^ x2 ;
  assign n116 = x6 ^ x4 ;
  assign n117 = x10 ^ x6 ;
  assign n118 = ~n116 & ~n117 ;
  assign n119 = ~n115 & n118 ;
  assign n120 = n114 & n119 ;
  assign n121 = n120 ^ n100 ;
  assign n122 = n110 ^ n106 ;
  assign n123 = ~n121 & n122 ;
  assign n124 = n123 ^ n100 ;
  assign n125 = ~n113 & n124 ;
  assign n126 = n125 ^ n100 ;
  assign n127 = n126 ^ n99 ;
  assign n128 = n127 ^ n100 ;
  assign n129 = ~x1 & n128 ;
  assign n130 = x2 & ~x10 ;
  assign n131 = n103 & n130 ;
  assign n132 = n78 & n81 ;
  assign n133 = n132 ^ n81 ;
  assign n134 = n131 & n133 ;
  assign n135 = ~n129 & ~n134 ;
  assign n136 = x3 & ~n135 ;
  assign n137 = n136 ^ n90 ;
  assign n138 = ~n90 & n137 ;
  assign n139 = n138 ^ n70 ;
  assign n140 = n139 ^ n90 ;
  assign n141 = n73 & n140 ;
  assign n142 = n141 ^ n138 ;
  assign n143 = n142 ^ n90 ;
  assign n144 = ~x13 & ~n143 ;
  assign n145 = n144 ^ x13 ;
  assign n146 = ~n35 & n145 ;
  assign n147 = ~x11 & ~n146 ;
  assign n148 = ~x12 & n147 ;
  assign y0 = n148 ;
endmodule
