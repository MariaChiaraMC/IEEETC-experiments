module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 ;
  output y0 ;
  wire n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 ;
  assign n23 = x3 & ~x5 ;
  assign n24 = ~x4 & ~n23 ;
  assign n25 = x1 ^ x0 ;
  assign n26 = x3 ^ x2 ;
  assign n27 = x2 ^ x1 ;
  assign n28 = n27 ^ x2 ;
  assign n29 = ~n26 & ~n28 ;
  assign n30 = n29 ^ x2 ;
  assign n31 = n25 & ~n30 ;
  assign n32 = n24 & n31 ;
  assign n33 = x14 & ~n32 ;
  assign n205 = ~x19 & ~x20 ;
  assign n34 = ~x12 & ~x13 ;
  assign n35 = ~x6 & ~x7 ;
  assign n36 = ~x8 & n35 ;
  assign n37 = x10 & ~x11 ;
  assign n38 = n36 & n37 ;
  assign n39 = ~x0 & x1 ;
  assign n40 = ~x3 & ~x4 ;
  assign n41 = n39 & n40 ;
  assign n42 = n38 & n41 ;
  assign n43 = ~x2 & x3 ;
  assign n44 = x0 & ~x1 ;
  assign n45 = ~x11 & n36 ;
  assign n46 = n44 & n45 ;
  assign n47 = x11 & n35 ;
  assign n48 = ~x10 & n47 ;
  assign n49 = ~x1 & n37 ;
  assign n50 = ~n48 & ~n49 ;
  assign n51 = ~x0 & ~x4 ;
  assign n52 = ~n50 & n51 ;
  assign n53 = x8 & n52 ;
  assign n54 = ~n46 & ~n53 ;
  assign n55 = n43 & ~n54 ;
  assign n56 = x8 & n37 ;
  assign n57 = n41 & n56 ;
  assign n58 = x0 & x2 ;
  assign n59 = ~x5 & n58 ;
  assign n60 = n40 & n59 ;
  assign n61 = x8 & n48 ;
  assign n62 = ~x1 & ~x10 ;
  assign n63 = n45 & ~n62 ;
  assign n64 = ~n61 & ~n63 ;
  assign n65 = n60 & ~n64 ;
  assign n66 = ~n57 & ~n65 ;
  assign n67 = ~n55 & n66 ;
  assign n68 = x9 & ~n67 ;
  assign n69 = ~n42 & ~n68 ;
  assign n70 = n34 & ~n69 ;
  assign n71 = ~x3 & x4 ;
  assign n72 = x10 & x11 ;
  assign n73 = x9 & ~x12 ;
  assign n74 = n72 & n73 ;
  assign n75 = ~x13 & ~n74 ;
  assign n76 = x0 & ~n75 ;
  assign n77 = ~x15 & n76 ;
  assign n78 = ~n58 & ~n77 ;
  assign n79 = n71 & ~n78 ;
  assign n80 = ~x3 & ~x21 ;
  assign n81 = x2 & ~n80 ;
  assign n82 = ~x0 & ~n81 ;
  assign n83 = ~x1 & ~x2 ;
  assign n84 = ~x16 & n83 ;
  assign n85 = ~n39 & ~n84 ;
  assign n86 = x3 & n34 ;
  assign n87 = n38 ^ x2 ;
  assign n88 = n87 ^ x9 ;
  assign n97 = n88 ^ n87 ;
  assign n89 = ~x8 & ~x9 ;
  assign n90 = n48 & n89 ;
  assign n91 = n90 ^ n88 ;
  assign n92 = n91 ^ n87 ;
  assign n93 = n88 ^ n38 ;
  assign n94 = n93 ^ n90 ;
  assign n95 = n94 ^ n92 ;
  assign n96 = n92 & ~n95 ;
  assign n98 = n97 ^ n96 ;
  assign n99 = n98 ^ n92 ;
  assign n100 = ~n45 & ~n61 ;
  assign n101 = ~n56 & n100 ;
  assign n102 = n101 ^ n87 ;
  assign n103 = n96 ^ n92 ;
  assign n104 = n102 & n103 ;
  assign n105 = n104 ^ n87 ;
  assign n106 = ~n99 & n105 ;
  assign n107 = n106 ^ n87 ;
  assign n108 = n107 ^ x2 ;
  assign n109 = n108 ^ n87 ;
  assign n110 = n86 & n109 ;
  assign n111 = n85 & ~n110 ;
  assign n112 = ~n82 & n111 ;
  assign n113 = ~x4 & ~n112 ;
  assign n114 = ~x9 & ~x10 ;
  assign n115 = ~n73 & ~n114 ;
  assign n116 = ~x10 & ~x11 ;
  assign n117 = ~x8 & ~n116 ;
  assign n118 = ~n115 & n117 ;
  assign n119 = ~x15 & ~n118 ;
  assign n120 = ~x6 & ~n119 ;
  assign n121 = x13 & ~n120 ;
  assign n122 = ~x9 & n35 ;
  assign n123 = x10 & ~x13 ;
  assign n124 = x16 & n123 ;
  assign n125 = n122 & n124 ;
  assign n126 = x7 & x16 ;
  assign n127 = ~x8 & x13 ;
  assign n128 = n114 & n127 ;
  assign n129 = n126 & n128 ;
  assign n130 = ~n125 & ~n129 ;
  assign n131 = x11 & ~n130 ;
  assign n132 = ~x13 & ~n36 ;
  assign n133 = x11 & ~x16 ;
  assign n134 = ~n123 & ~n133 ;
  assign n135 = ~n132 & ~n134 ;
  assign n136 = ~x15 & n135 ;
  assign n137 = ~n131 & ~n136 ;
  assign n138 = ~x12 & ~n137 ;
  assign n139 = ~n121 & ~n138 ;
  assign n140 = n56 ^ x11 ;
  assign n141 = x7 & n140 ;
  assign n142 = x6 & n141 ;
  assign n143 = x11 & ~x15 ;
  assign n144 = n143 ^ x8 ;
  assign n145 = n143 ^ x10 ;
  assign n146 = n145 ^ x10 ;
  assign n147 = n146 ^ n144 ;
  assign n148 = n35 & n116 ;
  assign n149 = n148 ^ n144 ;
  assign n150 = ~x13 & n149 ;
  assign n151 = n150 ^ x10 ;
  assign n152 = n147 & ~n151 ;
  assign n153 = n152 ^ n150 ;
  assign n154 = n144 & n153 ;
  assign n155 = n154 ^ n150 ;
  assign n156 = n155 ^ n152 ;
  assign n157 = n156 ^ n143 ;
  assign n158 = ~n142 & ~n157 ;
  assign n159 = n73 & ~n158 ;
  assign n160 = ~x16 & n122 ;
  assign n161 = n56 & n160 ;
  assign n162 = n72 & n89 ;
  assign n163 = ~x16 & n162 ;
  assign n164 = ~x12 & ~n163 ;
  assign n165 = x16 ^ x7 ;
  assign n166 = ~x6 & ~n165 ;
  assign n167 = ~n164 & n166 ;
  assign n168 = ~n161 & ~n167 ;
  assign n169 = ~x13 & ~n168 ;
  assign n170 = ~x17 & ~n169 ;
  assign n171 = ~n159 & n170 ;
  assign n172 = n139 & n171 ;
  assign n173 = n71 & ~n172 ;
  assign n174 = n173 ^ x3 ;
  assign n175 = n174 ^ n173 ;
  assign n176 = ~x0 & x15 ;
  assign n177 = n176 ^ n173 ;
  assign n178 = n177 ^ n173 ;
  assign n179 = n175 & ~n178 ;
  assign n180 = n179 ^ n173 ;
  assign n181 = ~x2 & n180 ;
  assign n182 = n181 ^ n173 ;
  assign n183 = n182 ^ x1 ;
  assign n184 = n183 ^ n182 ;
  assign n185 = x3 & n58 ;
  assign n186 = n185 ^ n182 ;
  assign n187 = n184 & n186 ;
  assign n188 = n187 ^ n182 ;
  assign n189 = ~n113 & ~n188 ;
  assign n190 = ~n79 & n189 ;
  assign n191 = x5 & ~n190 ;
  assign n192 = n23 ^ x1 ;
  assign n193 = n192 ^ n23 ;
  assign n194 = x5 & x15 ;
  assign n195 = n194 ^ n23 ;
  assign n196 = n195 ^ n23 ;
  assign n197 = ~n193 & ~n196 ;
  assign n198 = n197 ^ n23 ;
  assign n199 = ~x2 & n198 ;
  assign n200 = n199 ^ n23 ;
  assign n201 = x4 & n200 ;
  assign n202 = x0 & n201 ;
  assign n203 = ~n191 & ~n202 ;
  assign n204 = ~n70 & n203 ;
  assign n206 = n205 ^ n204 ;
  assign n207 = n206 ^ n204 ;
  assign n208 = n204 ^ x18 ;
  assign n209 = ~n207 & n208 ;
  assign n210 = n209 ^ n204 ;
  assign n211 = n33 & n210 ;
  assign y0 = ~n211 ;
endmodule
