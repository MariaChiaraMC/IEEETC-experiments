module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 ;
  assign n7 = ~x4 & ~x5 ;
  assign n8 = ~x3 & n7 ;
  assign n9 = x3 & ~n7 ;
  assign n10 = ~x2 & ~x4 ;
  assign n11 = x1 & ~n10 ;
  assign n12 = ~n9 & n11 ;
  assign n13 = ~n8 & n12 ;
  assign n14 = x1 & x3 ;
  assign n15 = n14 ^ x0 ;
  assign n16 = n15 ^ x0 ;
  assign n17 = x2 ^ x0 ;
  assign n18 = x4 ^ x3 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = x4 ^ x2 ;
  assign n22 = n21 ^ x5 ;
  assign n23 = x5 & ~n22 ;
  assign n24 = n23 ^ x2 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = ~n20 & ~n25 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = n27 ^ x5 ;
  assign n29 = ~n17 & n28 ;
  assign n30 = n29 ^ x2 ;
  assign n31 = n30 ^ x0 ;
  assign n32 = ~n16 & n31 ;
  assign n33 = n32 ^ x0 ;
  assign n34 = x2 & ~x3 ;
  assign n35 = ~x0 & n34 ;
  assign n36 = n35 ^ n13 ;
  assign n37 = ~n33 & ~n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = ~n13 & n38 ;
  assign n40 = n39 ^ n13 ;
  assign y0 = n40 ;
endmodule
