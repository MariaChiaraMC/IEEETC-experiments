module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 ;
  assign n24 = ~x6 & ~x7 ;
  assign n43 = ~x1 & n24 ;
  assign n44 = ~x4 & x5 ;
  assign n45 = ~x7 & n44 ;
  assign n46 = ~n43 & ~n45 ;
  assign n47 = ~x3 & ~n46 ;
  assign n48 = x6 ^ x4 ;
  assign n49 = n48 ^ x5 ;
  assign n57 = n49 ^ x6 ;
  assign n50 = n49 ^ x3 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = n51 ^ x6 ;
  assign n53 = n50 ^ x5 ;
  assign n54 = n53 ^ n50 ;
  assign n55 = n54 ^ n52 ;
  assign n56 = n52 & ~n55 ;
  assign n58 = n57 ^ n56 ;
  assign n59 = n58 ^ n52 ;
  assign n60 = x7 ^ x6 ;
  assign n61 = n60 ^ x6 ;
  assign n62 = n56 ^ n52 ;
  assign n63 = n61 & n62 ;
  assign n64 = n63 ^ x6 ;
  assign n65 = n59 & n64 ;
  assign n66 = n65 ^ x6 ;
  assign n67 = n66 ^ n48 ;
  assign n68 = n67 ^ x6 ;
  assign n69 = ~n47 & ~n68 ;
  assign n9 = x4 ^ x3 ;
  assign n10 = n9 ^ x1 ;
  assign n13 = n10 ^ x5 ;
  assign n11 = n10 ^ x1 ;
  assign n12 = n11 ^ x1 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n11 ^ x3 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n14 & ~n16 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = n13 ^ n11 ;
  assign n20 = n19 ^ n15 ;
  assign n25 = n24 ^ x1 ;
  assign n26 = n15 ^ n12 ;
  assign n27 = ~n25 & n26 ;
  assign n21 = x6 ^ x1 ;
  assign n22 = n21 ^ n13 ;
  assign n23 = n19 & n22 ;
  assign n28 = n27 ^ n23 ;
  assign n29 = n28 ^ x1 ;
  assign n30 = n29 ^ n11 ;
  assign n31 = n30 ^ n15 ;
  assign n32 = ~n20 & n31 ;
  assign n33 = n32 ^ n23 ;
  assign n34 = n33 ^ n11 ;
  assign n35 = n34 ^ n15 ;
  assign n36 = ~n18 & n35 ;
  assign n37 = n36 ^ n23 ;
  assign n38 = n37 ^ n17 ;
  assign n39 = n38 ^ n32 ;
  assign n40 = n39 ^ n11 ;
  assign n41 = n40 ^ n13 ;
  assign n42 = n41 ^ n15 ;
  assign n70 = n69 ^ n42 ;
  assign n71 = n70 ^ n42 ;
  assign n72 = ~x3 & ~x5 ;
  assign n73 = ~x6 & n72 ;
  assign n74 = x1 & ~n73 ;
  assign n75 = n74 ^ n42 ;
  assign n76 = n75 ^ n42 ;
  assign n77 = n71 & ~n76 ;
  assign n78 = n77 ^ n42 ;
  assign n79 = ~x2 & ~n78 ;
  assign n80 = n79 ^ n42 ;
  assign y0 = n80 ;
endmodule
