module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 ;
  assign n12 = x5 ^ x3 ;
  assign n13 = n12 ^ x5 ;
  assign n14 = ~x5 & x7 ;
  assign n15 = n14 ^ x5 ;
  assign n16 = ~n13 & n15 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = ~x6 & n17 ;
  assign n19 = x7 ^ x5 ;
  assign n20 = x5 ^ x2 ;
  assign n21 = n20 ^ x5 ;
  assign n22 = n19 & ~n21 ;
  assign n23 = n22 ^ x5 ;
  assign n24 = ~x6 & ~n23 ;
  assign n25 = n24 ^ x2 ;
  assign n26 = ~n18 & ~n25 ;
  assign n9 = x6 & x7 ;
  assign n10 = ~x4 & ~n9 ;
  assign n11 = x3 & ~n10 ;
  assign n27 = n26 ^ n11 ;
  assign n28 = n27 ^ x4 ;
  assign n37 = n28 ^ n27 ;
  assign n29 = ~x6 & ~x7 ;
  assign n30 = ~x5 & ~n29 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = n30 ^ n11 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = n32 & n35 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = n38 ^ n32 ;
  assign n40 = n27 ^ x2 ;
  assign n41 = n36 ^ n32 ;
  assign n42 = n40 & n41 ;
  assign n43 = n42 ^ n27 ;
  assign n44 = ~n39 & ~n43 ;
  assign n45 = n44 ^ n27 ;
  assign n46 = n45 ^ n11 ;
  assign n47 = n46 ^ n27 ;
  assign n48 = ~x1 & n47 ;
  assign n49 = x7 ^ x4 ;
  assign n50 = n19 ^ x4 ;
  assign n51 = n49 & ~n50 ;
  assign n52 = ~x6 & n51 ;
  assign n53 = n52 ^ n19 ;
  assign n54 = n53 ^ x1 ;
  assign n55 = n54 ^ n53 ;
  assign n56 = n55 ^ x3 ;
  assign n57 = ~x4 & ~x5 ;
  assign n58 = n57 ^ n10 ;
  assign n59 = ~n10 & n58 ;
  assign n60 = n59 ^ n53 ;
  assign n61 = n60 ^ n10 ;
  assign n62 = ~n56 & ~n61 ;
  assign n63 = n62 ^ n59 ;
  assign n64 = n63 ^ n10 ;
  assign n65 = ~x3 & ~n64 ;
  assign n66 = n65 ^ x3 ;
  assign n67 = ~x2 & ~n66 ;
  assign n68 = ~n48 & ~n67 ;
  assign n69 = ~x0 & ~n68 ;
  assign y0 = n69 ;
endmodule
