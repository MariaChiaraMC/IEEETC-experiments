module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 ;
  assign n9 = ~x2 & ~x3 ;
  assign n10 = ~x6 & ~x7 ;
  assign n11 = x5 & ~n10 ;
  assign n12 = n11 ^ x0 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = ~x1 & ~x4 ;
  assign n15 = n14 ^ x4 ;
  assign n16 = ~n11 & n15 ;
  assign n17 = n16 ^ x4 ;
  assign n18 = n13 & ~n17 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n19 ^ x4 ;
  assign n21 = n20 ^ n11 ;
  assign n22 = n9 & n21 ;
  assign n23 = x1 ^ x0 ;
  assign n26 = x1 & x4 ;
  assign n27 = n10 & ~n26 ;
  assign n28 = ~x5 & n27 ;
  assign n29 = n28 ^ x1 ;
  assign n30 = n29 ^ x1 ;
  assign n24 = x3 ^ x1 ;
  assign n25 = n24 ^ x1 ;
  assign n31 = n30 ^ n25 ;
  assign n32 = x2 & ~n14 ;
  assign n33 = n32 ^ x1 ;
  assign n34 = n33 ^ x1 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = ~n30 & ~n35 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = ~n31 & ~n37 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n39 ^ x1 ;
  assign n41 = n40 ^ n30 ;
  assign n42 = ~n23 & n41 ;
  assign n43 = n42 ^ x0 ;
  assign n44 = ~n22 & n43 ;
  assign y0 = n44 ;
endmodule
