module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n9 = x6 & ~x7 ;
  assign n10 = ~x3 & ~n9 ;
  assign n11 = ~x4 & ~x5 ;
  assign n12 = ~x2 & n11 ;
  assign n13 = x6 ^ x3 ;
  assign n14 = x0 & n13 ;
  assign n15 = n14 ^ x3 ;
  assign n16 = n12 & ~n15 ;
  assign n17 = ~n10 & n16 ;
  assign n18 = ~x0 & x3 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = n18 ^ x0 ;
  assign n22 = ~n20 & n21 ;
  assign n23 = n22 ^ n18 ;
  assign n24 = ~x5 & ~n18 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = ~n23 & n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = x4 & n27 ;
  assign n29 = n28 ^ x4 ;
  assign n30 = ~n17 & ~n29 ;
  assign n31 = ~x1 & ~n30 ;
  assign y0 = ~n31 ;
endmodule
