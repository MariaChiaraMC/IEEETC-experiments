module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 ;
  assign n9 = ~x0 & ~x6 ;
  assign n10 = x4 & x7 ;
  assign n11 = ~x1 & n10 ;
  assign n12 = x3 & ~x5 ;
  assign n13 = n11 & n12 ;
  assign n14 = n9 & n13 ;
  assign n15 = x4 & ~x5 ;
  assign n16 = x6 & ~x7 ;
  assign n17 = ~x0 & x1 ;
  assign n18 = n16 & n17 ;
  assign n19 = n15 & n18 ;
  assign n26 = ~x6 & x7 ;
  assign n27 = ~x1 & x5 ;
  assign n28 = x7 & ~n27 ;
  assign n29 = ~n26 & ~n28 ;
  assign n30 = ~x4 & x6 ;
  assign n31 = x5 ^ x1 ;
  assign n32 = n31 ^ x5 ;
  assign n33 = n15 ^ x5 ;
  assign n34 = n32 & n33 ;
  assign n35 = n34 ^ x5 ;
  assign n36 = ~n30 & ~n35 ;
  assign n37 = ~n29 & ~n36 ;
  assign n20 = x1 & ~x4 ;
  assign n21 = x5 & n20 ;
  assign n22 = ~x6 & n21 ;
  assign n23 = x7 ^ x6 ;
  assign n24 = n15 & n23 ;
  assign n25 = ~n22 & ~n24 ;
  assign n38 = n37 ^ n25 ;
  assign n39 = n38 ^ n25 ;
  assign n40 = ~x4 & n16 ;
  assign n41 = n27 & n40 ;
  assign n42 = n41 ^ n25 ;
  assign n43 = n42 ^ n25 ;
  assign n44 = ~n39 & ~n43 ;
  assign n45 = n44 ^ n25 ;
  assign n46 = x0 & n45 ;
  assign n47 = n46 ^ n25 ;
  assign n48 = n47 ^ x3 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = n49 ^ n19 ;
  assign n51 = ~x5 & n20 ;
  assign n52 = n16 & n51 ;
  assign n53 = x0 & ~n52 ;
  assign n54 = x5 & n10 ;
  assign n55 = ~x0 & ~n54 ;
  assign n56 = x1 & ~n55 ;
  assign n57 = x4 & ~x7 ;
  assign n58 = ~n20 & ~n57 ;
  assign n59 = ~x4 & x7 ;
  assign n60 = x5 & x6 ;
  assign n61 = ~n59 & n60 ;
  assign n62 = n58 & n61 ;
  assign n63 = ~n56 & ~n62 ;
  assign n64 = n63 ^ n53 ;
  assign n65 = ~n53 & n64 ;
  assign n66 = n65 ^ n47 ;
  assign n67 = n66 ^ n53 ;
  assign n68 = ~n50 & n67 ;
  assign n69 = n68 ^ n65 ;
  assign n70 = n69 ^ n53 ;
  assign n71 = ~n19 & ~n70 ;
  assign n72 = n71 ^ n19 ;
  assign n73 = n72 ^ x2 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = x5 & ~x6 ;
  assign n76 = n58 ^ x1 ;
  assign n77 = n76 ^ n58 ;
  assign n78 = n58 ^ n10 ;
  assign n79 = n78 ^ n58 ;
  assign n80 = n77 & n79 ;
  assign n81 = n80 ^ n58 ;
  assign n82 = ~x0 & ~n81 ;
  assign n83 = n82 ^ n58 ;
  assign n84 = n75 & ~n83 ;
  assign n85 = x7 ^ x5 ;
  assign n86 = n85 ^ x4 ;
  assign n87 = n86 ^ x0 ;
  assign n88 = n87 ^ x7 ;
  assign n97 = n88 ^ n85 ;
  assign n94 = x4 ^ x1 ;
  assign n98 = n97 ^ n94 ;
  assign n99 = n98 ^ n94 ;
  assign n90 = x7 ^ x0 ;
  assign n100 = n90 ^ n85 ;
  assign n101 = n100 ^ n94 ;
  assign n102 = ~n99 & n101 ;
  assign n89 = n85 ^ x7 ;
  assign n91 = n90 ^ n89 ;
  assign n92 = n91 ^ n85 ;
  assign n93 = n92 ^ n88 ;
  assign n95 = n94 ^ n93 ;
  assign n96 = n88 & n95 ;
  assign n103 = n102 ^ n96 ;
  assign n104 = n103 ^ n88 ;
  assign n105 = n96 ^ n94 ;
  assign n106 = n105 ^ n98 ;
  assign n107 = ~n94 & ~n106 ;
  assign n108 = n107 ^ n96 ;
  assign n109 = n104 & n108 ;
  assign n110 = n109 ^ n102 ;
  assign n111 = n110 ^ n107 ;
  assign n112 = n111 ^ n88 ;
  assign n113 = n112 ^ n94 ;
  assign n114 = n113 ^ n98 ;
  assign n115 = n114 ^ x6 ;
  assign n116 = n115 ^ n114 ;
  assign n117 = n116 ^ n84 ;
  assign n118 = x0 & ~x1 ;
  assign n119 = n118 ^ n59 ;
  assign n120 = n59 & n119 ;
  assign n121 = n120 ^ n114 ;
  assign n122 = n121 ^ n59 ;
  assign n123 = n117 & ~n122 ;
  assign n124 = n123 ^ n120 ;
  assign n125 = n124 ^ n59 ;
  assign n126 = ~n84 & n125 ;
  assign n127 = n126 ^ n84 ;
  assign n128 = ~x3 & n127 ;
  assign n129 = ~x1 & ~n30 ;
  assign n130 = x0 & ~n129 ;
  assign n131 = x6 ^ x5 ;
  assign n132 = x5 ^ x0 ;
  assign n133 = n132 ^ x5 ;
  assign n134 = n131 & ~n133 ;
  assign n135 = n134 ^ x5 ;
  assign n136 = ~n59 & n135 ;
  assign n137 = ~n130 & ~n136 ;
  assign n138 = x1 & ~n15 ;
  assign n139 = ~x0 & x4 ;
  assign n140 = ~x6 & ~n139 ;
  assign n141 = ~x5 & n140 ;
  assign n142 = ~n138 & ~n141 ;
  assign n143 = x7 & ~n142 ;
  assign n144 = x5 ^ x3 ;
  assign n145 = n57 ^ n20 ;
  assign n146 = n20 ^ x5 ;
  assign n147 = n146 ^ n20 ;
  assign n148 = n145 & n147 ;
  assign n149 = n148 ^ n20 ;
  assign n150 = ~n144 & n149 ;
  assign n151 = n150 ^ x3 ;
  assign n152 = ~n143 & n151 ;
  assign n153 = n137 & n152 ;
  assign n154 = ~n128 & ~n153 ;
  assign n155 = n154 ^ n72 ;
  assign n156 = n74 & ~n155 ;
  assign n157 = n156 ^ n72 ;
  assign n158 = ~n14 & ~n157 ;
  assign y0 = ~n158 ;
endmodule
