module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 ;
  assign n25 = ~x10 & ~x11 ;
  assign n37 = ~x7 & ~x8 ;
  assign n38 = x7 & x8 ;
  assign n39 = ~n37 & ~n38 ;
  assign n57 = x13 & ~n39 ;
  assign n58 = ~x14 & ~n57 ;
  assign n26 = x2 & ~x23 ;
  assign n27 = x3 & ~n26 ;
  assign n28 = x4 & ~n27 ;
  assign n29 = x1 & ~n28 ;
  assign n30 = ~x21 & x22 ;
  assign n31 = x19 & ~n30 ;
  assign n32 = x20 & ~n31 ;
  assign n33 = x17 & ~n32 ;
  assign n34 = x18 & ~n33 ;
  assign n35 = x16 & ~n34 ;
  assign n36 = ~n29 & ~n35 ;
  assign n40 = x5 & ~n39 ;
  assign n41 = x0 & ~n40 ;
  assign n42 = x14 & n41 ;
  assign n43 = n36 & n42 ;
  assign n59 = n58 ^ n43 ;
  assign n60 = n59 ^ n43 ;
  assign n44 = ~x2 & x23 ;
  assign n45 = ~x3 & ~n44 ;
  assign n46 = ~x4 & ~n45 ;
  assign n47 = ~x1 & ~n46 ;
  assign n48 = x21 & ~x22 ;
  assign n49 = ~x19 & ~n48 ;
  assign n50 = ~x20 & ~n49 ;
  assign n51 = ~x17 & ~n50 ;
  assign n52 = ~x18 & ~n51 ;
  assign n53 = ~x16 & ~n52 ;
  assign n54 = ~n47 & ~n53 ;
  assign n55 = n54 ^ n43 ;
  assign n56 = n55 ^ n43 ;
  assign n61 = n60 ^ n56 ;
  assign n62 = n43 ^ x0 ;
  assign n63 = n62 ^ n43 ;
  assign n64 = n63 ^ n60 ;
  assign n65 = n60 & ~n64 ;
  assign n66 = n65 ^ n60 ;
  assign n67 = n61 & n66 ;
  assign n68 = n67 ^ n65 ;
  assign n69 = n68 ^ n43 ;
  assign n70 = n69 ^ n60 ;
  assign n71 = x9 & n70 ;
  assign n72 = n71 ^ n43 ;
  assign n73 = n25 & n72 ;
  assign n74 = ~x6 & n73 ;
  assign n108 = ~x12 & x15 ;
  assign n109 = n36 & n108 ;
  assign n110 = x0 & n109 ;
  assign n111 = ~x0 & ~x15 ;
  assign n112 = x12 & n111 ;
  assign n113 = n54 & n112 ;
  assign n114 = ~n37 & ~n113 ;
  assign n115 = ~n110 & n114 ;
  assign n75 = x0 & ~x5 ;
  assign n76 = x13 & n75 ;
  assign n77 = n36 & n76 ;
  assign n78 = x5 & ~x13 ;
  assign n79 = ~x0 & n78 ;
  assign n80 = n54 & n79 ;
  assign n116 = n37 & ~n80 ;
  assign n117 = ~n77 & n116 ;
  assign n118 = ~n115 & ~n117 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n81 ^ n25 ;
  assign n83 = n82 ^ n77 ;
  assign n88 = n83 ^ n81 ;
  assign n89 = n88 ^ n77 ;
  assign n90 = n89 ^ n77 ;
  assign n91 = n81 ^ x9 ;
  assign n92 = n91 ^ n81 ;
  assign n93 = n92 ^ n77 ;
  assign n94 = ~n90 & ~n93 ;
  assign n84 = n81 ^ x14 ;
  assign n85 = n84 ^ n83 ;
  assign n86 = n85 ^ n77 ;
  assign n87 = ~n83 & n86 ;
  assign n95 = n94 ^ n87 ;
  assign n96 = n95 ^ n83 ;
  assign n97 = n87 ^ n77 ;
  assign n98 = n97 ^ n89 ;
  assign n99 = ~n77 & ~n98 ;
  assign n100 = n99 ^ n87 ;
  assign n101 = ~n96 & n100 ;
  assign n102 = n101 ^ n94 ;
  assign n103 = n102 ^ n99 ;
  assign n104 = n103 ^ n83 ;
  assign n105 = n104 ^ n77 ;
  assign n106 = n105 ^ n89 ;
  assign n107 = n106 ^ n80 ;
  assign n119 = n118 ^ n107 ;
  assign n120 = n119 ^ x6 ;
  assign n127 = n120 ^ n119 ;
  assign n121 = n120 ^ n37 ;
  assign n122 = n121 ^ n119 ;
  assign n123 = n120 ^ n118 ;
  assign n124 = n123 ^ n37 ;
  assign n125 = n124 ^ n122 ;
  assign n126 = ~n122 & ~n125 ;
  assign n128 = n127 ^ n126 ;
  assign n129 = n128 ^ n122 ;
  assign n130 = n119 ^ n38 ;
  assign n131 = n126 ^ n122 ;
  assign n132 = ~n130 & ~n131 ;
  assign n133 = n132 ^ n119 ;
  assign n134 = ~n129 & n133 ;
  assign n135 = n134 ^ n119 ;
  assign n136 = n135 ^ n107 ;
  assign n137 = n136 ^ n119 ;
  assign n138 = ~n74 & ~n137 ;
  assign y0 = ~n138 ;
endmodule
