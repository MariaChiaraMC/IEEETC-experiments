module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n12 = x7 ^ x6 ;
  assign n17 = n12 ^ x7 ;
  assign n18 = n17 ^ x7 ;
  assign n19 = ~n17 & ~n18 ;
  assign n9 = x7 ^ x4 ;
  assign n10 = n9 ^ x5 ;
  assign n11 = n10 ^ n9 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = n13 ^ x7 ;
  assign n15 = ~n11 & n14 ;
  assign n22 = n19 ^ n15 ;
  assign n16 = n15 ^ x2 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = ~n16 & ~n20 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = ~x2 & n23 ;
  assign n25 = n24 ^ n15 ;
  assign n26 = n25 ^ n19 ;
  assign n27 = n26 ^ n21 ;
  assign n28 = ~x1 & ~n27 ;
  assign n29 = ~x0 & ~n28 ;
  assign n30 = ~x3 & n29 ;
  assign y0 = n30 ;
endmodule
