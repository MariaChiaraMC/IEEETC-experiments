module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 ;
  assign n10 = ~x1 & ~x2 ;
  assign n11 = ~x3 & n10 ;
  assign n12 = ~x7 & x8 ;
  assign n13 = x4 & x5 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = n13 ^ x0 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = ~n15 & ~n17 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = x6 & n19 ;
  assign n21 = n20 ^ n13 ;
  assign n22 = n12 & n21 ;
  assign n23 = x0 & ~x8 ;
  assign n24 = x7 ^ x6 ;
  assign n25 = n24 ^ x7 ;
  assign n26 = ~x4 & ~x5 ;
  assign n27 = n26 ^ x7 ;
  assign n28 = n25 & ~n27 ;
  assign n29 = n28 ^ x7 ;
  assign n30 = n23 & ~n29 ;
  assign n31 = ~n22 & ~n30 ;
  assign n32 = n11 & ~n31 ;
  assign n34 = ~x4 & ~x8 ;
  assign n35 = x2 ^ x1 ;
  assign n36 = x1 ^ x0 ;
  assign n37 = n36 ^ n35 ;
  assign n39 = ~x3 & x5 ;
  assign n38 = x3 & ~x5 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = n39 ^ x2 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = n40 & n42 ;
  assign n44 = n43 ^ n39 ;
  assign n45 = n44 ^ n35 ;
  assign n46 = ~n37 & ~n45 ;
  assign n47 = n46 ^ n43 ;
  assign n48 = n47 ^ n39 ;
  assign n49 = n48 ^ n36 ;
  assign n50 = ~n35 & n49 ;
  assign n51 = n50 ^ n35 ;
  assign n52 = ~n34 & ~n51 ;
  assign n53 = x6 & x8 ;
  assign n54 = ~x3 & n53 ;
  assign n55 = x0 & n10 ;
  assign n56 = n54 & n55 ;
  assign n57 = ~n52 & ~n56 ;
  assign n33 = x7 ^ x0 ;
  assign n58 = n57 ^ n33 ;
  assign n59 = n58 ^ x7 ;
  assign n60 = n59 ^ n58 ;
  assign n61 = n60 ^ n33 ;
  assign n69 = ~x1 & ~x6 ;
  assign n70 = ~n54 & ~n69 ;
  assign n71 = ~x4 & x5 ;
  assign n72 = ~n70 & n71 ;
  assign n73 = x4 & x8 ;
  assign n74 = ~x5 & x6 ;
  assign n75 = x3 & x5 ;
  assign n76 = ~n74 & ~n75 ;
  assign n77 = n73 & ~n76 ;
  assign n78 = n77 ^ x1 ;
  assign n79 = n78 ^ n77 ;
  assign n80 = ~x5 & x8 ;
  assign n81 = ~x6 & ~n80 ;
  assign n82 = ~x4 & ~n53 ;
  assign n83 = ~n81 & n82 ;
  assign n84 = n83 ^ n77 ;
  assign n85 = n79 & n84 ;
  assign n86 = n85 ^ n77 ;
  assign n87 = ~n72 & ~n86 ;
  assign n88 = ~x7 & ~n87 ;
  assign n65 = x4 & ~x8 ;
  assign n89 = ~x3 & ~x5 ;
  assign n90 = n65 & n89 ;
  assign n91 = n69 & n90 ;
  assign n92 = ~n88 & ~n91 ;
  assign n62 = x1 & x6 ;
  assign n63 = ~n34 & ~n62 ;
  assign n64 = n39 & ~n63 ;
  assign n66 = x6 & n65 ;
  assign n67 = ~n38 & n66 ;
  assign n68 = ~n64 & ~n67 ;
  assign n93 = n92 ^ n68 ;
  assign n94 = n93 ^ n92 ;
  assign n95 = n92 ^ x7 ;
  assign n96 = n95 ^ n92 ;
  assign n97 = ~n94 & ~n96 ;
  assign n98 = n97 ^ n92 ;
  assign n99 = ~x2 & ~n98 ;
  assign n100 = n99 ^ n92 ;
  assign n101 = n100 ^ n58 ;
  assign n102 = n101 ^ n60 ;
  assign n103 = n102 ^ n61 ;
  assign n104 = n61 & ~n103 ;
  assign n105 = n104 ^ n100 ;
  assign n106 = ~x2 & x3 ;
  assign n107 = ~x5 & ~x8 ;
  assign n108 = n69 & n107 ;
  assign n109 = ~x8 & n26 ;
  assign n110 = n109 ^ x7 ;
  assign n111 = n110 ^ n109 ;
  assign n112 = n109 ^ x6 ;
  assign n113 = n112 ^ n110 ;
  assign n114 = n113 ^ x1 ;
  assign n115 = n114 ^ x1 ;
  assign n116 = n115 ^ n109 ;
  assign n117 = ~n111 & ~n116 ;
  assign n118 = n117 ^ n115 ;
  assign n119 = n115 ^ x4 ;
  assign n120 = n119 ^ x5 ;
  assign n121 = n120 ^ n119 ;
  assign n122 = n119 ^ n115 ;
  assign n123 = n122 ^ n114 ;
  assign n124 = n121 & ~n123 ;
  assign n125 = n124 ^ n115 ;
  assign n126 = n114 ^ n110 ;
  assign n127 = n126 ^ n109 ;
  assign n128 = n127 ^ n118 ;
  assign n129 = ~n125 & ~n128 ;
  assign n130 = n129 ^ n111 ;
  assign n131 = ~n118 & ~n130 ;
  assign n132 = n131 ^ n129 ;
  assign n133 = n132 ^ x7 ;
  assign n134 = n133 ^ n111 ;
  assign n135 = ~n108 & ~n134 ;
  assign n136 = n106 & ~n135 ;
  assign n137 = x5 & ~x8 ;
  assign n138 = ~n81 & ~n137 ;
  assign n139 = ~x4 & ~n138 ;
  assign n140 = x4 ^ x1 ;
  assign n141 = n140 ^ x5 ;
  assign n143 = n141 ^ x4 ;
  assign n142 = n141 ^ x6 ;
  assign n144 = n143 ^ n142 ;
  assign n150 = n144 ^ n141 ;
  assign n151 = n150 ^ n143 ;
  assign n152 = n151 ^ n143 ;
  assign n153 = n141 ^ x5 ;
  assign n154 = n153 ^ n141 ;
  assign n155 = n154 ^ n143 ;
  assign n156 = n152 & n155 ;
  assign n145 = ~x3 & ~x7 ;
  assign n146 = n145 ^ n141 ;
  assign n147 = n146 ^ n144 ;
  assign n148 = n147 ^ n143 ;
  assign n149 = n144 & ~n148 ;
  assign n157 = n156 ^ n149 ;
  assign n158 = n157 ^ n144 ;
  assign n159 = n149 ^ n143 ;
  assign n160 = n159 ^ n151 ;
  assign n161 = ~n143 & n160 ;
  assign n162 = n161 ^ n149 ;
  assign n163 = n158 & n162 ;
  assign n164 = n163 ^ n156 ;
  assign n165 = n164 ^ n161 ;
  assign n166 = n165 ^ n144 ;
  assign n167 = n166 ^ n143 ;
  assign n168 = n167 ^ n151 ;
  assign n169 = n168 ^ x4 ;
  assign n170 = ~n139 & ~n169 ;
  assign n171 = x7 ^ x5 ;
  assign n172 = x3 & ~n171 ;
  assign n173 = n172 ^ x5 ;
  assign n174 = n170 & n173 ;
  assign n175 = ~n136 & ~n174 ;
  assign n176 = n175 ^ n58 ;
  assign n177 = n176 ^ n60 ;
  assign n178 = n176 ^ n100 ;
  assign n179 = ~n177 & ~n178 ;
  assign n180 = n179 ^ n175 ;
  assign n181 = n180 ^ n61 ;
  assign n182 = x1 & ~x2 ;
  assign n183 = n107 & n182 ;
  assign n184 = ~x3 & n183 ;
  assign n185 = ~x2 & n13 ;
  assign n186 = ~n137 & ~n185 ;
  assign n187 = ~x1 & x3 ;
  assign n188 = ~n186 & n187 ;
  assign n189 = x2 & n137 ;
  assign n190 = ~n11 & ~n189 ;
  assign n191 = n190 ^ x4 ;
  assign n192 = n191 ^ n190 ;
  assign n193 = n192 ^ n188 ;
  assign n194 = n39 ^ n35 ;
  assign n195 = n38 ^ x2 ;
  assign n196 = n195 ^ n38 ;
  assign n197 = n196 ^ n194 ;
  assign n198 = n39 ^ x3 ;
  assign n199 = ~n39 & n198 ;
  assign n200 = n199 ^ n38 ;
  assign n201 = n200 ^ n39 ;
  assign n202 = ~n197 & n201 ;
  assign n203 = n202 ^ n199 ;
  assign n204 = n203 ^ n39 ;
  assign n205 = n194 & ~n204 ;
  assign n206 = n205 ^ x2 ;
  assign n207 = n206 ^ x8 ;
  assign n208 = x8 & n207 ;
  assign n209 = n208 ^ n190 ;
  assign n210 = n209 ^ x8 ;
  assign n211 = ~n193 & ~n210 ;
  assign n212 = n211 ^ n208 ;
  assign n213 = n212 ^ x8 ;
  assign n214 = ~n188 & n213 ;
  assign n215 = n214 ^ n188 ;
  assign n216 = ~n184 & ~n215 ;
  assign n217 = ~x6 & ~n216 ;
  assign n218 = n62 & n65 ;
  assign n219 = x3 & n218 ;
  assign n220 = n53 ^ x8 ;
  assign n221 = ~n26 & ~n220 ;
  assign n222 = n221 ^ x8 ;
  assign n223 = n182 & ~n222 ;
  assign n224 = n137 ^ n106 ;
  assign n225 = ~x1 & ~x4 ;
  assign n226 = n225 ^ n137 ;
  assign n227 = n226 ^ n225 ;
  assign n228 = ~x1 & x6 ;
  assign n229 = n80 & n228 ;
  assign n230 = n229 ^ n225 ;
  assign n231 = ~n227 & ~n230 ;
  assign n232 = n231 ^ n225 ;
  assign n233 = n224 & n232 ;
  assign n234 = n233 ^ n106 ;
  assign n235 = ~n223 & ~n234 ;
  assign n236 = x2 & x6 ;
  assign n237 = n225 ^ x8 ;
  assign n238 = n225 ^ n75 ;
  assign n239 = n238 ^ n75 ;
  assign n240 = n239 ^ n237 ;
  assign n241 = n39 ^ x4 ;
  assign n242 = n39 & n241 ;
  assign n243 = n242 ^ n75 ;
  assign n244 = n243 ^ n39 ;
  assign n245 = n240 & ~n244 ;
  assign n246 = n245 ^ n242 ;
  assign n247 = n246 ^ n39 ;
  assign n248 = ~n237 & n247 ;
  assign n249 = n248 ^ n225 ;
  assign n250 = n236 & n249 ;
  assign n251 = n235 & ~n250 ;
  assign n252 = ~n219 & n251 ;
  assign n253 = ~n217 & n252 ;
  assign n254 = n175 ^ n61 ;
  assign n255 = n253 & ~n254 ;
  assign n256 = n255 ^ n253 ;
  assign n257 = n256 ^ n100 ;
  assign n258 = n257 ^ n60 ;
  assign n259 = n258 ^ n61 ;
  assign n260 = ~n181 & n259 ;
  assign n261 = n260 ^ n60 ;
  assign n262 = n261 ^ n61 ;
  assign n263 = ~n105 & ~n262 ;
  assign n264 = n263 ^ n260 ;
  assign n265 = n264 ^ n60 ;
  assign n266 = n265 ^ n61 ;
  assign n267 = n266 ^ x0 ;
  assign n268 = ~n32 & ~n267 ;
  assign y0 = ~n268 ;
endmodule
