module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 ;
  assign n9 = ~x1 & ~x5 ;
  assign n10 = ~x4 & ~x7 ;
  assign n11 = ~x3 & ~n10 ;
  assign n12 = x6 ^ x4 ;
  assign n13 = x2 & n12 ;
  assign n14 = ~n11 & ~n13 ;
  assign n15 = n9 & ~n14 ;
  assign n16 = x6 & x7 ;
  assign n17 = x5 & n16 ;
  assign n18 = ~x3 & ~n17 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = x5 & ~x7 ;
  assign n22 = x6 & n21 ;
  assign n23 = n22 ^ n18 ;
  assign n24 = n23 ^ n18 ;
  assign n25 = ~n20 & n24 ;
  assign n26 = n25 ^ n18 ;
  assign n27 = ~x1 & ~n26 ;
  assign n28 = n27 ^ n18 ;
  assign n30 = x5 ^ x3 ;
  assign n29 = x4 ^ x1 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n31 ^ x1 ;
  assign n33 = n32 ^ n30 ;
  assign n37 = x7 ^ x1 ;
  assign n38 = n37 ^ n29 ;
  assign n39 = n38 ^ n29 ;
  assign n40 = n39 ^ x1 ;
  assign n34 = n29 ^ x5 ;
  assign n35 = n34 ^ x1 ;
  assign n36 = n35 ^ x1 ;
  assign n41 = n40 ^ n36 ;
  assign n42 = ~n33 & ~n41 ;
  assign n43 = n42 ^ n35 ;
  assign n44 = n43 ^ n36 ;
  assign n45 = x6 ^ x3 ;
  assign n46 = n45 ^ n30 ;
  assign n47 = n46 ^ n35 ;
  assign n48 = n47 ^ n33 ;
  assign n49 = n48 ^ n40 ;
  assign n50 = n46 ^ n30 ;
  assign n53 = n50 ^ n35 ;
  assign n54 = n49 & n53 ;
  assign n51 = n50 ^ n33 ;
  assign n52 = n49 & n51 ;
  assign n55 = n54 ^ n52 ;
  assign n56 = n55 ^ n30 ;
  assign n57 = ~n48 & n56 ;
  assign n58 = n57 ^ n52 ;
  assign n59 = n58 ^ n30 ;
  assign n60 = n59 ^ n35 ;
  assign n61 = n60 ^ n33 ;
  assign n62 = n61 ^ n40 ;
  assign n63 = ~n44 & ~n62 ;
  assign n64 = n63 ^ n30 ;
  assign n65 = n64 ^ n33 ;
  assign n66 = n65 ^ x4 ;
  assign n67 = n66 ^ n32 ;
  assign n68 = n28 & ~n67 ;
  assign n69 = n22 ^ x6 ;
  assign n70 = n69 ^ n22 ;
  assign n71 = ~x1 & ~x4 ;
  assign n72 = x7 & n71 ;
  assign n73 = ~n9 & ~n72 ;
  assign n74 = n73 ^ n22 ;
  assign n75 = n74 ^ n22 ;
  assign n76 = ~n70 & ~n75 ;
  assign n77 = n76 ^ n22 ;
  assign n78 = ~x3 & n77 ;
  assign n79 = n78 ^ n22 ;
  assign n80 = n68 & ~n79 ;
  assign n81 = n80 ^ x2 ;
  assign n82 = n81 ^ n80 ;
  assign n83 = x3 & x5 ;
  assign n84 = n71 & n83 ;
  assign n85 = n84 ^ n80 ;
  assign n86 = n82 & ~n85 ;
  assign n87 = n86 ^ n80 ;
  assign n88 = ~n15 & n87 ;
  assign n89 = ~x0 & ~n88 ;
  assign y0 = n89 ;
endmodule
