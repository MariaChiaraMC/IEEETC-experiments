module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 ;
  assign n9 = ~x1 & x4 ;
  assign n10 = x2 & x7 ;
  assign n11 = ~x6 & ~n10 ;
  assign n12 = n9 & ~n11 ;
  assign n13 = ~x5 & ~n12 ;
  assign n14 = x0 & ~x3 ;
  assign n15 = ~n13 & n14 ;
  assign n23 = x7 ^ x1 ;
  assign n16 = x6 ^ x1 ;
  assign n24 = n16 ^ x5 ;
  assign n25 = n23 & n24 ;
  assign n17 = n16 ^ x4 ;
  assign n18 = x2 ^ x1 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = n17 & n19 ;
  assign n31 = n25 ^ n20 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = n21 ^ n17 ;
  assign n26 = x4 ^ x1 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = n27 ^ n23 ;
  assign n29 = n28 ^ x5 ;
  assign n30 = n22 & n29 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = n32 ^ n26 ;
  assign n34 = n33 ^ n23 ;
  assign n35 = n34 ^ x5 ;
  assign n36 = x5 & n35 ;
  assign n37 = n36 ^ x5 ;
  assign n38 = n37 ^ x5 ;
  assign n39 = n38 ^ x5 ;
  assign n40 = n15 & ~n39 ;
  assign y0 = n40 ;
endmodule
