module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 ;
  assign n10 = ~x7 & ~x8 ;
  assign n11 = x6 & ~n10 ;
  assign n13 = x4 ^ x1 ;
  assign n12 = x5 ^ x4 ;
  assign n14 = n13 ^ n12 ;
  assign n16 = n14 ^ x0 ;
  assign n15 = n14 ^ x3 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n17 ^ x4 ;
  assign n23 = n18 ^ n16 ;
  assign n24 = n23 ^ n14 ;
  assign n19 = n14 ^ n12 ;
  assign n20 = n19 ^ x4 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = ~n18 & n21 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n25 ^ n20 ;
  assign n27 = n24 ^ x4 ;
  assign n28 = n27 ^ n18 ;
  assign n29 = n28 ^ n20 ;
  assign n31 = n12 ^ x2 ;
  assign n32 = n31 ^ n12 ;
  assign n33 = n32 ^ n12 ;
  assign n34 = ~n29 & ~n33 ;
  assign n30 = n12 & ~n29 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n35 ^ n12 ;
  assign n37 = n36 ^ n32 ;
  assign n38 = n37 ^ n20 ;
  assign n39 = ~x4 & n38 ;
  assign n40 = n39 ^ n34 ;
  assign n41 = n40 ^ n32 ;
  assign n42 = n41 ^ n20 ;
  assign n43 = ~n26 & n42 ;
  assign n44 = n43 ^ n30 ;
  assign n45 = n44 ^ n12 ;
  assign n46 = n45 ^ x5 ;
  assign n47 = ~n11 & ~n46 ;
  assign y0 = n47 ;
endmodule
