module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 ;
  assign n10 = ~x4 & x5 ;
  assign n11 = x4 & ~x8 ;
  assign n12 = ~n10 & ~n11 ;
  assign n13 = x2 & x6 ;
  assign n14 = x4 & x5 ;
  assign n15 = n14 ^ x1 ;
  assign n16 = n15 ^ x1 ;
  assign n17 = x8 ^ x1 ;
  assign n18 = n17 ^ x1 ;
  assign n19 = n16 & ~n18 ;
  assign n20 = n19 ^ x1 ;
  assign n21 = ~x7 & ~n20 ;
  assign n22 = n21 ^ x1 ;
  assign n23 = n13 & ~n22 ;
  assign n24 = ~n12 & n23 ;
  assign n25 = ~x2 & x6 ;
  assign n29 = x7 & x8 ;
  assign n26 = x4 & x7 ;
  assign n27 = ~x7 & x8 ;
  assign n28 = ~n26 & ~n27 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = x1 & ~n30 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = ~x5 & n32 ;
  assign n34 = x5 & ~x7 ;
  assign n35 = x4 & n34 ;
  assign n36 = ~x1 & n35 ;
  assign n37 = ~n33 & ~n36 ;
  assign n38 = n25 & ~n37 ;
  assign n39 = ~x6 & x8 ;
  assign n40 = ~x4 & ~x5 ;
  assign n41 = ~x7 & n40 ;
  assign n42 = x1 & x2 ;
  assign n43 = ~n41 & n42 ;
  assign n44 = n39 & n43 ;
  assign n45 = ~x4 & n34 ;
  assign n46 = n45 ^ x5 ;
  assign n47 = n44 & ~n46 ;
  assign n48 = ~n38 & ~n47 ;
  assign n49 = ~n24 & n48 ;
  assign n62 = ~x6 & ~x7 ;
  assign n138 = ~n26 & ~n62 ;
  assign n139 = x8 & ~n138 ;
  assign n140 = n139 ^ x4 ;
  assign n141 = n140 ^ n139 ;
  assign n55 = x7 & ~x8 ;
  assign n120 = ~x6 & n55 ;
  assign n142 = n139 ^ n120 ;
  assign n143 = n142 ^ n139 ;
  assign n144 = n141 & n143 ;
  assign n145 = n144 ^ n139 ;
  assign n146 = x2 & n145 ;
  assign n147 = n146 ^ n139 ;
  assign n148 = ~x5 & n147 ;
  assign n77 = x6 & ~x8 ;
  assign n78 = ~n14 & ~n41 ;
  assign n79 = n77 & ~n78 ;
  assign n56 = x5 & ~x6 ;
  assign n80 = ~n39 & ~n56 ;
  assign n81 = ~x2 & n34 ;
  assign n82 = ~x4 & ~n29 ;
  assign n83 = ~n81 & n82 ;
  assign n84 = ~n80 & n83 ;
  assign n85 = ~n79 & ~n84 ;
  assign n50 = ~x7 & ~x8 ;
  assign n51 = ~x5 & ~n50 ;
  assign n52 = n13 & ~n51 ;
  assign n53 = ~x2 & ~x5 ;
  assign n54 = x7 & n53 ;
  assign n57 = n55 & n56 ;
  assign n58 = ~n54 & ~n57 ;
  assign n59 = ~n52 & n58 ;
  assign n63 = n62 ^ n59 ;
  assign n64 = n63 ^ n59 ;
  assign n60 = n59 ^ x8 ;
  assign n61 = n60 ^ n59 ;
  assign n65 = n64 ^ n61 ;
  assign n66 = n59 ^ x2 ;
  assign n67 = n66 ^ n59 ;
  assign n68 = n67 ^ n64 ;
  assign n69 = n64 & ~n68 ;
  assign n70 = n69 ^ n64 ;
  assign n71 = ~n65 & n70 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = n72 ^ n59 ;
  assign n74 = n73 ^ n64 ;
  assign n75 = ~x4 & ~n74 ;
  assign n76 = n75 ^ n59 ;
  assign n86 = n85 ^ n76 ;
  assign n87 = n86 ^ n85 ;
  assign n88 = x4 ^ x2 ;
  assign n89 = n88 ^ x4 ;
  assign n90 = n89 ^ x8 ;
  assign n91 = n90 ^ x8 ;
  assign n92 = x8 ^ x6 ;
  assign n93 = n91 ^ n88 ;
  assign n94 = n93 ^ n91 ;
  assign n95 = n92 & ~n94 ;
  assign n96 = n95 ^ x8 ;
  assign n97 = x8 ^ x5 ;
  assign n98 = ~n93 & n97 ;
  assign n99 = n98 ^ n91 ;
  assign n100 = n99 ^ n93 ;
  assign n101 = ~n96 & ~n100 ;
  assign n102 = n91 & n101 ;
  assign n103 = n102 ^ n95 ;
  assign n104 = n103 ^ x2 ;
  assign n105 = x7 & n104 ;
  assign n106 = n105 ^ n85 ;
  assign n107 = n106 ^ n85 ;
  assign n108 = n87 & ~n107 ;
  assign n109 = n108 ^ n85 ;
  assign n110 = x1 & n109 ;
  assign n111 = n110 ^ n85 ;
  assign n112 = n35 & n77 ;
  assign n113 = x6 & ~x7 ;
  assign n114 = ~x5 & ~n113 ;
  assign n115 = ~n39 & ~n55 ;
  assign n116 = n114 & n115 ;
  assign n117 = n116 ^ x4 ;
  assign n118 = n117 ^ n116 ;
  assign n119 = n118 ^ n112 ;
  assign n121 = x6 & x8 ;
  assign n122 = x5 & n121 ;
  assign n123 = ~n120 & ~n122 ;
  assign n124 = n123 ^ x2 ;
  assign n125 = ~n123 & ~n124 ;
  assign n126 = n125 ^ n116 ;
  assign n127 = n126 ^ n123 ;
  assign n128 = n119 & ~n127 ;
  assign n129 = n128 ^ n125 ;
  assign n130 = n129 ^ n123 ;
  assign n131 = ~n112 & ~n130 ;
  assign n132 = n131 ^ n112 ;
  assign n133 = n111 & ~n132 ;
  assign n149 = n148 ^ n133 ;
  assign n150 = n149 ^ n133 ;
  assign n134 = n10 & n27 ;
  assign n135 = n25 & n134 ;
  assign n136 = n135 ^ n133 ;
  assign n137 = n136 ^ n133 ;
  assign n151 = n150 ^ n137 ;
  assign n184 = n26 ^ x2 ;
  assign n185 = n184 ^ x2 ;
  assign n186 = n185 ^ x5 ;
  assign n189 = ~n29 & ~n50 ;
  assign n190 = ~x4 & ~n189 ;
  assign n187 = x4 & ~x6 ;
  assign n188 = ~n55 & ~n187 ;
  assign n191 = n190 ^ n188 ;
  assign n192 = ~x2 & n191 ;
  assign n193 = n192 ^ n188 ;
  assign n194 = ~n186 & ~n193 ;
  assign n195 = n194 ^ n192 ;
  assign n196 = n195 ^ n188 ;
  assign n197 = n196 ^ x2 ;
  assign n198 = x5 & n197 ;
  assign n152 = ~n113 & ~n120 ;
  assign n153 = n10 & ~n121 ;
  assign n154 = ~n27 & n153 ;
  assign n155 = n152 & n154 ;
  assign n157 = n40 & ~n77 ;
  assign n156 = x7 ^ x6 ;
  assign n158 = n157 ^ n156 ;
  assign n159 = n157 ^ x7 ;
  assign n160 = n159 ^ x7 ;
  assign n161 = n160 ^ n158 ;
  assign n162 = x7 ^ x5 ;
  assign n163 = n162 ^ x4 ;
  assign n164 = x4 & ~n163 ;
  assign n165 = n164 ^ x7 ;
  assign n166 = n165 ^ x4 ;
  assign n167 = ~n161 & ~n166 ;
  assign n168 = n167 ^ n164 ;
  assign n169 = n168 ^ x4 ;
  assign n170 = n158 & n169 ;
  assign n171 = n170 ^ n157 ;
  assign n172 = n171 ^ x2 ;
  assign n173 = n172 ^ n171 ;
  assign n174 = n173 ^ n155 ;
  assign n175 = n62 ^ x5 ;
  assign n176 = ~x5 & ~n175 ;
  assign n177 = n176 ^ n171 ;
  assign n178 = n177 ^ x5 ;
  assign n179 = n174 & ~n178 ;
  assign n180 = n179 ^ n176 ;
  assign n181 = n180 ^ x5 ;
  assign n182 = ~n155 & ~n181 ;
  assign n183 = n182 ^ n155 ;
  assign n199 = n198 ^ n183 ;
  assign n200 = n199 ^ n183 ;
  assign n202 = n14 & n29 ;
  assign n203 = x2 & ~x4 ;
  assign n204 = n50 & n203 ;
  assign n205 = ~n202 & ~n204 ;
  assign n201 = ~x2 & ~x4 ;
  assign n206 = n205 ^ n201 ;
  assign n207 = n206 ^ n205 ;
  assign n208 = n205 ^ n55 ;
  assign n209 = n208 ^ n205 ;
  assign n210 = n207 & n209 ;
  assign n211 = n210 ^ n205 ;
  assign n212 = ~x6 & ~n211 ;
  assign n213 = n212 ^ n205 ;
  assign n214 = n213 ^ n183 ;
  assign n215 = n214 ^ n183 ;
  assign n216 = ~n200 & n215 ;
  assign n217 = n216 ^ n183 ;
  assign n218 = x1 & ~n217 ;
  assign n219 = n218 ^ n183 ;
  assign n220 = n219 ^ n133 ;
  assign n221 = n220 ^ n133 ;
  assign n222 = n221 ^ n150 ;
  assign n223 = ~n150 & n222 ;
  assign n224 = n223 ^ n150 ;
  assign n225 = n151 & ~n224 ;
  assign n226 = n225 ^ n223 ;
  assign n227 = n226 ^ n133 ;
  assign n228 = n227 ^ n150 ;
  assign n229 = x3 & ~n228 ;
  assign n230 = n229 ^ n133 ;
  assign n231 = n49 & n230 ;
  assign n232 = ~x0 & ~n231 ;
  assign n233 = ~x2 & ~x3 ;
  assign n234 = x6 & x7 ;
  assign n235 = n234 ^ x6 ;
  assign n236 = ~x5 & ~n235 ;
  assign n237 = n236 ^ x6 ;
  assign n238 = x0 & ~n237 ;
  assign n239 = n11 & n238 ;
  assign n240 = ~x6 & x7 ;
  assign n241 = x5 & ~n240 ;
  assign n242 = ~n189 & n241 ;
  assign n243 = ~n11 & ~n121 ;
  assign n244 = ~x7 & n243 ;
  assign n245 = ~n242 & ~n244 ;
  assign n246 = x0 & ~n245 ;
  assign n247 = n246 ^ n239 ;
  assign n248 = ~x0 & ~x5 ;
  assign n249 = ~n234 & ~n248 ;
  assign n250 = x8 & ~n249 ;
  assign n251 = n250 ^ x4 ;
  assign n252 = n251 ^ n250 ;
  assign n253 = n97 ^ x5 ;
  assign n254 = n56 ^ x5 ;
  assign n255 = n254 ^ x5 ;
  assign n256 = n253 & n255 ;
  assign n257 = n256 ^ x5 ;
  assign n258 = x7 & ~n257 ;
  assign n259 = n258 ^ x5 ;
  assign n260 = ~x0 & ~n259 ;
  assign n261 = n260 ^ n250 ;
  assign n262 = n252 & n261 ;
  assign n263 = n262 ^ n250 ;
  assign n264 = n263 ^ n239 ;
  assign n265 = n247 & n264 ;
  assign n266 = n265 ^ n262 ;
  assign n267 = n266 ^ n250 ;
  assign n268 = n267 ^ n246 ;
  assign n269 = ~n239 & n268 ;
  assign n270 = n269 ^ n239 ;
  assign n271 = n233 & n270 ;
  assign n272 = ~x1 & n271 ;
  assign n273 = ~n232 & ~n272 ;
  assign y0 = ~n273 ;
endmodule
