module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 ;
  assign n26 = x5 & ~x6 ;
  assign n11 = ~x3 & x9 ;
  assign n12 = ~x7 & n11 ;
  assign n27 = n26 ^ n12 ;
  assign n35 = n27 ^ n12 ;
  assign n13 = x1 & x4 ;
  assign n14 = n13 ^ x3 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = n13 ^ x0 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n15 & n17 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = x6 & n19 ;
  assign n21 = n20 ^ n13 ;
  assign n22 = ~x5 & n21 ;
  assign n23 = ~x7 & ~n22 ;
  assign n24 = ~x9 & ~n23 ;
  assign n25 = n24 ^ n12 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ n12 ;
  assign n31 = n28 ^ x8 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n30 & ~n33 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = ~x3 & x6 ;
  assign n39 = x4 & n38 ;
  assign n40 = x7 & ~n39 ;
  assign n41 = ~x5 & ~n40 ;
  assign n42 = n41 ^ n12 ;
  assign n43 = n34 ^ n30 ;
  assign n44 = ~n42 & n43 ;
  assign n45 = n44 ^ n12 ;
  assign n46 = n37 & ~n45 ;
  assign n47 = n46 ^ n12 ;
  assign n48 = n47 ^ n26 ;
  assign n49 = n48 ^ n12 ;
  assign n50 = ~x2 & n49 ;
  assign y0 = n50 ;
endmodule
