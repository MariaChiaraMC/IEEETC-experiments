module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 ;
  assign n23 = x13 ^ x0 ;
  assign n31 = n23 ^ x0 ;
  assign n32 = n31 ^ x0 ;
  assign n33 = ~n31 & ~n32 ;
  assign n22 = x12 ^ x0 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n24 ^ n23 ;
  assign n28 = n27 ^ x0 ;
  assign n29 = n26 & n28 ;
  assign n36 = n33 ^ n29 ;
  assign n30 = n29 ^ x6 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = ~n30 & ~n34 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = ~x6 & n37 ;
  assign n39 = n38 ^ n29 ;
  assign n40 = n39 ^ n33 ;
  assign n41 = n40 ^ n35 ;
  assign n42 = n41 ^ x13 ;
  assign n43 = ~x11 & ~n42 ;
  assign n44 = n43 ^ x3 ;
  assign n45 = n44 ^ n43 ;
  assign n15 = ~x12 & ~x13 ;
  assign n16 = x4 & ~x8 ;
  assign n17 = n15 & ~n16 ;
  assign n46 = n43 ^ n17 ;
  assign n47 = n46 ^ n43 ;
  assign n48 = n45 & n47 ;
  assign n49 = n48 ^ n43 ;
  assign n50 = ~x9 & ~n49 ;
  assign n51 = n50 ^ n43 ;
  assign n52 = n51 ^ x11 ;
  assign n18 = ~x9 & n17 ;
  assign n19 = ~x6 & x10 ;
  assign n20 = n18 & n19 ;
  assign n21 = n20 ^ x11 ;
  assign n53 = n52 ^ n21 ;
  assign n54 = n53 ^ x10 ;
  assign n55 = n54 ^ n53 ;
  assign n56 = n53 ^ n21 ;
  assign n57 = n56 ^ x11 ;
  assign n58 = ~n55 & ~n57 ;
  assign n59 = n58 ^ n21 ;
  assign n60 = x9 & n15 ;
  assign n61 = n21 & n60 ;
  assign n62 = n61 ^ x11 ;
  assign n63 = n59 & n62 ;
  assign n64 = n63 ^ n61 ;
  assign n65 = x11 & n64 ;
  assign n66 = n65 ^ n58 ;
  assign n67 = n66 ^ n20 ;
  assign n68 = n67 ^ n21 ;
  assign n69 = ~x5 & n68 ;
  assign y0 = n69 ;
endmodule
