module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 ;
  assign n17 = ~x3 & x4 ;
  assign n18 = ~x0 & ~n17 ;
  assign n19 = x5 ^ x2 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = x6 ^ x5 ;
  assign n22 = x5 ^ x3 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n21 & ~n23 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = n20 & ~n26 ;
  assign n28 = n27 ^ n24 ;
  assign n29 = n28 ^ n21 ;
  assign n30 = ~n18 & n29 ;
  assign n31 = n30 ^ n18 ;
  assign n8 = x5 & x6 ;
  assign n9 = n8 ^ x2 ;
  assign n10 = n9 ^ n8 ;
  assign n11 = n8 ^ x3 ;
  assign n12 = n11 ^ n8 ;
  assign n13 = ~n10 & n12 ;
  assign n14 = n13 ^ n8 ;
  assign n15 = x0 & n14 ;
  assign n16 = n15 ^ n8 ;
  assign n32 = n31 ^ n16 ;
  assign n33 = n32 ^ n16 ;
  assign n34 = x5 & ~x6 ;
  assign n35 = ~x4 & ~n34 ;
  assign n36 = ~x2 & ~n35 ;
  assign n37 = n36 ^ n16 ;
  assign n38 = n37 ^ n16 ;
  assign n39 = ~n33 & ~n38 ;
  assign n40 = n39 ^ n16 ;
  assign n41 = x1 & ~n40 ;
  assign n42 = n41 ^ n16 ;
  assign y0 = ~n42 ;
endmodule
