module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
  assign n17 = x13 & x14 ;
  assign n18 = ~x11 & ~x12 ;
  assign n19 = ~n17 & n18 ;
  assign n20 = x8 & x15 ;
  assign n21 = x9 ^ x8 ;
  assign n22 = x10 ^ x8 ;
  assign n23 = ~n21 & ~n22 ;
  assign n24 = n23 ^ n19 ;
  assign n25 = n20 & n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n19 & n26 ;
  assign n28 = n27 ^ n19 ;
  assign n30 = ~x13 & ~x14 ;
  assign n29 = ~x8 & ~x15 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n28 & n31 ;
  assign n33 = ~x7 & ~n32 ;
  assign n34 = ~x6 & ~n33 ;
  assign n35 = ~x0 & ~n34 ;
  assign y0 = ~n35 ;
endmodule
