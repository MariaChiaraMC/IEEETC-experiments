module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 ;
  assign n10 = ~x1 & x5 ;
  assign n11 = ~x6 & ~x8 ;
  assign n12 = n10 & n11 ;
  assign n13 = ~x0 & n12 ;
  assign n14 = x4 & x5 ;
  assign n15 = ~x8 & n14 ;
  assign n16 = x0 & ~x7 ;
  assign n17 = n15 & n16 ;
  assign n18 = x2 & x6 ;
  assign n19 = ~x1 & ~x7 ;
  assign n20 = n14 & n19 ;
  assign n21 = ~n18 & n20 ;
  assign n22 = ~n17 & ~n21 ;
  assign n23 = x1 & ~x5 ;
  assign n24 = ~x0 & ~n18 ;
  assign n25 = n23 & n24 ;
  assign n26 = ~x8 & n25 ;
  assign n27 = n22 & ~n26 ;
  assign n28 = ~n13 & n27 ;
  assign n29 = x6 & x8 ;
  assign n30 = x4 & n10 ;
  assign n31 = ~n29 & n30 ;
  assign n32 = ~x2 & n31 ;
  assign n33 = ~n10 & ~n23 ;
  assign n34 = x6 & ~n10 ;
  assign n35 = ~n33 & ~n34 ;
  assign n36 = ~x4 & n24 ;
  assign n37 = n35 & n36 ;
  assign n38 = ~n32 & ~n37 ;
  assign n39 = x4 & x8 ;
  assign n40 = ~x1 & ~x5 ;
  assign n41 = n39 & n40 ;
  assign n42 = x7 ^ x6 ;
  assign n43 = x2 & n42 ;
  assign n44 = n41 & n43 ;
  assign n45 = n38 & ~n44 ;
  assign n46 = x2 & x7 ;
  assign n56 = x0 & ~x4 ;
  assign n57 = n56 ^ n46 ;
  assign n48 = x4 & x7 ;
  assign n49 = ~x2 & ~x5 ;
  assign n50 = ~n48 & n49 ;
  assign n51 = ~x4 & ~x6 ;
  assign n52 = x5 & ~n51 ;
  assign n53 = n43 & n52 ;
  assign n54 = ~n50 & ~n53 ;
  assign n47 = x1 & x8 ;
  assign n55 = n54 ^ n47 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = n55 ^ n54 ;
  assign n60 = n59 ^ n46 ;
  assign n61 = ~n58 & n60 ;
  assign n62 = n61 ^ n54 ;
  assign n63 = ~x5 & ~x6 ;
  assign n64 = n54 & ~n63 ;
  assign n65 = n64 ^ n46 ;
  assign n66 = n62 & ~n65 ;
  assign n67 = n66 ^ n64 ;
  assign n68 = ~n46 & n67 ;
  assign n69 = n68 ^ n61 ;
  assign n70 = n69 ^ n47 ;
  assign n71 = n70 ^ n54 ;
  assign n72 = n45 & ~n71 ;
  assign n73 = n28 & n72 ;
  assign n74 = ~x3 & ~n73 ;
  assign n75 = ~x6 & ~x7 ;
  assign n76 = ~x5 & n47 ;
  assign n78 = n76 ^ x2 ;
  assign n77 = n76 ^ n10 ;
  assign n79 = n78 ^ n77 ;
  assign n80 = n79 ^ x4 ;
  assign n81 = n78 ^ x8 ;
  assign n82 = n78 ^ n76 ;
  assign n83 = n82 ^ n81 ;
  assign n84 = n81 & n83 ;
  assign n85 = n84 ^ n78 ;
  assign n86 = n85 ^ n81 ;
  assign n87 = ~n80 & ~n86 ;
  assign n88 = n87 ^ n84 ;
  assign n89 = n88 ^ n81 ;
  assign n90 = x4 & n89 ;
  assign n91 = n90 ^ n76 ;
  assign n92 = n75 & n91 ;
  assign n93 = x3 & x6 ;
  assign n94 = ~x7 & n93 ;
  assign n96 = x1 & n39 ;
  assign n97 = x5 & ~n96 ;
  assign n95 = x2 ^ x1 ;
  assign n98 = n97 ^ n95 ;
  assign n99 = n94 & ~n98 ;
  assign n100 = n99 ^ n94 ;
  assign n101 = ~x5 & x8 ;
  assign n102 = n101 ^ n99 ;
  assign n103 = n95 & ~n102 ;
  assign n104 = n103 ^ n95 ;
  assign n105 = n104 ^ n97 ;
  assign n106 = n100 & ~n105 ;
  assign n107 = ~n92 & ~n106 ;
  assign n108 = n19 & n49 ;
  assign n109 = x2 & x4 ;
  assign n110 = n23 & n109 ;
  assign n111 = n46 ^ x1 ;
  assign n112 = ~x8 & n111 ;
  assign n113 = n112 ^ x1 ;
  assign n114 = ~x4 & ~n113 ;
  assign n115 = ~n110 & ~n114 ;
  assign n116 = ~n108 & n115 ;
  assign n117 = n93 & ~n116 ;
  assign n118 = n15 & n75 ;
  assign n119 = n29 & n48 ;
  assign n120 = ~n33 & n119 ;
  assign n121 = ~n118 & ~n120 ;
  assign n122 = x5 ^ x2 ;
  assign n123 = n122 ^ x4 ;
  assign n124 = n123 ^ n122 ;
  assign n125 = n124 ^ x7 ;
  assign n126 = x6 ^ x2 ;
  assign n127 = ~x6 & ~n126 ;
  assign n128 = n127 ^ n122 ;
  assign n129 = n128 ^ x6 ;
  assign n130 = ~n125 & ~n129 ;
  assign n131 = n130 ^ n127 ;
  assign n132 = n131 ^ x6 ;
  assign n133 = x7 & ~n132 ;
  assign n134 = n133 ^ x8 ;
  assign n135 = n134 ^ n133 ;
  assign n136 = ~x1 & ~x4 ;
  assign n137 = x3 & ~n136 ;
  assign n138 = n33 ^ x2 ;
  assign n139 = n33 ^ x6 ;
  assign n140 = n139 ^ n138 ;
  assign n141 = n10 ^ x7 ;
  assign n142 = ~x6 & ~n141 ;
  assign n143 = n142 ^ n10 ;
  assign n144 = n140 & n143 ;
  assign n145 = n144 ^ n142 ;
  assign n146 = n145 ^ n10 ;
  assign n147 = n146 ^ x6 ;
  assign n148 = n138 & ~n147 ;
  assign n149 = ~n51 & ~n148 ;
  assign n150 = n137 & ~n149 ;
  assign n151 = n150 ^ n133 ;
  assign n152 = n135 & n151 ;
  assign n153 = n152 ^ n133 ;
  assign n154 = n121 & ~n153 ;
  assign n155 = ~n117 & n154 ;
  assign n156 = n155 ^ x0 ;
  assign n157 = n156 ^ n155 ;
  assign n158 = x5 ^ x1 ;
  assign n159 = ~x2 & ~x4 ;
  assign n160 = ~n11 & ~n159 ;
  assign n161 = n160 ^ x5 ;
  assign n162 = n161 ^ n160 ;
  assign n163 = n162 ^ n158 ;
  assign n164 = ~n18 & ~n39 ;
  assign n165 = n164 ^ n109 ;
  assign n166 = ~n109 & ~n165 ;
  assign n167 = n166 ^ n160 ;
  assign n168 = n167 ^ n109 ;
  assign n169 = n163 & n168 ;
  assign n170 = n169 ^ n166 ;
  assign n171 = n170 ^ n109 ;
  assign n172 = n158 & ~n171 ;
  assign n173 = ~x7 & n172 ;
  assign n174 = n41 & n93 ;
  assign n175 = ~x2 & ~x6 ;
  assign n176 = ~n33 & n175 ;
  assign n177 = ~n174 & ~n176 ;
  assign n178 = x3 & x7 ;
  assign n179 = n164 & ~n178 ;
  assign n180 = x6 & x7 ;
  assign n181 = ~x3 & ~x6 ;
  assign n182 = x2 & ~n181 ;
  assign n183 = ~n180 & ~n182 ;
  assign n184 = n33 & ~n183 ;
  assign n185 = ~n179 & n184 ;
  assign n186 = n177 & ~n185 ;
  assign n187 = ~n173 & n186 ;
  assign n188 = n187 ^ n155 ;
  assign n189 = ~n157 & n188 ;
  assign n190 = n189 ^ n155 ;
  assign n191 = n107 & n190 ;
  assign n192 = ~n74 & n191 ;
  assign y0 = ~n192 ;
endmodule
