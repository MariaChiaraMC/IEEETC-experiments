module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 ;
  assign n105 = x11 ^ x10 ;
  assign n91 = ~x10 & ~x11 ;
  assign n20 = ~x2 & ~x3 ;
  assign n81 = ~x4 & ~x9 ;
  assign n82 = n20 & n81 ;
  assign n83 = ~x10 & ~n82 ;
  assign n84 = x1 ^ x0 ;
  assign n85 = ~x1 & x8 ;
  assign n86 = ~n84 & n85 ;
  assign n87 = n86 ^ n84 ;
  assign n88 = ~n83 & ~n87 ;
  assign n89 = ~x11 & ~n88 ;
  assign n16 = x9 ^ x4 ;
  assign n17 = ~x1 & n16 ;
  assign n21 = x6 & x7 ;
  assign n22 = n20 & ~n21 ;
  assign n18 = ~x3 & ~x5 ;
  assign n19 = ~x6 & n18 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n22 ^ x9 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n25 ^ n17 ;
  assign n27 = n23 & ~n26 ;
  assign n28 = n27 ^ n19 ;
  assign n29 = n17 & n28 ;
  assign n30 = n29 ^ x9 ;
  assign n39 = x3 ^ x2 ;
  assign n40 = n39 ^ x4 ;
  assign n41 = n40 ^ x5 ;
  assign n46 = n41 ^ n40 ;
  assign n47 = n46 ^ x3 ;
  assign n48 = n47 ^ x3 ;
  assign n49 = n40 ^ x4 ;
  assign n50 = n49 ^ n40 ;
  assign n51 = n50 ^ x3 ;
  assign n52 = ~n48 & ~n51 ;
  assign n42 = n40 ^ x6 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = n43 ^ x3 ;
  assign n45 = ~n41 & ~n44 ;
  assign n53 = n52 ^ n45 ;
  assign n54 = n53 ^ n41 ;
  assign n55 = n45 ^ x3 ;
  assign n56 = n55 ^ n47 ;
  assign n57 = x3 & ~n56 ;
  assign n58 = n57 ^ n45 ;
  assign n59 = ~n54 & n58 ;
  assign n60 = n59 ^ n52 ;
  assign n61 = n60 ^ n57 ;
  assign n62 = n61 ^ n41 ;
  assign n63 = n62 ^ x3 ;
  assign n64 = n63 ^ n47 ;
  assign n65 = n64 ^ x2 ;
  assign n66 = x1 & ~n65 ;
  assign n67 = x6 & ~x7 ;
  assign n68 = ~x2 & n67 ;
  assign n69 = n18 & n68 ;
  assign n70 = ~n66 & ~n69 ;
  assign n31 = x5 & x6 ;
  assign n32 = x5 & x9 ;
  assign n33 = ~x1 & ~n32 ;
  assign n34 = ~n31 & n33 ;
  assign n35 = x4 & ~x6 ;
  assign n36 = x2 & n18 ;
  assign n37 = ~n35 & n36 ;
  assign n38 = ~n34 & ~n37 ;
  assign n71 = n70 ^ n38 ;
  assign n72 = n71 ^ n38 ;
  assign n73 = ~x1 & ~n39 ;
  assign n74 = n73 ^ n38 ;
  assign n75 = n74 ^ n38 ;
  assign n76 = n72 & ~n75 ;
  assign n77 = n76 ^ n38 ;
  assign n78 = x0 & n77 ;
  assign n79 = n78 ^ n38 ;
  assign n80 = ~n30 & n79 ;
  assign n90 = n89 ^ n80 ;
  assign n92 = n91 ^ n90 ;
  assign n93 = n92 ^ n90 ;
  assign n94 = n93 ^ x13 ;
  assign n95 = n90 ^ n80 ;
  assign n96 = n95 ^ x14 ;
  assign n97 = ~x14 & n96 ;
  assign n98 = n97 ^ n90 ;
  assign n99 = n98 ^ x14 ;
  assign n100 = n94 & ~n99 ;
  assign n101 = n100 ^ n97 ;
  assign n102 = n101 ^ x14 ;
  assign n103 = ~x13 & ~n102 ;
  assign n104 = n103 ^ n89 ;
  assign n106 = n105 ^ n104 ;
  assign n108 = n106 ^ x13 ;
  assign n109 = n108 ^ n106 ;
  assign n107 = n106 ^ n104 ;
  assign n110 = n109 ^ n107 ;
  assign n111 = n106 ^ x10 ;
  assign n112 = n111 ^ n106 ;
  assign n113 = n112 ^ n109 ;
  assign n114 = ~n109 & ~n113 ;
  assign n115 = n114 ^ n109 ;
  assign n116 = ~n110 & ~n115 ;
  assign n117 = n116 ^ n114 ;
  assign n118 = n117 ^ n106 ;
  assign n119 = n118 ^ n109 ;
  assign n120 = x12 & n119 ;
  assign n121 = n120 ^ n104 ;
  assign y0 = ~n121 ;
endmodule
