module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 ;
  assign n20 = ~x0 & ~x15 ;
  assign n21 = x6 & ~x8 ;
  assign n22 = x14 & x18 ;
  assign n23 = ~n21 & n22 ;
  assign n24 = x16 & n23 ;
  assign n25 = x16 & ~x18 ;
  assign n26 = x9 & ~x14 ;
  assign n27 = ~x6 & x8 ;
  assign n28 = n26 & n27 ;
  assign n29 = n25 & n28 ;
  assign n30 = x4 & n29 ;
  assign n31 = ~n22 & ~n30 ;
  assign n32 = x7 & ~n31 ;
  assign n33 = x12 & x13 ;
  assign n34 = x11 & n33 ;
  assign n35 = ~x11 & ~x12 ;
  assign n36 = x1 & ~n35 ;
  assign n37 = x3 & ~x5 ;
  assign n38 = ~x10 & ~x18 ;
  assign n39 = n37 & n38 ;
  assign n40 = n36 & n39 ;
  assign n41 = ~x14 & ~x16 ;
  assign n42 = n40 & n41 ;
  assign n43 = ~n34 & n42 ;
  assign n44 = ~n32 & ~n43 ;
  assign n45 = ~x6 & ~x8 ;
  assign n46 = ~x16 & x18 ;
  assign n47 = ~n45 & n46 ;
  assign n48 = ~n25 & ~n47 ;
  assign n49 = x14 & ~n48 ;
  assign n50 = n49 ^ x7 ;
  assign n51 = n21 & n25 ;
  assign n56 = n51 ^ x9 ;
  assign n67 = n56 ^ n51 ;
  assign n52 = ~x6 & x16 ;
  assign n53 = x6 & ~x16 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = n54 ^ n51 ;
  assign n57 = n56 ^ n55 ;
  assign n58 = n57 ^ n56 ;
  assign n59 = n58 ^ n51 ;
  assign n60 = x18 & ~n26 ;
  assign n61 = ~x8 & n60 ;
  assign n62 = n61 ^ x18 ;
  assign n63 = n62 ^ n57 ;
  assign n64 = n63 ^ n57 ;
  assign n65 = n64 ^ n59 ;
  assign n66 = n59 & n65 ;
  assign n68 = n67 ^ n66 ;
  assign n69 = n68 ^ n59 ;
  assign n70 = n51 ^ x8 ;
  assign n71 = n66 ^ n59 ;
  assign n72 = n70 & n71 ;
  assign n73 = n72 ^ n51 ;
  assign n74 = ~n69 & ~n73 ;
  assign n75 = n74 ^ n51 ;
  assign n76 = n75 ^ x9 ;
  assign n77 = n76 ^ n51 ;
  assign n78 = x4 & ~n77 ;
  assign n79 = n78 ^ n49 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = n27 & ~n46 ;
  assign n82 = n81 ^ n78 ;
  assign n83 = n80 & n82 ;
  assign n84 = n83 ^ n78 ;
  assign n85 = ~n50 & ~n84 ;
  assign n86 = n85 ^ x7 ;
  assign n87 = n44 & n86 ;
  assign n88 = n87 ^ x17 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = x16 ^ x6 ;
  assign n91 = n90 ^ x18 ;
  assign n92 = x18 ^ x16 ;
  assign n93 = n92 ^ x16 ;
  assign n94 = ~x7 & x8 ;
  assign n95 = n94 ^ x16 ;
  assign n96 = ~n93 & ~n95 ;
  assign n97 = n96 ^ x16 ;
  assign n98 = ~n91 & ~n97 ;
  assign n99 = n98 ^ x18 ;
  assign n100 = x14 & ~n99 ;
  assign n101 = x7 & ~x8 ;
  assign n102 = n22 & ~n101 ;
  assign n103 = x9 ^ x8 ;
  assign n104 = n103 ^ x18 ;
  assign n105 = x9 ^ x7 ;
  assign n106 = n105 ^ x7 ;
  assign n107 = n106 ^ n104 ;
  assign n108 = x18 ^ x7 ;
  assign n109 = n108 ^ x14 ;
  assign n110 = ~x14 & n109 ;
  assign n111 = n110 ^ x7 ;
  assign n112 = n111 ^ x14 ;
  assign n113 = ~n107 & ~n112 ;
  assign n114 = n113 ^ n110 ;
  assign n115 = n114 ^ x14 ;
  assign n116 = ~n104 & ~n115 ;
  assign n117 = n54 & n116 ;
  assign n118 = x4 & n117 ;
  assign n119 = ~n102 & ~n118 ;
  assign n120 = ~n100 & n119 ;
  assign n121 = n120 ^ n87 ;
  assign n122 = n89 & n121 ;
  assign n123 = n122 ^ n87 ;
  assign n124 = ~n24 & n123 ;
  assign n125 = n20 & ~n124 ;
  assign y0 = n125 ;
endmodule
