module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 ;
  assign n13 = x7 & x8 ;
  assign n107 = ~x10 & n13 ;
  assign n14 = x0 & x3 ;
  assign n15 = x10 & n14 ;
  assign n16 = ~x1 & n15 ;
  assign n17 = n13 & n16 ;
  assign n18 = x5 & ~x6 ;
  assign n19 = x0 & x5 ;
  assign n20 = ~n18 & ~n19 ;
  assign n21 = ~n14 & ~n20 ;
  assign n22 = ~x10 & ~n21 ;
  assign n23 = ~x1 & n22 ;
  assign n24 = x8 ^ x1 ;
  assign n25 = x8 ^ x0 ;
  assign n26 = n25 ^ x0 ;
  assign n27 = n20 ^ x0 ;
  assign n28 = n26 & n27 ;
  assign n29 = n28 ^ x0 ;
  assign n30 = n24 & ~n29 ;
  assign n31 = n30 ^ x1 ;
  assign n32 = ~n23 & ~n31 ;
  assign n33 = x1 & ~x3 ;
  assign n34 = x0 & ~x4 ;
  assign n35 = n33 & n34 ;
  assign n36 = x10 & n35 ;
  assign n37 = ~n15 & ~n36 ;
  assign n38 = ~n32 & n37 ;
  assign n39 = ~x3 & x10 ;
  assign n40 = x4 & n39 ;
  assign n41 = ~x7 & ~n40 ;
  assign n42 = ~n38 & n41 ;
  assign n43 = ~x10 & ~x11 ;
  assign n44 = x4 & n20 ;
  assign n45 = n44 ^ n19 ;
  assign n46 = ~x7 & ~n45 ;
  assign n47 = n39 & ~n46 ;
  assign n48 = n14 ^ x10 ;
  assign n49 = n48 ^ n14 ;
  assign n50 = ~x7 & ~n18 ;
  assign n51 = ~x0 & ~n50 ;
  assign n52 = n51 ^ n14 ;
  assign n53 = n49 & ~n52 ;
  assign n54 = n53 ^ n14 ;
  assign n55 = ~x1 & n54 ;
  assign n56 = ~n47 & n55 ;
  assign n57 = x8 & ~n56 ;
  assign n58 = ~n43 & n57 ;
  assign n59 = ~n42 & ~n58 ;
  assign n60 = n59 ^ x2 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = n61 ^ n17 ;
  assign n63 = ~x6 & ~x8 ;
  assign n64 = ~x5 & n63 ;
  assign n65 = ~x3 & n64 ;
  assign n66 = x0 & ~x1 ;
  assign n67 = ~n39 & n66 ;
  assign n68 = n67 ^ x10 ;
  assign n69 = n67 ^ x7 ;
  assign n70 = n69 ^ x7 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = x11 ^ x8 ;
  assign n73 = ~x11 & ~n72 ;
  assign n74 = n73 ^ x7 ;
  assign n75 = n74 ^ x11 ;
  assign n76 = n71 & n75 ;
  assign n77 = n76 ^ n73 ;
  assign n78 = n77 ^ x11 ;
  assign n79 = ~n68 & ~n78 ;
  assign n80 = n79 ^ n67 ;
  assign n81 = ~n65 & n80 ;
  assign n82 = x6 ^ x4 ;
  assign n83 = x5 & ~n82 ;
  assign n84 = n83 ^ x4 ;
  assign n85 = ~x7 & ~x10 ;
  assign n86 = x1 ^ x0 ;
  assign n87 = n86 ^ n85 ;
  assign n88 = x5 ^ x3 ;
  assign n89 = ~x1 & ~n88 ;
  assign n90 = n89 ^ x3 ;
  assign n91 = ~n87 & n90 ;
  assign n92 = n91 ^ n89 ;
  assign n93 = n92 ^ x3 ;
  assign n94 = n93 ^ x1 ;
  assign n95 = n85 & ~n94 ;
  assign n96 = n84 & n95 ;
  assign n97 = ~x8 & ~n96 ;
  assign n98 = n97 ^ n81 ;
  assign n99 = ~n81 & n98 ;
  assign n100 = n99 ^ n59 ;
  assign n101 = n100 ^ n81 ;
  assign n102 = ~n62 & n101 ;
  assign n103 = n102 ^ n99 ;
  assign n104 = n103 ^ n81 ;
  assign n105 = ~n17 & ~n104 ;
  assign n106 = n105 ^ n17 ;
  assign n108 = n107 ^ n106 ;
  assign n109 = x9 & n108 ;
  assign n110 = n109 ^ n106 ;
  assign y0 = n110 ;
endmodule
