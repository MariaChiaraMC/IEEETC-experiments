module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 ;
  assign n8 = ~x2 & ~x3 ;
  assign n9 = x1 & ~x6 ;
  assign n10 = n8 & ~n9 ;
  assign n11 = ~x0 & ~n10 ;
  assign n12 = x3 ^ x2 ;
  assign n13 = x5 ^ x3 ;
  assign n14 = n12 & n13 ;
  assign n15 = n14 ^ x3 ;
  assign n16 = ~x4 & x6 ;
  assign n17 = ~x3 & n16 ;
  assign n18 = n17 ^ x1 ;
  assign n19 = ~n15 & n18 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = x1 & n20 ;
  assign n22 = n21 ^ x1 ;
  assign n23 = n11 & ~n22 ;
  assign y0 = n23 ;
endmodule
