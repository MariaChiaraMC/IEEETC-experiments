module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 ;
  output y0 ;
  wire n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 ;
  assign n14 = x4 & ~x9 ;
  assign n15 = ~x8 & ~n14 ;
  assign n16 = x3 & ~x7 ;
  assign n17 = x2 & ~x6 ;
  assign n18 = x1 & ~x5 ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = ~n16 & n19 ;
  assign n21 = ~x12 & n20 ;
  assign n22 = ~x6 & ~x7 ;
  assign n23 = ~x5 & ~x11 ;
  assign n24 = n22 & n23 ;
  assign n25 = ~x2 & ~x3 ;
  assign n26 = ~x1 & n25 ;
  assign n27 = ~n24 & ~n26 ;
  assign n28 = ~n21 & n27 ;
  assign n29 = ~n15 & ~n28 ;
  assign n30 = ~x1 & ~x6 ;
  assign n31 = x3 & x7 ;
  assign n32 = ~x11 & ~n31 ;
  assign n33 = n30 & n32 ;
  assign n34 = x2 & x6 ;
  assign n35 = n23 & ~n34 ;
  assign n36 = ~n31 & n35 ;
  assign n37 = x6 & x7 ;
  assign n38 = x11 & ~n37 ;
  assign n39 = ~x5 & x11 ;
  assign n40 = ~x12 & ~n39 ;
  assign n41 = ~n38 & n40 ;
  assign n42 = ~n36 & ~n41 ;
  assign n43 = ~x2 & ~x7 ;
  assign n44 = ~x11 & n43 ;
  assign n45 = ~n25 & ~n44 ;
  assign n46 = ~x1 & ~n45 ;
  assign n47 = n42 & ~n46 ;
  assign n48 = ~n33 & n47 ;
  assign n49 = ~x10 & ~n48 ;
  assign n50 = n49 ^ x11 ;
  assign n51 = n50 ^ x4 ;
  assign n66 = n51 ^ n50 ;
  assign n53 = ~x2 & ~x5 ;
  assign n54 = ~n30 & ~n53 ;
  assign n55 = ~n31 & ~n54 ;
  assign n56 = ~x1 & n43 ;
  assign n57 = ~x3 & ~x6 ;
  assign n58 = ~x5 & n57 ;
  assign n59 = ~n56 & ~n58 ;
  assign n60 = ~n55 & n59 ;
  assign n61 = x8 & ~n60 ;
  assign n52 = n51 ^ n49 ;
  assign n62 = n61 ^ n52 ;
  assign n63 = n61 ^ n51 ;
  assign n64 = n63 ^ n50 ;
  assign n65 = n62 & n64 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = ~x9 & ~x12 ;
  assign n69 = n68 ^ n51 ;
  assign n70 = ~n66 & n69 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = ~n67 & n71 ;
  assign n73 = n72 ^ n65 ;
  assign n74 = n73 ^ n51 ;
  assign n75 = n74 ^ x11 ;
  assign n76 = n75 ^ n50 ;
  assign n77 = ~n29 & ~n76 ;
  assign n78 = ~x0 & ~n77 ;
  assign n79 = ~x4 & x8 ;
  assign n80 = n36 & n79 ;
  assign n81 = x10 ^ x9 ;
  assign n82 = ~x6 & n81 ;
  assign n83 = n82 ^ x9 ;
  assign n84 = ~n45 & ~n83 ;
  assign n85 = ~n80 & ~n84 ;
  assign n86 = ~x5 & ~x10 ;
  assign n87 = x5 & ~x9 ;
  assign n88 = ~n86 & ~n87 ;
  assign n89 = n26 & ~n88 ;
  assign n90 = ~x7 & n81 ;
  assign n91 = n90 ^ x9 ;
  assign n92 = ~x3 & ~n91 ;
  assign n93 = ~n89 & ~n92 ;
  assign n94 = n85 & n93 ;
  assign n98 = ~n43 & ~n57 ;
  assign n97 = ~n22 & ~n25 ;
  assign n99 = n98 ^ n97 ;
  assign n108 = n99 ^ n98 ;
  assign n100 = n98 ^ n79 ;
  assign n101 = n100 ^ n99 ;
  assign n102 = n101 ^ n99 ;
  assign n103 = n102 ^ n98 ;
  assign n104 = n101 ^ n86 ;
  assign n105 = n104 ^ n101 ;
  assign n106 = n105 ^ n103 ;
  assign n107 = ~n103 & n106 ;
  assign n109 = n108 ^ n107 ;
  assign n110 = n109 ^ n103 ;
  assign n111 = n98 ^ n87 ;
  assign n112 = n107 ^ n103 ;
  assign n113 = n111 & ~n112 ;
  assign n114 = n113 ^ n98 ;
  assign n115 = ~n110 & ~n114 ;
  assign n116 = n115 ^ n98 ;
  assign n117 = n116 ^ n97 ;
  assign n118 = n117 ^ n98 ;
  assign n119 = ~x11 & ~n118 ;
  assign n95 = x12 ^ x1 ;
  assign n120 = n119 ^ n95 ;
  assign n96 = n95 ^ x12 ;
  assign n121 = n120 ^ n96 ;
  assign n122 = n121 ^ n120 ;
  assign n123 = n122 ^ n95 ;
  assign n124 = x4 & n20 ;
  assign n125 = x11 & ~n124 ;
  assign n126 = x8 & ~n125 ;
  assign n127 = n126 ^ n120 ;
  assign n128 = n127 ^ n122 ;
  assign n129 = n128 ^ n123 ;
  assign n130 = n123 & ~n129 ;
  assign n131 = n130 ^ n126 ;
  assign n132 = ~x2 & x7 ;
  assign n133 = ~n83 & n132 ;
  assign n134 = n133 ^ n120 ;
  assign n135 = n134 ^ n122 ;
  assign n136 = n134 ^ n126 ;
  assign n137 = ~n135 & ~n136 ;
  assign n138 = n137 ^ n133 ;
  assign n139 = n138 ^ n123 ;
  assign n140 = ~n38 & ~n88 ;
  assign n141 = ~x3 & x6 ;
  assign n142 = ~n132 & ~n141 ;
  assign n143 = n87 & ~n142 ;
  assign n144 = ~n140 & ~n143 ;
  assign n145 = n133 ^ n123 ;
  assign n146 = n144 & n145 ;
  assign n147 = n146 ^ n144 ;
  assign n148 = n147 ^ n126 ;
  assign n149 = n148 ^ n122 ;
  assign n150 = n149 ^ n123 ;
  assign n151 = n139 & n150 ;
  assign n152 = n151 ^ n122 ;
  assign n153 = n152 ^ n123 ;
  assign n154 = n131 & n153 ;
  assign n155 = n154 ^ n151 ;
  assign n156 = n155 ^ n122 ;
  assign n157 = n156 ^ n123 ;
  assign n158 = n157 ^ x12 ;
  assign n159 = n94 & n158 ;
  assign n160 = ~n78 & n159 ;
  assign y0 = ~n160 ;
endmodule
