module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 ;
  assign n75 = x7 ^ x4 ;
  assign n16 = ~x3 & ~x5 ;
  assign n17 = x1 & ~n16 ;
  assign n76 = n17 ^ x7 ;
  assign n77 = n76 ^ n17 ;
  assign n78 = ~x1 & ~x3 ;
  assign n79 = n78 ^ n17 ;
  assign n80 = ~n77 & n79 ;
  assign n81 = n80 ^ n17 ;
  assign n82 = n75 & n81 ;
  assign n83 = x6 & n82 ;
  assign n84 = ~x1 & x3 ;
  assign n85 = x5 & ~x7 ;
  assign n86 = n84 & n85 ;
  assign n87 = x4 & n86 ;
  assign n88 = ~n83 & ~n87 ;
  assign n89 = x2 & ~n88 ;
  assign n90 = ~x1 & x2 ;
  assign n91 = x6 ^ x4 ;
  assign n92 = x4 & x7 ;
  assign n93 = n92 ^ x3 ;
  assign n94 = ~n91 & n93 ;
  assign n95 = ~x1 & n94 ;
  assign n96 = ~n90 & ~n95 ;
  assign n97 = x3 & ~x7 ;
  assign n98 = ~x4 & x6 ;
  assign n99 = n97 & n98 ;
  assign n25 = ~x3 & x7 ;
  assign n100 = ~x6 & n25 ;
  assign n101 = x2 & ~n100 ;
  assign n102 = ~n99 & n101 ;
  assign n103 = ~n96 & ~n102 ;
  assign n105 = ~x7 & n98 ;
  assign n104 = x1 & ~x2 ;
  assign n106 = n105 ^ n104 ;
  assign n107 = x3 & n92 ;
  assign n108 = n107 ^ n104 ;
  assign n109 = n108 ^ n107 ;
  assign n110 = ~x3 & ~n90 ;
  assign n111 = n110 ^ n107 ;
  assign n112 = ~n109 & ~n111 ;
  assign n113 = n112 ^ n107 ;
  assign n114 = n106 & n113 ;
  assign n115 = n114 ^ n105 ;
  assign n116 = ~n103 & ~n115 ;
  assign n117 = n116 ^ x2 ;
  assign n118 = n117 ^ n116 ;
  assign n18 = ~x4 & ~x6 ;
  assign n26 = n18 & n25 ;
  assign n27 = x1 & n26 ;
  assign n119 = ~x4 & x7 ;
  assign n120 = n84 & n119 ;
  assign n121 = ~n25 & ~n97 ;
  assign n122 = x4 & ~n121 ;
  assign n123 = x1 & n122 ;
  assign n124 = ~n120 & ~n123 ;
  assign n125 = x6 & ~n124 ;
  assign n126 = ~n27 & ~n125 ;
  assign n127 = n126 ^ n116 ;
  assign n128 = n127 ^ n116 ;
  assign n129 = ~n118 & ~n128 ;
  assign n130 = n129 ^ n116 ;
  assign n131 = x5 & ~n130 ;
  assign n132 = n131 ^ n116 ;
  assign n133 = ~n89 & n132 ;
  assign n9 = ~x2 & x5 ;
  assign n10 = ~x1 & ~x6 ;
  assign n11 = n9 & ~n10 ;
  assign n12 = x4 ^ x1 ;
  assign n13 = ~x3 & n12 ;
  assign n14 = n13 ^ x1 ;
  assign n15 = n11 & ~n14 ;
  assign n19 = x3 & x5 ;
  assign n20 = x2 & ~n19 ;
  assign n21 = n18 & n20 ;
  assign n22 = ~n17 & n21 ;
  assign n23 = ~n15 & ~n22 ;
  assign n24 = ~x7 & ~n23 ;
  assign n28 = x2 & x5 ;
  assign n29 = ~x2 & ~x5 ;
  assign n30 = ~n28 & ~n29 ;
  assign n31 = n27 & ~n30 ;
  assign n32 = x7 ^ x3 ;
  assign n33 = x7 ^ x5 ;
  assign n34 = x5 ^ x1 ;
  assign n35 = n34 ^ x5 ;
  assign n36 = ~n33 & ~n35 ;
  assign n37 = n36 ^ x5 ;
  assign n38 = ~n32 & ~n37 ;
  assign n39 = n38 ^ x5 ;
  assign n40 = x2 & ~n39 ;
  assign n41 = x6 & ~n40 ;
  assign n42 = ~n19 & ~n28 ;
  assign n43 = n42 ^ n17 ;
  assign n44 = n43 ^ n17 ;
  assign n45 = x2 & x3 ;
  assign n46 = ~x1 & ~n45 ;
  assign n47 = n46 ^ n17 ;
  assign n48 = ~n44 & n47 ;
  assign n49 = n48 ^ n17 ;
  assign n50 = x7 & n49 ;
  assign n51 = x5 ^ x2 ;
  assign n52 = n32 ^ x7 ;
  assign n53 = n33 ^ x7 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = n54 ^ x7 ;
  assign n56 = n51 & ~n55 ;
  assign n57 = n56 ^ x7 ;
  assign n58 = n57 ^ x1 ;
  assign n59 = n58 ^ n57 ;
  assign n60 = n59 ^ x6 ;
  assign n61 = n29 ^ x3 ;
  assign n62 = n29 & ~n61 ;
  assign n63 = n62 ^ n57 ;
  assign n64 = n63 ^ n29 ;
  assign n65 = n60 & ~n64 ;
  assign n66 = n65 ^ n62 ;
  assign n67 = n66 ^ n29 ;
  assign n68 = ~x6 & n67 ;
  assign n69 = n68 ^ x6 ;
  assign n70 = ~n50 & ~n69 ;
  assign n71 = x4 & ~n70 ;
  assign n72 = ~n41 & n71 ;
  assign n73 = ~n31 & ~n72 ;
  assign n74 = ~n24 & n73 ;
  assign n134 = n133 ^ n74 ;
  assign n135 = ~x0 & n134 ;
  assign n136 = n135 ^ n133 ;
  assign y0 = ~n136 ;
endmodule
