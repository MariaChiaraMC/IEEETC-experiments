module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 ;
  assign n8 = ~x0 & ~x1 ;
  assign n9 = ~x3 & ~n8 ;
  assign n10 = x5 & x6 ;
  assign n11 = ~x1 & x3 ;
  assign n12 = n10 & ~n11 ;
  assign n13 = ~n9 & n12 ;
  assign n14 = x2 & n13 ;
  assign n15 = x0 & x1 ;
  assign n16 = ~x2 & ~n15 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = n17 ^ n8 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = n17 ^ n16 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n19 & n21 ;
  assign n23 = n22 ^ n17 ;
  assign n24 = ~x6 & n23 ;
  assign n25 = n24 ^ n17 ;
  assign n26 = x3 & n25 ;
  assign n27 = ~x3 & n10 ;
  assign n28 = n27 ^ x2 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = ~x3 & ~x6 ;
  assign n31 = x3 ^ x1 ;
  assign n32 = n31 ^ x5 ;
  assign n33 = n32 ^ n31 ;
  assign n36 = x1 ^ x0 ;
  assign n37 = n36 ^ n31 ;
  assign n38 = ~n31 & n37 ;
  assign n34 = x1 & x6 ;
  assign n41 = n38 ^ n34 ;
  assign n35 = n34 ^ n33 ;
  assign n39 = n38 ^ n31 ;
  assign n40 = n35 & ~n39 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = n33 & n42 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = n44 ^ n40 ;
  assign n46 = n45 ^ x1 ;
  assign n47 = ~n30 & ~n46 ;
  assign n48 = n47 ^ n27 ;
  assign n49 = n29 & ~n48 ;
  assign n50 = n49 ^ n27 ;
  assign n51 = ~n26 & ~n50 ;
  assign n52 = n51 ^ x4 ;
  assign n53 = n52 ^ n51 ;
  assign n56 = x2 ^ x0 ;
  assign n57 = n56 ^ x0 ;
  assign n58 = n57 ^ x6 ;
  assign n62 = n58 ^ n56 ;
  assign n54 = x6 ^ x3 ;
  assign n55 = n54 ^ x3 ;
  assign n59 = n58 ^ x3 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = n55 & ~n60 ;
  assign n63 = n62 ^ n61 ;
  assign n64 = n63 ^ x5 ;
  assign n65 = n56 ^ x1 ;
  assign n66 = n62 ^ x5 ;
  assign n67 = ~n65 & ~n66 ;
  assign n68 = n67 ^ n61 ;
  assign n69 = n68 ^ n56 ;
  assign n70 = n69 ^ n65 ;
  assign n71 = n70 ^ n62 ;
  assign n72 = x5 & n71 ;
  assign n73 = ~n64 & n72 ;
  assign n74 = x5 ^ x2 ;
  assign n75 = n74 ^ n11 ;
  assign n86 = x1 & ~x3 ;
  assign n87 = x6 & ~n86 ;
  assign n76 = n30 ^ x3 ;
  assign n77 = n76 ^ x0 ;
  assign n78 = x2 ^ x1 ;
  assign n79 = x3 & n78 ;
  assign n80 = n79 ^ x1 ;
  assign n81 = ~n77 & ~n80 ;
  assign n82 = n81 ^ n79 ;
  assign n83 = n82 ^ x1 ;
  assign n84 = n83 ^ x3 ;
  assign n85 = ~x0 & ~n84 ;
  assign n88 = n87 ^ n85 ;
  assign n89 = n85 ^ x5 ;
  assign n90 = n89 ^ n85 ;
  assign n91 = n88 & n90 ;
  assign n92 = n91 ^ n85 ;
  assign n93 = n75 & ~n92 ;
  assign n94 = n93 ^ x5 ;
  assign n95 = ~n73 & n94 ;
  assign n96 = n95 ^ n51 ;
  assign n97 = ~n53 & n96 ;
  assign n98 = n97 ^ n51 ;
  assign n99 = ~n14 & n98 ;
  assign y0 = ~n99 ;
endmodule
