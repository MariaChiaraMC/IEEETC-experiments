module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 ;
  assign n9 = ~x6 & ~x7 ;
  assign n10 = x2 & x4 ;
  assign n11 = ~x5 & n10 ;
  assign n12 = n9 & n11 ;
  assign n13 = x1 & ~x6 ;
  assign n14 = ~x4 & x5 ;
  assign n15 = x1 & ~n14 ;
  assign n16 = ~n13 & ~n15 ;
  assign n17 = ~n12 & ~n16 ;
  assign n18 = x6 & x7 ;
  assign n19 = ~x5 & ~n18 ;
  assign n20 = x4 & ~n19 ;
  assign n21 = ~x1 & ~n20 ;
  assign n22 = x5 & ~n9 ;
  assign n23 = ~x1 & ~x2 ;
  assign n24 = ~n22 & n23 ;
  assign n25 = ~x3 & ~n24 ;
  assign n26 = ~n21 & n25 ;
  assign n27 = ~n17 & n26 ;
  assign n28 = x3 & ~x4 ;
  assign n29 = n19 & n28 ;
  assign n30 = n23 & n29 ;
  assign n31 = ~n27 & ~n30 ;
  assign n32 = x0 & ~n31 ;
  assign n39 = x6 ^ x1 ;
  assign n33 = x6 ^ x0 ;
  assign n34 = n33 ^ x1 ;
  assign n35 = x7 ^ x0 ;
  assign n36 = n35 ^ x0 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = ~n34 & n37 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = n40 ^ n34 ;
  assign n42 = x2 ^ x1 ;
  assign n43 = n42 ^ x1 ;
  assign n44 = n38 ^ n34 ;
  assign n45 = n43 & ~n44 ;
  assign n46 = n45 ^ x1 ;
  assign n47 = ~n41 & n46 ;
  assign n48 = n47 ^ x1 ;
  assign n49 = n48 ^ x1 ;
  assign n50 = n49 ^ x5 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = n51 ^ x4 ;
  assign n53 = n9 ^ x0 ;
  assign n54 = ~n9 & n53 ;
  assign n55 = n54 ^ n49 ;
  assign n56 = n55 ^ n9 ;
  assign n57 = n52 & ~n56 ;
  assign n58 = n57 ^ n54 ;
  assign n59 = n58 ^ n9 ;
  assign n60 = ~x4 & ~n59 ;
  assign n61 = ~x3 & n60 ;
  assign n62 = ~n32 & ~n61 ;
  assign y0 = ~n62 ;
endmodule
