module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 ;
  assign n10 = ~x2 & ~x3 ;
  assign n11 = ~x1 & n10 ;
  assign n12 = x5 & ~n11 ;
  assign n13 = n12 ^ x6 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n14 ^ x7 ;
  assign n16 = ~x2 & x3 ;
  assign n17 = x5 & ~n16 ;
  assign n18 = x1 & n17 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = ~n18 & ~n19 ;
  assign n21 = n20 ^ n12 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = ~n15 & ~n22 ;
  assign n24 = n23 ^ n20 ;
  assign n25 = n24 ^ n18 ;
  assign n26 = x7 & ~n25 ;
  assign n27 = n26 ^ x7 ;
  assign y0 = ~n27 ;
endmodule
