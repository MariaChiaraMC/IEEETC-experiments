module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 ;
  assign n24 = ~x0 & ~x2 ;
  assign n25 = x4 & ~n24 ;
  assign n26 = n25 ^ x2 ;
  assign n27 = n25 ^ x5 ;
  assign n28 = n26 & n27 ;
  assign n29 = n28 ^ n25 ;
  assign n30 = x6 & n25 ;
  assign n31 = n30 ^ x3 ;
  assign n32 = n29 & n31 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = x3 & n33 ;
  assign n35 = n34 ^ x3 ;
  assign n36 = n35 ^ x3 ;
  assign n8 = x2 ^ x0 ;
  assign n9 = x3 ^ x2 ;
  assign n10 = n9 ^ x2 ;
  assign n11 = n10 ^ n8 ;
  assign n12 = x4 ^ x2 ;
  assign n13 = x5 & x6 ;
  assign n14 = n13 ^ x2 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n12 & n15 ;
  assign n17 = n16 ^ x2 ;
  assign n18 = n17 ^ n12 ;
  assign n19 = ~n11 & ~n18 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = n20 ^ n12 ;
  assign n22 = n8 & n21 ;
  assign n23 = n22 ^ x2 ;
  assign n37 = n36 ^ n23 ;
  assign n38 = n37 ^ n23 ;
  assign n39 = x0 & x2 ;
  assign n40 = n39 ^ n23 ;
  assign n41 = n40 ^ n23 ;
  assign n42 = ~n38 & ~n41 ;
  assign n43 = n42 ^ n23 ;
  assign n44 = ~x1 & n43 ;
  assign n45 = n44 ^ n23 ;
  assign y0 = ~n45 ;
endmodule
