module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 ;
  assign n34 = ~x3 & ~x4 ;
  assign n10 = x4 ^ x3 ;
  assign n9 = x5 ^ x4 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = n10 ^ x5 ;
  assign n13 = n12 ^ x6 ;
  assign n14 = n13 ^ n10 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = ~n11 & n15 ;
  assign n17 = n16 ^ n10 ;
  assign n18 = n17 ^ n11 ;
  assign n19 = n10 ^ x7 ;
  assign n20 = n19 ^ x1 ;
  assign n21 = ~x7 & ~n20 ;
  assign n22 = n21 ^ x7 ;
  assign n23 = n22 ^ n10 ;
  assign n24 = x7 ^ x6 ;
  assign n25 = n19 & n24 ;
  assign n26 = n25 ^ x6 ;
  assign n27 = n26 ^ x1 ;
  assign n28 = n23 & n27 ;
  assign n29 = n28 ^ x1 ;
  assign n30 = n18 & ~n29 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n31 ^ x1 ;
  assign n33 = n32 ^ x1 ;
  assign n35 = n34 ^ n33 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = n33 ^ x1 ;
  assign n38 = n37 ^ n33 ;
  assign n39 = ~n36 & ~n38 ;
  assign n40 = n39 ^ n33 ;
  assign n41 = x2 & ~n40 ;
  assign n42 = n41 ^ n33 ;
  assign y0 = ~n42 ;
endmodule
