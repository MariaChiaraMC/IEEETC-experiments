module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 ;
  assign n17 = x15 ^ x14 ;
  assign n18 = ~x13 & ~n17 ;
  assign n19 = x6 & ~n18 ;
  assign n20 = x7 & ~x8 ;
  assign n21 = x5 & n20 ;
  assign n22 = x4 & n21 ;
  assign n23 = ~x14 & ~x15 ;
  assign n24 = x13 & ~n23 ;
  assign n25 = x10 ^ x9 ;
  assign n26 = ~n24 & n25 ;
  assign n27 = n22 & n26 ;
  assign n28 = n19 & n27 ;
  assign n29 = ~x9 & x10 ;
  assign n30 = ~x13 & n29 ;
  assign n31 = ~x5 & ~x7 ;
  assign n32 = ~x4 & x8 ;
  assign n33 = n31 & n32 ;
  assign n34 = n23 & n33 ;
  assign n35 = n30 & n34 ;
  assign n36 = ~n28 & ~n35 ;
  assign n37 = x1 & ~x12 ;
  assign n38 = ~x2 & n37 ;
  assign n39 = ~x3 & ~x11 ;
  assign n40 = ~x0 & n39 ;
  assign n41 = n38 & n40 ;
  assign n42 = ~n36 & n41 ;
  assign y0 = n42 ;
endmodule
