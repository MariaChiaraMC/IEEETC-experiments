// Benchmark "./pla/mlp4.pla_res_7NonExact" written by ABC on Fri Nov 20 10:27:01 2020

module \./pla/mlp4.pla_res_7NonExact  ( 
    x0, x1,
    z0  );
  input  x0, x1;
  output z0;
  assign z0 = x0 & x1;
endmodule


