module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 ;
  output y0 ;
  wire n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 ;
  assign n24 = x8 & ~x9 ;
  assign n25 = x7 & ~n24 ;
  assign n26 = ~x15 & ~x16 ;
  assign n27 = x10 & ~n26 ;
  assign n28 = ~x19 & ~x21 ;
  assign n29 = x13 & ~x14 ;
  assign n30 = n28 & n29 ;
  assign n31 = ~x20 & n30 ;
  assign n32 = ~n27 & ~n31 ;
  assign n33 = x20 & x21 ;
  assign n34 = ~x13 & x14 ;
  assign n35 = ~x16 & n34 ;
  assign n36 = ~n33 & n35 ;
  assign n37 = x15 & ~n36 ;
  assign n38 = ~x0 & ~x8 ;
  assign n39 = ~n37 & n38 ;
  assign n40 = ~x4 & ~x18 ;
  assign n41 = ~x2 & ~x3 ;
  assign n42 = n40 & n41 ;
  assign n43 = ~x5 & ~x9 ;
  assign n44 = n42 & n43 ;
  assign n45 = ~x12 & x22 ;
  assign n46 = ~x1 & n45 ;
  assign n47 = n46 ^ n44 ;
  assign n48 = x11 & x16 ;
  assign n49 = n48 ^ x10 ;
  assign n50 = n49 ^ n48 ;
  assign n51 = x16 & ~n34 ;
  assign n52 = ~x11 & ~x17 ;
  assign n53 = ~n51 & n52 ;
  assign n54 = n53 ^ n48 ;
  assign n55 = n50 & n54 ;
  assign n56 = n55 ^ n48 ;
  assign n57 = n56 ^ n44 ;
  assign n58 = n47 & n57 ;
  assign n59 = n58 ^ n55 ;
  assign n60 = n59 ^ n48 ;
  assign n61 = n60 ^ n46 ;
  assign n62 = n44 & n61 ;
  assign n63 = n62 ^ n44 ;
  assign n64 = n39 & n63 ;
  assign n65 = ~n32 & n64 ;
  assign n66 = ~n25 & ~n65 ;
  assign n67 = ~x6 & ~n66 ;
  assign y0 = n67 ;
endmodule
