module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 ;
  assign n25 = ~x6 & ~x11 ;
  assign n26 = ~x10 & n25 ;
  assign n30 = x9 & n26 ;
  assign n17 = ~x7 & ~x8 ;
  assign n18 = x6 & ~n17 ;
  assign n31 = x12 & n18 ;
  assign n20 = x8 ^ x7 ;
  assign n21 = x8 & ~n20 ;
  assign n22 = x6 & n21 ;
  assign n23 = n22 ^ n20 ;
  assign n32 = x5 & ~n23 ;
  assign n33 = ~n31 & ~n32 ;
  assign n34 = ~n30 & n33 ;
  assign n19 = x15 & n18 ;
  assign n24 = x13 & ~n23 ;
  assign n27 = x14 & n26 ;
  assign n28 = ~n24 & ~n27 ;
  assign n29 = ~n19 & n28 ;
  assign n35 = n34 ^ n29 ;
  assign n36 = n29 ^ x0 ;
  assign n37 = n36 ^ n35 ;
  assign n41 = x2 & ~x3 ;
  assign n42 = ~x4 & ~n41 ;
  assign n43 = ~x1 & ~n42 ;
  assign n38 = ~x2 & x3 ;
  assign n39 = x4 & ~n38 ;
  assign n40 = x1 & ~n39 ;
  assign n44 = n43 ^ n40 ;
  assign n45 = ~x0 & n44 ;
  assign n46 = n45 ^ n40 ;
  assign n47 = n37 & n46 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = n48 ^ n40 ;
  assign n50 = n49 ^ x0 ;
  assign n51 = n35 & ~n50 ;
  assign n52 = n51 ^ n34 ;
  assign y0 = ~n52 ;
endmodule
