module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 ;
  assign n11 = ~x0 & x6 ;
  assign n12 = x7 & x9 ;
  assign n13 = x2 & ~x3 ;
  assign n14 = ~x1 & x4 ;
  assign n15 = n13 & n14 ;
  assign n16 = n12 & n15 ;
  assign n17 = ~x8 & n16 ;
  assign n18 = x8 & ~x9 ;
  assign n19 = x4 & x7 ;
  assign n20 = n18 & ~n19 ;
  assign n21 = x1 & ~x2 ;
  assign n22 = ~x4 & ~x7 ;
  assign n23 = ~x3 & ~n22 ;
  assign n24 = n21 & n23 ;
  assign n25 = n20 & n24 ;
  assign n26 = x8 & x9 ;
  assign n27 = x3 & n26 ;
  assign n28 = x4 & ~x7 ;
  assign n29 = n21 & n28 ;
  assign n30 = n27 & n29 ;
  assign n31 = ~n25 & ~n30 ;
  assign n32 = ~n17 & n31 ;
  assign n33 = n11 & ~n32 ;
  assign n34 = ~x8 & x9 ;
  assign n35 = x0 & ~x6 ;
  assign n36 = n34 & n35 ;
  assign n37 = ~x3 & n29 ;
  assign n38 = n36 & n37 ;
  assign n39 = n38 ^ n33 ;
  assign n40 = x0 & ~x8 ;
  assign n41 = ~x6 & ~x7 ;
  assign n42 = n21 & n41 ;
  assign n43 = ~x4 & n42 ;
  assign n44 = x4 & x6 ;
  assign n45 = x7 & n44 ;
  assign n46 = ~x1 & x2 ;
  assign n47 = n45 & n46 ;
  assign n48 = ~n43 & ~n47 ;
  assign n49 = x3 & ~n48 ;
  assign n50 = n40 & n49 ;
  assign n51 = ~x0 & x7 ;
  assign n52 = x1 & x3 ;
  assign n53 = n51 & ~n52 ;
  assign n54 = x2 & x3 ;
  assign n55 = ~x3 & ~x4 ;
  assign n56 = ~n54 & ~n55 ;
  assign n57 = ~n14 & n56 ;
  assign n58 = n53 & n57 ;
  assign n59 = ~x1 & ~x3 ;
  assign n60 = ~x2 & ~x4 ;
  assign n61 = ~x7 & n60 ;
  assign n62 = ~n59 & n61 ;
  assign n63 = ~n15 & ~n62 ;
  assign n64 = x0 & ~n63 ;
  assign n65 = ~x0 & x2 ;
  assign n66 = ~x2 & x3 ;
  assign n67 = ~n65 & ~n66 ;
  assign n68 = n14 & n67 ;
  assign n69 = x7 & n68 ;
  assign n70 = ~n64 & ~n69 ;
  assign n71 = ~n58 & n70 ;
  assign n72 = ~x6 & ~n71 ;
  assign n73 = x0 & ~x7 ;
  assign n74 = ~x1 & ~x2 ;
  assign n75 = n73 & n74 ;
  assign n76 = x3 & n44 ;
  assign n77 = n75 & n76 ;
  assign n78 = ~x1 & ~n35 ;
  assign n79 = n22 & n78 ;
  assign n80 = n67 & n79 ;
  assign n81 = ~x9 & ~n80 ;
  assign n82 = ~n77 & n81 ;
  assign n83 = ~n72 & n82 ;
  assign n104 = ~n13 & ~n66 ;
  assign n84 = x4 ^ x2 ;
  assign n85 = n84 ^ x7 ;
  assign n86 = x7 ^ x0 ;
  assign n87 = n86 ^ n85 ;
  assign n88 = x7 ^ x4 ;
  assign n89 = n88 ^ x4 ;
  assign n90 = x4 ^ x3 ;
  assign n91 = n90 ^ x4 ;
  assign n92 = ~n89 & n91 ;
  assign n93 = n92 ^ x4 ;
  assign n94 = n93 ^ n85 ;
  assign n95 = n87 & ~n94 ;
  assign n96 = n95 ^ n92 ;
  assign n97 = n96 ^ x4 ;
  assign n98 = n97 ^ n86 ;
  assign n99 = n85 & ~n98 ;
  assign n100 = n99 ^ n85 ;
  assign n105 = n104 ^ n100 ;
  assign n106 = n105 ^ n100 ;
  assign n101 = ~x7 & ~n65 ;
  assign n102 = n101 ^ n100 ;
  assign n103 = n102 ^ n100 ;
  assign n107 = n106 ^ n103 ;
  assign n108 = n100 ^ x4 ;
  assign n109 = n108 ^ n100 ;
  assign n110 = n109 ^ n106 ;
  assign n111 = ~n106 & ~n110 ;
  assign n112 = n111 ^ n106 ;
  assign n113 = n107 & ~n112 ;
  assign n114 = n113 ^ n111 ;
  assign n115 = n114 ^ n100 ;
  assign n116 = n115 ^ n106 ;
  assign n117 = ~x1 & ~n116 ;
  assign n118 = n117 ^ n100 ;
  assign n119 = n118 ^ x6 ;
  assign n120 = n119 ^ n118 ;
  assign n121 = n120 ^ x9 ;
  assign n122 = x7 ^ x1 ;
  assign n123 = n122 ^ n84 ;
  assign n124 = x4 ^ x0 ;
  assign n125 = ~n86 & ~n124 ;
  assign n126 = n125 ^ x0 ;
  assign n127 = n126 ^ n122 ;
  assign n128 = ~n123 & n127 ;
  assign n129 = n128 ^ n125 ;
  assign n130 = n129 ^ x0 ;
  assign n131 = n130 ^ n84 ;
  assign n132 = ~n122 & ~n131 ;
  assign n133 = n132 ^ n122 ;
  assign n134 = n133 ^ x3 ;
  assign n135 = ~n133 & ~n134 ;
  assign n136 = n135 ^ n118 ;
  assign n137 = n136 ^ n133 ;
  assign n138 = ~n121 & ~n137 ;
  assign n139 = n138 ^ n135 ;
  assign n140 = n139 ^ n133 ;
  assign n141 = x9 & ~n140 ;
  assign n142 = n141 ^ x9 ;
  assign n143 = ~n83 & ~n142 ;
  assign n144 = n143 ^ x8 ;
  assign n145 = n144 ^ n143 ;
  assign n150 = ~x6 & x7 ;
  assign n151 = ~x2 & n150 ;
  assign n152 = n55 & n151 ;
  assign n146 = ~x4 & ~x6 ;
  assign n147 = n54 & n146 ;
  assign n148 = ~x3 & n45 ;
  assign n149 = ~n147 & ~n148 ;
  assign n153 = n152 ^ n149 ;
  assign n154 = n153 ^ n149 ;
  assign n155 = n44 & n54 ;
  assign n156 = ~x7 & n155 ;
  assign n157 = n156 ^ n149 ;
  assign n158 = n157 ^ n149 ;
  assign n159 = ~n154 & ~n158 ;
  assign n160 = n159 ^ n149 ;
  assign n161 = x1 & n160 ;
  assign n162 = n161 ^ n149 ;
  assign n163 = n162 ^ x0 ;
  assign n164 = n163 ^ n162 ;
  assign n165 = ~x3 & x7 ;
  assign n166 = ~n28 & ~n165 ;
  assign n167 = x3 & ~x4 ;
  assign n168 = x6 & ~n167 ;
  assign n169 = n46 & n168 ;
  assign n170 = n166 & n169 ;
  assign n171 = ~x4 & x7 ;
  assign n172 = x1 & x2 ;
  assign n173 = n171 & n172 ;
  assign n174 = ~x6 & n173 ;
  assign n175 = x3 & x4 ;
  assign n176 = ~n55 & ~n175 ;
  assign n177 = n42 & ~n176 ;
  assign n178 = ~n174 & ~n177 ;
  assign n179 = ~n170 & n178 ;
  assign n180 = n179 ^ n162 ;
  assign n181 = ~n164 & n180 ;
  assign n182 = n181 ^ n162 ;
  assign n183 = ~n77 & n182 ;
  assign n184 = ~x9 & ~n183 ;
  assign n185 = ~x2 & n12 ;
  assign n186 = n146 ^ n52 ;
  assign n187 = n186 ^ n52 ;
  assign n188 = n187 ^ x0 ;
  assign n189 = n59 ^ n44 ;
  assign n190 = ~n44 & ~n189 ;
  assign n191 = n190 ^ n52 ;
  assign n192 = n191 ^ n44 ;
  assign n193 = n188 & ~n192 ;
  assign n194 = n193 ^ n190 ;
  assign n195 = n194 ^ n44 ;
  assign n196 = ~x0 & ~n195 ;
  assign n197 = n196 ^ x0 ;
  assign n198 = n185 & n197 ;
  assign n199 = n198 ^ x0 ;
  assign n200 = n167 & n172 ;
  assign n201 = n41 & n200 ;
  assign n202 = n46 & n150 ;
  assign n203 = ~n176 & n202 ;
  assign n204 = x9 & n203 ;
  assign n205 = ~n201 & ~n204 ;
  assign n206 = n205 ^ n198 ;
  assign n207 = n206 ^ n205 ;
  assign n208 = x3 ^ x1 ;
  assign n209 = n44 ^ x3 ;
  assign n210 = n209 ^ n44 ;
  assign n211 = n146 ^ n44 ;
  assign n212 = ~n210 & n211 ;
  assign n213 = n212 ^ n44 ;
  assign n214 = ~n208 & n213 ;
  assign n215 = n214 ^ n205 ;
  assign n216 = n207 & n215 ;
  assign n217 = n216 ^ n205 ;
  assign n218 = ~n199 & n217 ;
  assign n219 = n218 ^ x0 ;
  assign n220 = ~n184 & n219 ;
  assign n221 = n220 ^ n143 ;
  assign n222 = n145 & ~n221 ;
  assign n223 = n222 ^ n143 ;
  assign n224 = ~n50 & ~n223 ;
  assign n225 = n224 ^ x5 ;
  assign n226 = n225 ^ n224 ;
  assign n227 = ~x6 & n13 ;
  assign n228 = ~x0 & ~x8 ;
  assign n229 = n22 & n228 ;
  assign n230 = n227 & n229 ;
  assign n231 = x7 ^ x2 ;
  assign n232 = n231 ^ x8 ;
  assign n233 = n232 ^ x9 ;
  assign n235 = x8 ^ x7 ;
  assign n234 = x9 ^ x8 ;
  assign n236 = n235 ^ n234 ;
  assign n237 = n236 ^ n233 ;
  assign n238 = n235 ^ x6 ;
  assign n239 = n235 ^ x9 ;
  assign n240 = n239 ^ n238 ;
  assign n241 = n238 & ~n240 ;
  assign n242 = n241 ^ n235 ;
  assign n243 = n242 ^ n238 ;
  assign n244 = n237 & ~n243 ;
  assign n245 = n244 ^ n241 ;
  assign n246 = n245 ^ n238 ;
  assign n247 = n233 & n246 ;
  assign n248 = n167 & n247 ;
  assign n249 = ~x8 & ~x9 ;
  assign n250 = x4 & n249 ;
  assign n251 = ~n26 & ~n250 ;
  assign n252 = n151 & ~n251 ;
  assign n253 = x3 & n252 ;
  assign n254 = n249 ^ n26 ;
  assign n255 = n26 ^ x4 ;
  assign n256 = n255 ^ n26 ;
  assign n257 = n254 & ~n256 ;
  assign n258 = n257 ^ n26 ;
  assign n259 = x6 & n258 ;
  assign n260 = n259 ^ x2 ;
  assign n261 = n260 ^ n259 ;
  assign n262 = x4 & ~x6 ;
  assign n263 = n18 & n262 ;
  assign n264 = n263 ^ n259 ;
  assign n265 = n261 & n264 ;
  assign n266 = n265 ^ n259 ;
  assign n267 = n165 & n266 ;
  assign n268 = ~n253 & ~n267 ;
  assign n269 = ~n248 & n268 ;
  assign n270 = ~x0 & ~n269 ;
  assign n271 = ~x7 & n249 ;
  assign n272 = n147 & n271 ;
  assign n273 = ~x4 & x6 ;
  assign n274 = n34 & n273 ;
  assign n275 = ~n263 & ~n274 ;
  assign n276 = n54 & ~n275 ;
  assign n277 = ~x3 & x6 ;
  assign n278 = n18 & n277 ;
  assign n279 = x3 & ~x6 ;
  assign n280 = n26 & n279 ;
  assign n281 = ~n278 & ~n280 ;
  assign n282 = n60 & ~n281 ;
  assign n283 = ~n276 & ~n282 ;
  assign n284 = n73 & ~n283 ;
  assign n285 = x4 & n54 ;
  assign n286 = n36 & n285 ;
  assign n287 = ~n284 & ~n286 ;
  assign n288 = ~n272 & n287 ;
  assign n289 = ~n270 & n288 ;
  assign n290 = n289 ^ x1 ;
  assign n291 = n290 ^ n289 ;
  assign n292 = ~x8 & n171 ;
  assign n293 = n18 & n73 ;
  assign n294 = ~n292 & ~n293 ;
  assign n295 = n227 & ~n294 ;
  assign n296 = n11 & ~n13 ;
  assign n297 = x7 & n249 ;
  assign n298 = n176 & n297 ;
  assign n299 = n296 & n298 ;
  assign n300 = n26 ^ x6 ;
  assign n301 = ~n22 & ~n51 ;
  assign n302 = n301 ^ x3 ;
  assign n303 = n302 ^ n301 ;
  assign n304 = n301 ^ n28 ;
  assign n305 = ~n303 & ~n304 ;
  assign n306 = n305 ^ n301 ;
  assign n307 = n306 ^ n26 ;
  assign n308 = n300 & ~n307 ;
  assign n309 = n308 ^ n305 ;
  assign n310 = n309 ^ n301 ;
  assign n311 = n310 ^ x6 ;
  assign n312 = n26 & ~n311 ;
  assign n313 = n312 ^ n26 ;
  assign n314 = x2 & n313 ;
  assign n315 = x2 & x4 ;
  assign n316 = ~n165 & n315 ;
  assign n317 = n40 & n316 ;
  assign n318 = x6 & x7 ;
  assign n319 = n318 ^ n316 ;
  assign n320 = ~x3 & x9 ;
  assign n321 = n320 ^ n317 ;
  assign n322 = ~n319 & n321 ;
  assign n323 = n322 ^ n320 ;
  assign n324 = n317 & n323 ;
  assign n325 = ~n314 & ~n324 ;
  assign n326 = ~n299 & n325 ;
  assign n327 = n26 & ~n176 ;
  assign n328 = x0 & ~n327 ;
  assign n329 = n175 & n271 ;
  assign n330 = ~n73 & ~n329 ;
  assign n331 = ~n328 & ~n330 ;
  assign n332 = n34 & n51 ;
  assign n333 = n167 & n332 ;
  assign n334 = ~n331 & ~n333 ;
  assign n335 = n334 ^ x2 ;
  assign n336 = n335 ^ n334 ;
  assign n337 = n336 ^ x6 ;
  assign n338 = n18 & n51 ;
  assign n339 = n175 ^ x6 ;
  assign n340 = n338 & n339 ;
  assign n341 = n340 ^ n334 ;
  assign n342 = ~n337 & ~n341 ;
  assign n343 = n342 ^ n340 ;
  assign n344 = x6 & n343 ;
  assign n345 = n344 ^ n340 ;
  assign n346 = n345 ^ n342 ;
  assign n347 = n326 & ~n346 ;
  assign n348 = ~n295 & n347 ;
  assign n349 = n348 ^ n289 ;
  assign n350 = n291 & n349 ;
  assign n351 = n350 ^ n289 ;
  assign n352 = ~n230 & n351 ;
  assign n353 = n352 ^ n224 ;
  assign n354 = n226 & n353 ;
  assign n355 = n354 ^ n224 ;
  assign n356 = n355 ^ n33 ;
  assign n357 = n39 & ~n356 ;
  assign n358 = n357 ^ n354 ;
  assign n359 = n358 ^ n224 ;
  assign n360 = n359 ^ n38 ;
  assign n361 = ~n33 & ~n360 ;
  assign n362 = n361 ^ n33 ;
  assign y0 = n362 ;
endmodule
