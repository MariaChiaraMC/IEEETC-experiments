module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n7 = x4 ^ x3 ;
  assign n8 = n7 ^ x2 ;
  assign n9 = n8 ^ x1 ;
  assign n15 = n9 ^ n7 ;
  assign n10 = n8 ^ x4 ;
  assign n11 = n10 ^ x5 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = n12 ^ x1 ;
  assign n14 = n13 ^ n9 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n10 ^ n7 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n18 ^ n9 ;
  assign n21 = n19 & ~n20 ;
  assign n22 = n21 ^ n13 ;
  assign n23 = n22 ^ n15 ;
  assign n24 = n7 ^ x1 ;
  assign n25 = n24 ^ n17 ;
  assign n26 = n25 ^ n13 ;
  assign n27 = ~n9 & ~n26 ;
  assign n28 = n27 ^ n9 ;
  assign n29 = n28 ^ n15 ;
  assign n30 = n23 & ~n29 ;
  assign n31 = ~n16 & n30 ;
  assign n32 = n31 ^ n21 ;
  assign n33 = n32 ^ n27 ;
  assign n34 = n33 ^ n17 ;
  assign n35 = n34 ^ n13 ;
  assign n36 = n35 ^ n15 ;
  assign n37 = n36 ^ x2 ;
  assign y0 = n37 ;
endmodule
