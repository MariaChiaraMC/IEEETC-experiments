module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 ;
  assign n8 = ~x0 & x4 ;
  assign n9 = x1 & x5 ;
  assign n10 = ~n8 & ~n9 ;
  assign n11 = x3 & x6 ;
  assign n12 = ~x0 & x1 ;
  assign n13 = n11 & ~n12 ;
  assign n14 = ~n10 & n13 ;
  assign n15 = ~x4 & ~x5 ;
  assign n16 = n15 ^ x6 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n17 ^ x0 ;
  assign n19 = x1 & ~x3 ;
  assign n20 = n15 ^ x0 ;
  assign n21 = ~n17 & n20 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = n19 & n22 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n18 & n24 ;
  assign n26 = n25 ^ n21 ;
  assign n32 = x5 ^ x3 ;
  assign n28 = x5 ^ x4 ;
  assign n27 = x5 ^ x0 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ x5 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ x5 ;
  assign n46 = n34 ^ n30 ;
  assign n37 = n30 ^ n27 ;
  assign n38 = n37 ^ n32 ;
  assign n42 = n38 ^ n34 ;
  assign n47 = n42 ^ n30 ;
  assign n48 = ~n46 & n47 ;
  assign n55 = n48 ^ n34 ;
  assign n56 = n55 ^ n38 ;
  assign n35 = x6 ^ x5 ;
  assign n36 = n35 ^ n34 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n39 ^ n30 ;
  assign n57 = n56 ^ n40 ;
  assign n43 = n42 ^ n40 ;
  assign n44 = n40 ^ n38 ;
  assign n45 = ~n43 & ~n44 ;
  assign n58 = n45 ^ n34 ;
  assign n59 = n58 ^ n38 ;
  assign n60 = n59 ^ n30 ;
  assign n61 = ~n57 & n60 ;
  assign n31 = n30 ^ x6 ;
  assign n41 = n40 ^ n31 ;
  assign n49 = n48 ^ n45 ;
  assign n50 = n49 ^ n34 ;
  assign n51 = n50 ^ n38 ;
  assign n52 = n51 ^ n30 ;
  assign n53 = n52 ^ n40 ;
  assign n54 = ~n41 & n53 ;
  assign n62 = n61 ^ n54 ;
  assign n63 = n62 ^ n30 ;
  assign n64 = n63 ^ n40 ;
  assign n65 = n64 ^ x0 ;
  assign n66 = n65 ^ x5 ;
  assign n67 = n66 ^ x1 ;
  assign n68 = n67 ^ n66 ;
  assign n69 = n68 ^ n26 ;
  assign n70 = x4 & x6 ;
  assign n71 = n70 ^ x0 ;
  assign n72 = n71 ^ x5 ;
  assign n73 = ~x5 & n72 ;
  assign n74 = n73 ^ n66 ;
  assign n75 = n74 ^ x5 ;
  assign n76 = ~n69 & ~n75 ;
  assign n77 = n76 ^ n73 ;
  assign n78 = n77 ^ x5 ;
  assign n79 = ~n26 & ~n78 ;
  assign n80 = n79 ^ n26 ;
  assign n81 = n80 ^ x2 ;
  assign n82 = n81 ^ n80 ;
  assign n83 = x3 & x5 ;
  assign n84 = ~x0 & ~n83 ;
  assign n85 = ~x3 & x6 ;
  assign n86 = x0 & ~n85 ;
  assign n87 = n86 ^ x1 ;
  assign n88 = n86 ^ x4 ;
  assign n89 = n88 ^ x4 ;
  assign n90 = n15 ^ x4 ;
  assign n91 = n89 & n90 ;
  assign n92 = n91 ^ x4 ;
  assign n93 = n87 & n92 ;
  assign n94 = n93 ^ x1 ;
  assign n95 = ~n84 & n94 ;
  assign n96 = x1 & ~x5 ;
  assign n97 = n96 ^ x5 ;
  assign n98 = n97 ^ x5 ;
  assign n99 = n28 ^ x5 ;
  assign n100 = n98 & n99 ;
  assign n101 = n100 ^ x5 ;
  assign n102 = x6 & n101 ;
  assign n103 = n102 ^ x5 ;
  assign n104 = ~x0 & n103 ;
  assign n105 = ~x0 & ~n70 ;
  assign n106 = ~x5 & x6 ;
  assign n107 = ~x4 & ~n106 ;
  assign n108 = n105 & ~n107 ;
  assign n109 = ~x1 & n108 ;
  assign n110 = ~x1 & ~n15 ;
  assign n111 = ~n8 & n85 ;
  assign n112 = n110 & n111 ;
  assign n113 = ~n109 & ~n112 ;
  assign n114 = ~n104 & n113 ;
  assign n115 = ~n95 & n114 ;
  assign n116 = n115 ^ n80 ;
  assign n117 = n82 & ~n116 ;
  assign n118 = n117 ^ n80 ;
  assign n119 = ~n14 & ~n118 ;
  assign y0 = ~n119 ;
endmodule
