module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;
  assign n9 = x5 ^ x3 ;
  assign n10 = x6 ^ x5 ;
  assign n11 = x4 & ~x7 ;
  assign n12 = n11 ^ x5 ;
  assign n13 = n12 ^ x5 ;
  assign n14 = n10 & n13 ;
  assign n15 = n14 ^ x5 ;
  assign n16 = ~n9 & n15 ;
  assign n17 = n16 ^ x3 ;
  assign n18 = ~x1 & ~x3 ;
  assign n19 = x7 ^ x6 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = x5 ^ x4 ;
  assign n22 = ~x6 & n21 ;
  assign n23 = n22 ^ x4 ;
  assign n24 = ~n20 & ~n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = n26 ^ x6 ;
  assign n28 = n18 & n27 ;
  assign n29 = ~n17 & ~n28 ;
  assign n30 = ~x2 & ~n29 ;
  assign n31 = x2 & ~x3 ;
  assign n32 = x5 & x7 ;
  assign n33 = n31 & n32 ;
  assign n34 = x2 ^ x1 ;
  assign n35 = x5 & x6 ;
  assign n36 = ~x4 & ~n35 ;
  assign n37 = n36 ^ x1 ;
  assign n38 = n34 & ~n37 ;
  assign n39 = ~x3 & n38 ;
  assign n40 = n39 ^ x1 ;
  assign n41 = ~x0 & ~n40 ;
  assign n42 = ~n33 & n41 ;
  assign n43 = ~n30 & n42 ;
  assign y0 = n43 ;
endmodule
