module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 ;
  assign n9 = x2 ^ x1 ;
  assign n10 = n9 ^ x2 ;
  assign n11 = x4 & ~x5 ;
  assign n12 = x3 & ~n11 ;
  assign n13 = x3 ^ x2 ;
  assign n14 = n13 ^ x3 ;
  assign n15 = x5 ^ x4 ;
  assign n16 = n15 ^ x3 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n17 ^ x6 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = n20 ^ x3 ;
  assign n22 = ~n14 & n21 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n20 ^ x4 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n18 ^ x6 ;
  assign n27 = n26 ^ x7 ;
  assign n28 = n27 ^ x7 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = ~n20 & ~n29 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = ~n25 & ~n32 ;
  assign n34 = n33 ^ n20 ;
  assign n35 = ~n23 & ~n34 ;
  assign n36 = n35 ^ n22 ;
  assign n37 = n36 ^ n20 ;
  assign n38 = n37 ^ x2 ;
  assign n39 = ~n12 & ~n38 ;
  assign n40 = n39 ^ x2 ;
  assign n41 = ~n10 & ~n40 ;
  assign n42 = n41 ^ x2 ;
  assign n43 = ~x5 & ~x6 ;
  assign n44 = ~x7 & ~n43 ;
  assign n45 = x5 & x6 ;
  assign n46 = ~x3 & x4 ;
  assign n47 = ~n45 & n46 ;
  assign n48 = ~n44 & n47 ;
  assign n49 = x2 & n48 ;
  assign n50 = n49 ^ x0 ;
  assign n51 = n42 & ~n50 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = ~x0 & n52 ;
  assign n54 = n53 ^ x0 ;
  assign y0 = ~n54 ;
endmodule
