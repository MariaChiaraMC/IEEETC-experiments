// Benchmark "./addm4.pla" written by ABC on Thu Apr 23 10:59:45 2020

module \./addm4.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8,
    z7  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8;
  output z7;
  assign z7 = ~x0 | x4;
endmodule


