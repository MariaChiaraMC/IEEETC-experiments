module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 ;
  assign n17 = x9 & x15 ;
  assign n18 = x4 & x12 ;
  assign n19 = x10 & n18 ;
  assign n20 = x11 & x13 ;
  assign n21 = x14 & n20 ;
  assign n22 = x15 & ~n21 ;
  assign n23 = ~x2 & ~n22 ;
  assign n25 = x3 & ~x6 ;
  assign n24 = x7 & x8 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = n25 ^ x0 ;
  assign n29 = n28 ^ n25 ;
  assign n30 = n27 & ~n29 ;
  assign n31 = n30 ^ n25 ;
  assign n32 = x1 & n31 ;
  assign n33 = n32 ^ n25 ;
  assign n34 = n23 & n33 ;
  assign n35 = ~x14 & x15 ;
  assign n36 = ~x11 & ~n35 ;
  assign n37 = x13 & ~n36 ;
  assign n38 = x2 ^ x0 ;
  assign n39 = x3 ^ x2 ;
  assign n40 = n39 ^ x3 ;
  assign n41 = x7 ^ x3 ;
  assign n42 = n40 & ~n41 ;
  assign n43 = n42 ^ x3 ;
  assign n44 = n38 & ~n43 ;
  assign n45 = ~n37 & n44 ;
  assign n46 = ~x1 & n45 ;
  assign n47 = ~n34 & ~n46 ;
  assign n48 = n47 ^ x5 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = ~x0 & x1 ;
  assign n51 = x15 ^ x11 ;
  assign n52 = n51 ^ x13 ;
  assign n53 = n52 ^ n51 ;
  assign n56 = n51 ^ x3 ;
  assign n57 = n51 & n56 ;
  assign n54 = x14 & x15 ;
  assign n60 = n57 ^ n54 ;
  assign n55 = n54 ^ n53 ;
  assign n58 = n57 ^ n51 ;
  assign n59 = ~n55 & n58 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = ~n53 & n61 ;
  assign n63 = n62 ^ n57 ;
  assign n64 = n63 ^ n59 ;
  assign n65 = n64 ^ x15 ;
  assign n66 = n50 & ~n65 ;
  assign n67 = x2 & n66 ;
  assign n68 = n67 ^ n47 ;
  assign n69 = n49 & ~n68 ;
  assign n70 = n69 ^ n47 ;
  assign n71 = n19 & ~n70 ;
  assign n72 = ~n17 & ~n71 ;
  assign y0 = ~n72 ;
endmodule
