module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 ;
  assign n15 = x3 ^ x1 ;
  assign n16 = n15 ^ x3 ;
  assign n17 = x4 & ~x5 ;
  assign n18 = n17 ^ x3 ;
  assign n19 = ~n16 & ~n18 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = ~x6 & n20 ;
  assign n22 = n21 ^ x1 ;
  assign n23 = ~x2 & ~n22 ;
  assign n24 = x4 ^ x3 ;
  assign n25 = n24 ^ x6 ;
  assign n26 = n25 ^ x6 ;
  assign n30 = x3 ^ x2 ;
  assign n27 = x5 ^ x3 ;
  assign n32 = n30 ^ n27 ;
  assign n28 = n27 ^ x6 ;
  assign n29 = n28 ^ x3 ;
  assign n31 = n30 ^ n29 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = ~n26 & ~n33 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n35 ^ n29 ;
  assign n37 = n36 ^ x3 ;
  assign n38 = n37 ^ n32 ;
  assign n39 = n32 ^ x3 ;
  assign n40 = x6 ^ x1 ;
  assign n41 = n40 ^ x3 ;
  assign n42 = n41 ^ n26 ;
  assign n43 = ~n39 & n42 ;
  assign n44 = n43 ^ n29 ;
  assign n45 = n44 ^ n26 ;
  assign n46 = n45 ^ n32 ;
  assign n47 = n32 ^ n26 ;
  assign n48 = n29 ^ n26 ;
  assign n49 = n48 ^ n32 ;
  assign n50 = n47 & ~n49 ;
  assign n51 = n50 ^ n26 ;
  assign n52 = ~n46 & ~n51 ;
  assign n53 = n52 ^ n30 ;
  assign n54 = n53 ^ n32 ;
  assign n55 = ~n38 & n54 ;
  assign n56 = n55 ^ n52 ;
  assign n57 = n56 ^ n30 ;
  assign n58 = n57 ^ n32 ;
  assign n59 = n58 ^ x3 ;
  assign n60 = ~n23 & n59 ;
  assign n61 = ~x1 & x3 ;
  assign n62 = x1 & ~x6 ;
  assign n63 = ~x2 & ~n62 ;
  assign n64 = ~n61 & ~n63 ;
  assign n65 = n64 ^ x4 ;
  assign n66 = n65 ^ n64 ;
  assign n67 = n66 ^ x5 ;
  assign n68 = ~x7 & ~x9 ;
  assign n69 = ~x11 & ~x12 ;
  assign n70 = ~n68 & n69 ;
  assign n71 = x3 & ~x8 ;
  assign n72 = x2 & ~x10 ;
  assign n73 = ~x13 & n72 ;
  assign n74 = n71 & n73 ;
  assign n75 = n70 & n74 ;
  assign n76 = x1 & ~n75 ;
  assign n77 = x6 & ~n76 ;
  assign n78 = n77 ^ n62 ;
  assign n79 = ~n62 & n78 ;
  assign n80 = n79 ^ n64 ;
  assign n81 = n80 ^ n62 ;
  assign n82 = n67 & ~n81 ;
  assign n83 = n82 ^ n79 ;
  assign n84 = n83 ^ n62 ;
  assign n85 = x5 & ~n84 ;
  assign n86 = n85 ^ x5 ;
  assign n87 = n60 & ~n86 ;
  assign n88 = ~x0 & ~n87 ;
  assign y0 = n88 ;
endmodule
