module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 ;
  assign n16 = x1 & x6 ;
  assign n15 = x3 ^ x2 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n15 ^ x3 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n21 ^ n15 ;
  assign n23 = n22 ^ n15 ;
  assign n24 = n18 & n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n22 ^ x4 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = ~x10 & ~x11 ;
  assign n29 = x9 & ~x12 ;
  assign n30 = n28 & n29 ;
  assign n31 = ~x8 & ~x13 ;
  assign n32 = n30 & n31 ;
  assign n33 = ~x7 & n32 ;
  assign n34 = n33 ^ x1 ;
  assign n35 = ~n22 & ~n34 ;
  assign n36 = n35 ^ x1 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = ~n27 & ~n37 ;
  assign n39 = n38 ^ n22 ;
  assign n40 = ~n25 & ~n39 ;
  assign n41 = n40 ^ n24 ;
  assign n42 = n41 ^ n22 ;
  assign n43 = n42 ^ x3 ;
  assign n44 = x2 & ~x3 ;
  assign n45 = n44 ^ x5 ;
  assign n46 = n45 ^ x0 ;
  assign n47 = ~x4 & ~x6 ;
  assign n48 = ~x3 & ~n47 ;
  assign n49 = n48 ^ n44 ;
  assign n50 = n49 ^ n48 ;
  assign n51 = x4 & ~n16 ;
  assign n52 = n51 ^ n48 ;
  assign n53 = n50 & n52 ;
  assign n54 = n53 ^ n48 ;
  assign n55 = n54 ^ n45 ;
  assign n56 = n46 & n55 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n57 ^ n48 ;
  assign n59 = n58 ^ x0 ;
  assign n60 = ~n45 & n59 ;
  assign n61 = n60 ^ n45 ;
  assign n62 = n61 ^ x0 ;
  assign n63 = n43 & n62 ;
  assign y0 = n63 ;
endmodule
