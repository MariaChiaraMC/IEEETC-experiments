module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
  assign n11 = ~x2 & ~x3 ;
  assign n12 = ~x0 & n11 ;
  assign n13 = ~x4 & ~x5 ;
  assign n14 = ~x1 & n13 ;
  assign n15 = n14 ^ x6 ;
  assign n16 = x7 & x8 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = x8 & ~x9 ;
  assign n20 = ~x8 & x9 ;
  assign n21 = n20 ^ x7 ;
  assign n22 = n13 & n21 ;
  assign n23 = ~n19 & n22 ;
  assign n24 = ~x7 & n20 ;
  assign n25 = ~n16 & ~n24 ;
  assign n26 = ~x4 & ~n25 ;
  assign n27 = ~x5 & n21 ;
  assign n28 = ~n26 & ~n27 ;
  assign n29 = ~x1 & ~n28 ;
  assign n30 = ~n23 & ~n29 ;
  assign n31 = n30 ^ n16 ;
  assign n32 = ~n18 & ~n31 ;
  assign n33 = n32 ^ n16 ;
  assign n34 = ~n15 & n33 ;
  assign n35 = n12 & n34 ;
  assign y0 = n35 ;
endmodule
