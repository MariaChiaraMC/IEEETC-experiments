module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
  assign n11 = x5 ^ x4 ;
  assign n12 = x7 & x8 ;
  assign n13 = ~x2 & x9 ;
  assign n14 = n12 & n13 ;
  assign n15 = n14 ^ x4 ;
  assign n16 = n15 ^ x4 ;
  assign n17 = n16 ^ n11 ;
  assign n18 = ~n11 & ~n17 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = n19 ^ n11 ;
  assign n21 = x3 & ~x6 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = n22 ^ x0 ;
  assign n24 = n21 & n23 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = n21 ^ x1 ;
  assign n28 = ~n22 & n27 ;
  assign n29 = n28 ^ x1 ;
  assign n30 = n29 ^ x0 ;
  assign n31 = ~n26 & ~n30 ;
  assign n32 = n31 ^ x0 ;
  assign n33 = n20 & ~n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n34 ^ x0 ;
  assign y0 = ~n35 ;
endmodule
