module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 ;
  assign n9 = ~x1 & ~x3 ;
  assign n10 = x4 & n9 ;
  assign n11 = x2 & ~n10 ;
  assign n12 = ~x2 & x6 ;
  assign n13 = x4 & ~n12 ;
  assign n15 = ~x3 & ~x6 ;
  assign n14 = ~x6 & ~x7 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n15 ^ x3 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n17 & ~n19 ;
  assign n21 = n20 ^ n15 ;
  assign n22 = ~x1 & ~n21 ;
  assign n23 = n22 ^ n15 ;
  assign n24 = ~n13 & n23 ;
  assign n25 = ~x3 & ~x7 ;
  assign n26 = ~x4 & n25 ;
  assign n27 = ~x1 & ~n26 ;
  assign n28 = n27 ^ x5 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ n24 ;
  assign n31 = ~x3 & x4 ;
  assign n32 = ~n25 & ~n31 ;
  assign n33 = ~n14 & ~n15 ;
  assign n34 = n33 ^ n32 ;
  assign n35 = n32 & n34 ;
  assign n36 = n35 ^ n27 ;
  assign n37 = n36 ^ n32 ;
  assign n38 = ~n30 & ~n37 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n39 ^ n32 ;
  assign n41 = n24 & n40 ;
  assign n42 = n41 ^ n24 ;
  assign n43 = ~n11 & ~n42 ;
  assign n44 = x6 & n9 ;
  assign n45 = n44 ^ x5 ;
  assign n46 = n45 ^ n44 ;
  assign n47 = ~x1 & ~x7 ;
  assign n48 = x3 & ~n47 ;
  assign n49 = ~x6 & ~n9 ;
  assign n50 = ~n48 & n49 ;
  assign n51 = ~x4 & n50 ;
  assign n52 = n51 ^ n44 ;
  assign n53 = ~n46 & n52 ;
  assign n54 = n53 ^ n44 ;
  assign n55 = x2 & n54 ;
  assign n56 = ~n43 & ~n55 ;
  assign n57 = ~x0 & ~n56 ;
  assign y0 = n57 ;
endmodule
