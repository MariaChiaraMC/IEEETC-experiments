module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 ;
  assign n9 = ~x0 & ~x1 ;
  assign n13 = x3 ^ x2 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = n14 ^ x2 ;
  assign n10 = x5 ^ x4 ;
  assign n11 = n10 ^ x2 ;
  assign n12 = n11 ^ x2 ;
  assign n16 = n15 ^ n12 ;
  assign n24 = n14 ^ x6 ;
  assign n25 = n24 ^ n10 ;
  assign n18 = x5 ^ x2 ;
  assign n19 = n18 ^ n14 ;
  assign n26 = n25 ^ n19 ;
  assign n20 = n19 ^ n10 ;
  assign n21 = n20 ^ n14 ;
  assign n22 = n21 ^ x2 ;
  assign n17 = n12 ^ n11 ;
  assign n23 = n22 ^ n17 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = ~n16 & n27 ;
  assign n29 = n28 ^ n11 ;
  assign n30 = n29 ^ n15 ;
  assign n31 = n22 ^ n15 ;
  assign n32 = n26 & n31 ;
  assign n33 = n32 ^ n15 ;
  assign n34 = n33 ^ n12 ;
  assign n35 = n14 ^ x7 ;
  assign n36 = n35 ^ n19 ;
  assign n37 = n36 ^ n15 ;
  assign n38 = n37 ^ n12 ;
  assign n39 = ~n22 & n38 ;
  assign n40 = n39 ^ n11 ;
  assign n41 = n40 ^ n15 ;
  assign n42 = n41 ^ n12 ;
  assign n43 = ~n34 & n42 ;
  assign n44 = n43 ^ n11 ;
  assign n45 = n44 ^ n15 ;
  assign n46 = n45 ^ n12 ;
  assign n47 = n30 & n46 ;
  assign n48 = n47 ^ x2 ;
  assign n49 = n9 & ~n48 ;
  assign y0 = n49 ;
endmodule
