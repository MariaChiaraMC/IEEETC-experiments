module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 ;
  assign n10 = x1 & x3 ;
  assign n11 = x5 & x7 ;
  assign n12 = ~n10 & ~n11 ;
  assign n13 = ~x0 & ~x8 ;
  assign n14 = ~n12 & n13 ;
  assign n15 = ~x2 & ~x6 ;
  assign n18 = n15 ^ x3 ;
  assign n19 = n18 ^ x5 ;
  assign n16 = n15 ^ x7 ;
  assign n17 = n16 ^ x1 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n20 ^ n15 ;
  assign n22 = n19 ^ x1 ;
  assign n23 = n22 ^ n15 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n24 ^ n17 ;
  assign n26 = ~n19 & ~n25 ;
  assign n27 = n26 ^ n15 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = n23 ^ n19 ;
  assign n30 = n29 ^ n21 ;
  assign n31 = ~n15 & n30 ;
  assign n32 = n31 ^ n19 ;
  assign n33 = ~n28 & ~n32 ;
  assign n34 = n21 & n33 ;
  assign n35 = n34 ^ n26 ;
  assign n36 = n35 ^ n31 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ n15 ;
  assign n39 = ~n14 & ~n38 ;
  assign n40 = x4 & ~n39 ;
  assign y0 = n40 ;
endmodule
