// Benchmark "./pla/pdc.pla_res_14NonExact" written by ABC on Fri Nov 20 10:29:06 2020

module \./pla/pdc.pla_res_14NonExact  ( 
    x0, x1,
    z0  );
  input  x0, x1;
  output z0;
  assign z0 = x0 & ~x1;
endmodule


