module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 ;
  output y0 ;
  wire n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 ;
  assign n24 = ~x12 & ~x13 ;
  assign n25 = x14 & ~x17 ;
  assign n26 = n24 & n25 ;
  assign n27 = x16 ^ x15 ;
  assign n28 = x20 & x21 ;
  assign n29 = ~x16 & n28 ;
  assign n30 = n27 & n29 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n26 & n31 ;
  assign n33 = ~x11 & ~n32 ;
  assign n34 = ~x4 & ~x7 ;
  assign n35 = x11 & x18 ;
  assign n36 = ~x12 & n35 ;
  assign n37 = n34 & ~n36 ;
  assign n38 = ~x2 & ~x3 ;
  assign n39 = ~x9 & ~x19 ;
  assign n40 = ~x0 & ~x1 ;
  assign n41 = n39 & n40 ;
  assign n42 = n38 & n41 ;
  assign n43 = ~x5 & x22 ;
  assign n44 = ~x6 & n43 ;
  assign n45 = ~x8 & n44 ;
  assign n46 = n42 & n45 ;
  assign n47 = n37 & n46 ;
  assign n48 = n47 ^ n33 ;
  assign n49 = x12 & ~x13 ;
  assign n50 = n49 ^ x10 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = ~x15 & x16 ;
  assign n53 = x13 & n52 ;
  assign n54 = ~x14 & n53 ;
  assign n55 = x12 & ~n54 ;
  assign n56 = n55 ^ n49 ;
  assign n57 = n51 & ~n56 ;
  assign n58 = n57 ^ n49 ;
  assign n59 = n58 ^ n33 ;
  assign n60 = ~n48 & ~n59 ;
  assign n61 = n60 ^ n57 ;
  assign n62 = n61 ^ n49 ;
  assign n63 = n62 ^ n47 ;
  assign n64 = ~n33 & n63 ;
  assign n65 = n64 ^ n33 ;
  assign y0 = ~n65 ;
endmodule
