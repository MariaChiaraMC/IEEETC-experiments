module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n9 = x5 ^ x0 ;
  assign n10 = x5 & n9 ;
  assign n11 = n10 ^ x5 ;
  assign n15 = x6 ^ x1 ;
  assign n12 = x6 ^ x2 ;
  assign n13 = n12 ^ x5 ;
  assign n14 = x2 & n13 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = n17 ^ x0 ;
  assign n20 = x7 ^ x6 ;
  assign n19 = n15 ^ x2 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = n15 & n21 ;
  assign n23 = n22 ^ x2 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n18 & n24 ;
  assign n26 = n25 ^ x6 ;
  assign n27 = n26 ^ x5 ;
  assign n28 = n27 ^ x0 ;
  assign n29 = n11 & n28 ;
  assign y0 = ~n29 ;
endmodule
