module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 ;
  assign n17 = x6 ^ x5 ;
  assign n18 = n17 ^ x7 ;
  assign n19 = x7 ^ x6 ;
  assign n20 = n19 ^ x7 ;
  assign n21 = x5 ^ x4 ;
  assign n22 = n21 ^ x6 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n20 & n23 ;
  assign n25 = n24 ^ n19 ;
  assign n26 = ~x8 & ~x9 ;
  assign n27 = x11 ^ x10 ;
  assign n28 = n26 & n27 ;
  assign n29 = ~n19 & n28 ;
  assign n30 = n29 ^ n18 ;
  assign n31 = ~n25 & ~n30 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = ~n18 & n32 ;
  assign n34 = n33 ^ n22 ;
  assign n35 = n34 ^ n18 ;
  assign n36 = x15 ^ x14 ;
  assign n37 = x13 ^ x12 ;
  assign n38 = ~n36 & ~n37 ;
  assign n39 = ~n35 & ~n38 ;
  assign n40 = x12 & ~x13 ;
  assign n41 = x10 & ~x11 ;
  assign n42 = n40 & n41 ;
  assign n43 = x14 & ~x15 ;
  assign n44 = x4 & x6 ;
  assign n45 = x5 & n44 ;
  assign n46 = n43 & n45 ;
  assign n47 = n42 & n46 ;
  assign n48 = ~n39 & ~n47 ;
  assign n49 = ~n40 & ~n43 ;
  assign n50 = x10 & n45 ;
  assign n51 = ~n49 & n50 ;
  assign n52 = ~x5 & x6 ;
  assign n53 = ~x4 & ~x10 ;
  assign n54 = n52 & n53 ;
  assign n55 = x4 & x7 ;
  assign n56 = x14 & x15 ;
  assign n57 = n55 & n56 ;
  assign n58 = n40 & n57 ;
  assign n59 = ~n54 & ~n58 ;
  assign n60 = ~n38 & ~n59 ;
  assign n61 = x5 & ~x6 ;
  assign n62 = ~x4 & x7 ;
  assign n63 = ~x13 & n43 ;
  assign n64 = ~x12 & n63 ;
  assign n65 = ~n62 & ~n64 ;
  assign n66 = n61 & ~n65 ;
  assign n67 = ~n60 & ~n66 ;
  assign n68 = ~n51 & n67 ;
  assign n69 = ~x11 & ~n68 ;
  assign n70 = ~x10 & x11 ;
  assign n71 = n37 & n56 ;
  assign n72 = x12 & x13 ;
  assign n73 = n36 & n72 ;
  assign n74 = ~n71 & ~n73 ;
  assign n75 = n45 & ~n74 ;
  assign n76 = n70 & n75 ;
  assign n77 = ~n69 & ~n76 ;
  assign n78 = x9 ^ x8 ;
  assign n79 = ~n77 & n78 ;
  assign n80 = n48 & ~n79 ;
  assign n81 = ~x0 & ~x3 ;
  assign n82 = ~x1 & n81 ;
  assign n83 = ~x2 & n82 ;
  assign n84 = ~n80 & n83 ;
  assign y0 = n84 ;
endmodule
