module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 ;
  assign n12 = ~x6 & ~x10 ;
  assign n13 = x3 & ~n12 ;
  assign n14 = x2 ^ x0 ;
  assign n15 = n14 ^ x9 ;
  assign n16 = x10 ^ x6 ;
  assign n17 = x2 & n16 ;
  assign n18 = n17 ^ x10 ;
  assign n19 = n15 & ~n18 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n20 ^ x10 ;
  assign n22 = n21 ^ x2 ;
  assign n23 = x9 & ~n22 ;
  assign n24 = ~n13 & ~n23 ;
  assign n25 = ~x8 & ~n24 ;
  assign n26 = ~x7 & n25 ;
  assign n30 = ~x7 & ~x9 ;
  assign n27 = x9 & x10 ;
  assign n28 = x3 & ~n27 ;
  assign n29 = ~x8 & ~n28 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = n32 ^ x6 ;
  assign n34 = x0 & ~n12 ;
  assign n35 = x0 & ~x3 ;
  assign n36 = x8 & ~n35 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = ~n34 & n37 ;
  assign n39 = n38 ^ n29 ;
  assign n40 = n39 ^ n34 ;
  assign n41 = ~n33 & ~n40 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = n42 ^ n34 ;
  assign n44 = ~x6 & ~n43 ;
  assign n45 = n44 ^ x6 ;
  assign n46 = ~n26 & n45 ;
  assign n47 = x4 & ~n46 ;
  assign n48 = ~x2 & ~x9 ;
  assign n49 = ~x5 & n48 ;
  assign n50 = ~x3 & n12 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = x1 & ~x7 ;
  assign n53 = n52 ^ x8 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = n52 ^ x7 ;
  assign n56 = n54 & n55 ;
  assign n57 = n56 ^ n52 ;
  assign n58 = n57 ^ n49 ;
  assign n59 = n51 & n58 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = n60 ^ n52 ;
  assign n62 = n61 ^ n50 ;
  assign n63 = n49 & n62 ;
  assign n64 = n63 ^ n49 ;
  assign n65 = ~n47 & ~n64 ;
  assign y0 = ~n65 ;
endmodule
