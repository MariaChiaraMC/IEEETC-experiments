module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 ;
  assign n16 = ~x10 & ~x11 ;
  assign n17 = ~x3 & x14 ;
  assign n18 = ~x9 & ~n17 ;
  assign n19 = ~x7 & ~x8 ;
  assign n20 = ~x4 & ~x5 ;
  assign n21 = ~x13 & n20 ;
  assign n22 = ~x0 & x9 ;
  assign n23 = x14 & ~n22 ;
  assign n24 = x6 & ~n23 ;
  assign n25 = n21 & n24 ;
  assign n26 = ~n19 & n25 ;
  assign n27 = ~n18 & ~n26 ;
  assign n28 = n16 & ~n27 ;
  assign n60 = x9 & ~x13 ;
  assign n82 = x7 & ~x14 ;
  assign n127 = ~n60 & ~n82 ;
  assign n128 = n16 & ~n127 ;
  assign n100 = x9 & ~x10 ;
  assign n130 = ~x13 & n100 ;
  assign n120 = ~x7 & x8 ;
  assign n129 = ~x5 & n120 ;
  assign n131 = n130 ^ n129 ;
  assign n132 = n131 ^ x14 ;
  assign n43 = x10 & x13 ;
  assign n44 = ~x11 & n43 ;
  assign n62 = ~x4 & ~x6 ;
  assign n136 = n44 & n62 ;
  assign n133 = x7 & ~x8 ;
  assign n134 = ~x3 & ~x6 ;
  assign n135 = ~n133 & n134 ;
  assign n137 = n136 ^ n135 ;
  assign n138 = n130 & n137 ;
  assign n139 = n138 ^ n136 ;
  assign n140 = n132 & n139 ;
  assign n141 = n140 ^ n138 ;
  assign n142 = n141 ^ n136 ;
  assign n143 = n142 ^ n130 ;
  assign n144 = x14 & n143 ;
  assign n145 = ~n128 & ~n144 ;
  assign n29 = x13 & ~x14 ;
  assign n30 = x4 & x7 ;
  assign n31 = ~x5 & n30 ;
  assign n32 = x1 & x3 ;
  assign n33 = n31 & n32 ;
  assign n34 = n29 & ~n33 ;
  assign n35 = ~x11 & n34 ;
  assign n36 = x5 & x6 ;
  assign n37 = x1 & x5 ;
  assign n38 = ~n36 & ~n37 ;
  assign n39 = ~x13 & x14 ;
  assign n40 = ~x0 & n39 ;
  assign n41 = ~n38 & n40 ;
  assign n42 = x5 & ~x7 ;
  assign n45 = ~x0 & ~x3 ;
  assign n46 = ~n36 & ~n45 ;
  assign n47 = n44 & ~n46 ;
  assign n48 = ~n42 & n47 ;
  assign n49 = ~n41 & ~n48 ;
  assign n50 = x4 & ~n49 ;
  assign n51 = x1 & x13 ;
  assign n52 = ~x10 & ~n51 ;
  assign n53 = ~n50 & ~n52 ;
  assign n54 = ~n35 & n53 ;
  assign n55 = ~x9 & ~n54 ;
  assign n81 = ~x5 & n62 ;
  assign n83 = x8 & n82 ;
  assign n84 = n81 & n83 ;
  assign n85 = x4 & x5 ;
  assign n86 = ~x9 & ~n85 ;
  assign n87 = ~n18 & ~n86 ;
  assign n88 = ~x0 & n87 ;
  assign n89 = ~n84 & ~n88 ;
  assign n90 = ~x6 & ~x8 ;
  assign n91 = x10 & n20 ;
  assign n92 = ~x0 & ~x7 ;
  assign n93 = n91 & n92 ;
  assign n94 = ~n90 & n93 ;
  assign n95 = x9 & ~n94 ;
  assign n96 = ~n89 & ~n95 ;
  assign n97 = ~x13 & n96 ;
  assign n56 = x10 & ~n31 ;
  assign n57 = x13 & n22 ;
  assign n58 = ~n56 & n57 ;
  assign n59 = ~n22 & n46 ;
  assign n61 = x14 & ~n60 ;
  assign n63 = n19 & n62 ;
  assign n64 = x10 & ~n63 ;
  assign n65 = ~n61 & n64 ;
  assign n66 = ~n59 & n65 ;
  assign n67 = x9 & ~x14 ;
  assign n68 = n67 ^ x4 ;
  assign n69 = n67 ^ n42 ;
  assign n70 = n69 ^ n42 ;
  assign n71 = ~x7 & ~x13 ;
  assign n72 = x6 & ~n71 ;
  assign n73 = ~x5 & ~n72 ;
  assign n74 = n73 ^ n42 ;
  assign n75 = n70 & n74 ;
  assign n76 = n75 ^ n42 ;
  assign n77 = n68 & n76 ;
  assign n78 = n77 ^ x4 ;
  assign n79 = n66 & n78 ;
  assign n80 = ~n58 & ~n79 ;
  assign n98 = n97 ^ n80 ;
  assign n99 = n98 ^ n80 ;
  assign n101 = ~x1 & x14 ;
  assign n102 = n101 ^ x13 ;
  assign n103 = x13 ^ x0 ;
  assign n104 = n103 ^ x14 ;
  assign n105 = n104 ^ x13 ;
  assign n106 = n105 ^ n100 ;
  assign n107 = n106 ^ x10 ;
  assign n108 = ~n102 & n107 ;
  assign n109 = n108 ^ x13 ;
  assign n110 = n100 & ~n109 ;
  assign n111 = n110 ^ n100 ;
  assign n112 = n111 ^ x10 ;
  assign n113 = n112 ^ n80 ;
  assign n114 = n113 ^ n80 ;
  assign n115 = ~n99 & n114 ;
  assign n116 = n115 ^ n80 ;
  assign n117 = x11 & n116 ;
  assign n118 = n117 ^ n80 ;
  assign n119 = ~n55 & n118 ;
  assign n146 = n145 ^ n119 ;
  assign n147 = n146 ^ n119 ;
  assign n121 = x6 & n120 ;
  assign n122 = ~x11 & ~n121 ;
  assign n123 = x13 & n100 ;
  assign n124 = ~n122 & n123 ;
  assign n125 = n124 ^ n119 ;
  assign n126 = n125 ^ n119 ;
  assign n148 = n147 ^ n126 ;
  assign n149 = x13 ^ x4 ;
  assign n150 = n149 ^ x4 ;
  assign n151 = ~x3 & ~x14 ;
  assign n152 = n31 & n151 ;
  assign n153 = n152 ^ x1 ;
  assign n154 = n153 ^ x4 ;
  assign n155 = ~n150 & n154 ;
  assign n156 = n155 ^ x1 ;
  assign n157 = n156 ^ n152 ;
  assign n158 = n157 ^ n150 ;
  assign n159 = x4 ^ x0 ;
  assign n160 = n159 ^ n149 ;
  assign n161 = n160 ^ n149 ;
  assign n162 = n161 ^ x4 ;
  assign n163 = n162 ^ n158 ;
  assign n164 = ~x2 & ~n38 ;
  assign n165 = n164 ^ x1 ;
  assign n166 = n162 ^ n150 ;
  assign n167 = n165 & ~n166 ;
  assign n168 = n167 ^ x1 ;
  assign n169 = n163 & n168 ;
  assign n170 = n169 ^ n150 ;
  assign n171 = n158 & ~n170 ;
  assign n172 = n171 ^ x13 ;
  assign n173 = x11 & ~n172 ;
  assign n174 = n81 & n133 ;
  assign n175 = n39 & n174 ;
  assign n176 = ~n173 & ~n175 ;
  assign n177 = n176 ^ x4 ;
  assign n178 = n177 ^ n176 ;
  assign n179 = n176 ^ x11 ;
  assign n180 = n179 ^ n176 ;
  assign n181 = n178 & ~n180 ;
  assign n182 = n181 ^ n176 ;
  assign n183 = ~x10 & ~n182 ;
  assign n184 = n183 ^ n176 ;
  assign n185 = ~x9 & ~n184 ;
  assign n186 = n185 ^ n119 ;
  assign n187 = n186 ^ n119 ;
  assign n188 = n187 ^ n147 ;
  assign n189 = n147 & ~n188 ;
  assign n190 = n189 ^ n147 ;
  assign n191 = ~n148 & n190 ;
  assign n192 = n191 ^ n189 ;
  assign n193 = n192 ^ n119 ;
  assign n194 = n193 ^ n147 ;
  assign n195 = x12 & n194 ;
  assign n196 = n195 ^ n119 ;
  assign n197 = ~n28 & n196 ;
  assign y0 = ~n197 ;
endmodule
