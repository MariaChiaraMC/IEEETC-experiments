module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 ;
  assign n33 = ~x25 & ~x31 ;
  assign n34 = ~x27 & ~x29 ;
  assign n35 = n33 & n34 ;
  assign n36 = ~x26 & ~x28 ;
  assign n37 = ~x24 & ~x30 ;
  assign n38 = n36 & n37 ;
  assign n39 = n35 & n38 ;
  assign n40 = ~x20 & ~x23 ;
  assign n41 = ~x17 & ~x18 ;
  assign n42 = n40 & n41 ;
  assign n43 = ~x16 & ~x19 ;
  assign n44 = ~x21 & ~x22 ;
  assign n45 = n43 & n44 ;
  assign n46 = n42 & n45 ;
  assign n47 = ~n39 & n46 ;
  assign n48 = ~x11 & ~x13 ;
  assign n49 = ~x9 & ~x15 ;
  assign n50 = ~x10 & ~x12 ;
  assign n51 = ~x8 & ~x14 ;
  assign n52 = n50 & n51 ;
  assign n53 = n49 & n52 ;
  assign n54 = n48 & n53 ;
  assign n55 = ~n47 & n54 ;
  assign y0 = ~n55 ;
endmodule
