module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 ;
  assign n8 = ~x4 & ~x5 ;
  assign n9 = n8 ^ x2 ;
  assign n10 = x2 ^ x1 ;
  assign n11 = n10 ^ x2 ;
  assign n12 = n11 ^ x2 ;
  assign n13 = n9 & ~n12 ;
  assign n14 = n13 ^ x2 ;
  assign n15 = ~x2 & x6 ;
  assign n16 = n15 ^ x3 ;
  assign n17 = ~n14 & ~n16 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = ~x3 & n18 ;
  assign n20 = n19 ^ n10 ;
  assign n21 = n20 ^ x3 ;
  assign n22 = x0 & n21 ;
  assign n24 = ~x1 & x2 ;
  assign n34 = x3 & n24 ;
  assign n25 = x4 & n24 ;
  assign n23 = x3 ^ x0 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n26 ^ x3 ;
  assign n35 = n34 ^ n27 ;
  assign n39 = n35 ^ n26 ;
  assign n40 = n39 ^ n23 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = n28 ^ n23 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = n26 ^ n8 ;
  assign n32 = n31 ^ n23 ;
  assign n33 = n30 & n32 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = n36 ^ n23 ;
  assign n38 = n29 & ~n37 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n41 ^ n29 ;
  assign n43 = x1 & ~x2 ;
  assign n44 = n43 ^ n23 ;
  assign n45 = n40 ^ n37 ;
  assign n46 = n45 ^ n29 ;
  assign n47 = ~n44 & ~n46 ;
  assign n48 = n47 ^ n23 ;
  assign n49 = n42 & n48 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = n50 ^ n23 ;
  assign n52 = n51 ^ x0 ;
  assign n53 = ~n22 & n52 ;
  assign y0 = ~n53 ;
endmodule
