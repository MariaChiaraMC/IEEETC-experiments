module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 ;
  assign n15 = x5 & x7 ;
  assign n16 = x8 & n15 ;
  assign n17 = ~x0 & ~x2 ;
  assign n18 = x3 & n17 ;
  assign n19 = ~x6 & n18 ;
  assign n20 = n16 & n19 ;
  assign n11 = x2 & x6 ;
  assign n21 = x0 & x5 ;
  assign n22 = n11 & n21 ;
  assign n23 = x3 & ~x8 ;
  assign n12 = ~x3 & x8 ;
  assign n24 = n23 ^ n12 ;
  assign n25 = x7 & n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n22 & n26 ;
  assign n28 = ~n20 & ~n27 ;
  assign n29 = ~x5 & ~x6 ;
  assign n30 = n29 ^ n17 ;
  assign n31 = ~x7 & x8 ;
  assign n32 = n31 ^ x3 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = n31 ^ x8 ;
  assign n35 = ~n33 & ~n34 ;
  assign n36 = n35 ^ n31 ;
  assign n37 = n36 ^ n17 ;
  assign n38 = n30 & n37 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n39 ^ n31 ;
  assign n41 = n40 ^ n29 ;
  assign n42 = n17 & n41 ;
  assign n43 = n42 ^ n17 ;
  assign n44 = n28 & ~n43 ;
  assign n13 = x7 & n12 ;
  assign n14 = n11 & n13 ;
  assign n45 = n44 ^ n14 ;
  assign n46 = n45 ^ n44 ;
  assign n47 = x0 & ~x5 ;
  assign n48 = n47 ^ n44 ;
  assign n49 = n48 ^ n44 ;
  assign n50 = n46 & n49 ;
  assign n51 = n50 ^ n44 ;
  assign n52 = ~x4 & ~n51 ;
  assign n53 = n52 ^ n44 ;
  assign n54 = x9 & ~n53 ;
  assign n55 = ~x3 & ~x4 ;
  assign n56 = x8 & n29 ;
  assign n57 = n55 & n56 ;
  assign n58 = ~x4 & ~x6 ;
  assign n59 = n23 & n58 ;
  assign n60 = x5 & n59 ;
  assign n61 = ~n57 & ~n60 ;
  assign n62 = ~x7 & ~x9 ;
  assign n63 = ~x2 & n62 ;
  assign n64 = ~n61 & n63 ;
  assign n65 = n11 & ~n55 ;
  assign n66 = ~n12 & n65 ;
  assign n67 = x5 & n62 ;
  assign n68 = ~n23 & n67 ;
  assign n69 = n66 & n68 ;
  assign n70 = ~n64 & ~n69 ;
  assign n71 = ~x2 & x7 ;
  assign n72 = n57 & n71 ;
  assign n85 = x6 & ~x7 ;
  assign n86 = ~n15 & ~n85 ;
  assign n87 = ~x8 & ~n29 ;
  assign n88 = n86 & n87 ;
  assign n89 = x2 & ~n88 ;
  assign n90 = x3 & ~n89 ;
  assign n73 = x5 & n31 ;
  assign n74 = ~x2 & ~x3 ;
  assign n75 = n73 & n74 ;
  assign n76 = ~x5 & x6 ;
  assign n77 = n71 ^ n23 ;
  assign n78 = n77 ^ n71 ;
  assign n79 = x2 & ~x7 ;
  assign n80 = n79 ^ n71 ;
  assign n81 = ~n78 & n80 ;
  assign n82 = n81 ^ n71 ;
  assign n83 = n76 & n82 ;
  assign n84 = ~n75 & ~n83 ;
  assign n91 = n90 ^ n84 ;
  assign n92 = n91 ^ n84 ;
  assign n93 = x6 & n73 ;
  assign n94 = ~x2 & ~n93 ;
  assign n95 = n94 ^ n84 ;
  assign n96 = n95 ^ n84 ;
  assign n97 = n92 & ~n96 ;
  assign n98 = n97 ^ n84 ;
  assign n99 = ~x4 & ~n98 ;
  assign n100 = n99 ^ n84 ;
  assign n101 = ~n72 & n100 ;
  assign n102 = x9 & ~n101 ;
  assign n103 = x3 & x4 ;
  assign n104 = x6 & ~x9 ;
  assign n105 = n103 & n104 ;
  assign n106 = n16 & n105 ;
  assign n107 = x4 & ~x7 ;
  assign n108 = ~x2 & n29 ;
  assign n109 = n107 & n108 ;
  assign n110 = n23 & n109 ;
  assign n111 = ~n106 & ~n110 ;
  assign n112 = ~n102 & n111 ;
  assign n113 = n70 & n112 ;
  assign n114 = ~x0 & ~n113 ;
  assign n115 = x4 & x6 ;
  assign n116 = ~x8 & x9 ;
  assign n117 = ~x2 & ~x7 ;
  assign n118 = ~x3 & x5 ;
  assign n119 = n117 & n118 ;
  assign n120 = n116 & n119 ;
  assign n121 = x2 & x3 ;
  assign n122 = x9 ^ x8 ;
  assign n123 = n15 ^ x9 ;
  assign n124 = n123 ^ n15 ;
  assign n125 = ~x5 & x7 ;
  assign n126 = n125 ^ n15 ;
  assign n127 = ~n124 & n126 ;
  assign n128 = n127 ^ n15 ;
  assign n129 = ~n122 & n128 ;
  assign n130 = n121 & n129 ;
  assign n131 = ~n120 & ~n130 ;
  assign n132 = n115 & ~n131 ;
  assign n133 = x4 ^ x3 ;
  assign n134 = x9 & n71 ;
  assign n135 = x9 ^ x4 ;
  assign n136 = n79 & n135 ;
  assign n137 = n136 ^ n133 ;
  assign n138 = n134 & n137 ;
  assign n139 = n138 ^ n136 ;
  assign n140 = n133 & n139 ;
  assign n141 = n76 & n140 ;
  assign n142 = x4 & ~x9 ;
  assign n143 = ~x4 & x9 ;
  assign n144 = ~n142 & ~n143 ;
  assign n145 = x2 & ~n115 ;
  assign n146 = n125 & n145 ;
  assign n147 = n144 & n146 ;
  assign n148 = x2 & ~x3 ;
  assign n149 = ~n142 & n148 ;
  assign n150 = n149 ^ x6 ;
  assign n151 = x7 ^ x4 ;
  assign n152 = n151 ^ x7 ;
  assign n153 = n67 ^ x7 ;
  assign n154 = ~n152 & n153 ;
  assign n155 = n154 ^ x7 ;
  assign n156 = n155 ^ n149 ;
  assign n157 = ~n150 & n156 ;
  assign n158 = n157 ^ n154 ;
  assign n159 = n158 ^ x7 ;
  assign n160 = n159 ^ x6 ;
  assign n161 = n149 & ~n160 ;
  assign n162 = n161 ^ n149 ;
  assign n163 = ~n147 & ~n162 ;
  assign n164 = ~n141 & n163 ;
  assign n165 = n164 ^ x8 ;
  assign n166 = n165 ^ n164 ;
  assign n167 = n166 ^ x0 ;
  assign n168 = x3 & ~x5 ;
  assign n169 = x9 & n168 ;
  assign n170 = ~x6 & x7 ;
  assign n171 = n170 ^ n85 ;
  assign n172 = ~x4 & n171 ;
  assign n173 = n172 ^ n85 ;
  assign n174 = n169 & n173 ;
  assign n175 = x5 & n105 ;
  assign n176 = n118 & n170 ;
  assign n177 = n144 & n176 ;
  assign n178 = ~n175 & ~n177 ;
  assign n179 = ~n174 & n178 ;
  assign n182 = n179 ^ x4 ;
  assign n183 = n182 ^ n179 ;
  assign n180 = n179 ^ x7 ;
  assign n181 = n180 ^ n179 ;
  assign n184 = n183 ^ n181 ;
  assign n185 = n168 ^ x9 ;
  assign n186 = n185 ^ n168 ;
  assign n187 = n168 ^ n118 ;
  assign n188 = n187 ^ n168 ;
  assign n189 = ~n186 & ~n188 ;
  assign n190 = n189 ^ n168 ;
  assign n191 = x6 & n190 ;
  assign n192 = n191 ^ n168 ;
  assign n193 = n192 ^ n179 ;
  assign n194 = n193 ^ n179 ;
  assign n195 = n194 ^ n183 ;
  assign n196 = ~n183 & ~n195 ;
  assign n197 = n196 ^ n183 ;
  assign n198 = n184 & ~n197 ;
  assign n199 = n198 ^ n196 ;
  assign n200 = n199 ^ n179 ;
  assign n201 = n200 ^ n183 ;
  assign n202 = x2 & n201 ;
  assign n203 = n202 ^ n179 ;
  assign n204 = x2 & x7 ;
  assign n205 = n142 & n204 ;
  assign n206 = n58 & n62 ;
  assign n207 = ~n205 & ~n206 ;
  assign n208 = n168 & ~n207 ;
  assign n209 = n208 ^ n203 ;
  assign n210 = n203 & ~n209 ;
  assign n211 = n210 ^ n164 ;
  assign n212 = n211 ^ n203 ;
  assign n213 = ~n167 & n212 ;
  assign n214 = n213 ^ n210 ;
  assign n215 = n214 ^ n203 ;
  assign n216 = x0 & n215 ;
  assign n217 = n216 ^ x0 ;
  assign n218 = ~n132 & ~n217 ;
  assign n219 = ~n114 & n218 ;
  assign n220 = n219 ^ x1 ;
  assign n221 = n220 ^ n219 ;
  assign n222 = ~x4 & n47 ;
  assign n223 = n85 & n222 ;
  assign n224 = x3 & n116 ;
  assign n225 = n223 & n224 ;
  assign n226 = x7 ^ x5 ;
  assign n227 = n116 & ~n226 ;
  assign n228 = x0 & ~n227 ;
  assign n229 = n15 ^ x8 ;
  assign n230 = n229 ^ n15 ;
  assign n231 = ~x0 & ~n125 ;
  assign n232 = n231 ^ n15 ;
  assign n233 = n232 ^ n15 ;
  assign n234 = ~n230 & ~n233 ;
  assign n235 = n234 ^ n15 ;
  assign n236 = x9 & n235 ;
  assign n237 = n236 ^ n15 ;
  assign n238 = ~x6 & n237 ;
  assign n239 = ~n228 & n238 ;
  assign n240 = ~x8 & ~x9 ;
  assign n241 = x6 & n21 ;
  assign n242 = n240 & n241 ;
  assign n243 = x7 & n242 ;
  assign n244 = ~n239 & ~n243 ;
  assign n245 = n103 & ~n244 ;
  assign n246 = ~x7 & x9 ;
  assign n247 = ~n55 & ~n246 ;
  assign n248 = ~n143 & ~n247 ;
  assign n249 = n241 & n248 ;
  assign n250 = ~x8 & n249 ;
  assign n251 = ~n245 & ~n250 ;
  assign n252 = ~n225 & n251 ;
  assign n253 = x2 & ~n252 ;
  assign n254 = ~x9 & n223 ;
  assign n255 = n143 ^ x0 ;
  assign n256 = n143 ^ n67 ;
  assign n257 = n256 ^ n67 ;
  assign n258 = n67 ^ n15 ;
  assign n259 = n257 & ~n258 ;
  assign n260 = n259 ^ n67 ;
  assign n261 = n255 & ~n260 ;
  assign n262 = n261 ^ x0 ;
  assign n263 = ~x6 & n262 ;
  assign n264 = ~n254 & ~n263 ;
  assign n265 = n74 & ~n264 ;
  assign n266 = n265 ^ x8 ;
  assign n267 = n266 ^ n265 ;
  assign n268 = ~x4 & n170 ;
  assign n269 = n18 & n268 ;
  assign n270 = x0 & x4 ;
  assign n271 = n148 & n270 ;
  assign n272 = n85 & n271 ;
  assign n273 = ~n269 & ~n272 ;
  assign n274 = ~x9 & ~n273 ;
  assign n275 = ~n58 & ~n270 ;
  assign n276 = ~x3 & ~n275 ;
  assign n277 = ~x2 & n115 ;
  assign n278 = n277 ^ x6 ;
  assign n279 = ~n55 & n278 ;
  assign n280 = n79 ^ x6 ;
  assign n281 = n103 ^ x2 ;
  assign n282 = n79 ^ x2 ;
  assign n283 = n282 ^ x2 ;
  assign n284 = ~n281 & n283 ;
  assign n285 = n284 ^ x2 ;
  assign n286 = n280 & n285 ;
  assign n287 = n286 ^ x6 ;
  assign n288 = ~n279 & n287 ;
  assign n289 = ~x9 & ~n11 ;
  assign n290 = x3 ^ x0 ;
  assign n291 = n290 ^ x3 ;
  assign n292 = x9 & ~n117 ;
  assign n293 = n292 ^ x3 ;
  assign n294 = n291 & ~n293 ;
  assign n295 = n294 ^ x3 ;
  assign n296 = ~n289 & ~n295 ;
  assign n297 = n288 & n296 ;
  assign n298 = ~n276 & n297 ;
  assign n299 = ~n274 & ~n298 ;
  assign n300 = x5 & ~n299 ;
  assign n301 = ~x3 & n142 ;
  assign n302 = x6 & n143 ;
  assign n303 = ~n301 & ~n302 ;
  assign n304 = n47 & n204 ;
  assign n305 = ~n303 & n304 ;
  assign n306 = ~x5 & ~x7 ;
  assign n307 = ~x6 & x9 ;
  assign n308 = n55 & n307 ;
  assign n309 = ~n105 & ~n308 ;
  assign n310 = n306 & ~n309 ;
  assign n311 = n17 & n310 ;
  assign n312 = ~n305 & ~n311 ;
  assign n313 = ~n300 & n312 ;
  assign n314 = n313 ^ n265 ;
  assign n315 = n267 & ~n314 ;
  assign n316 = n315 ^ n265 ;
  assign n317 = ~n253 & ~n316 ;
  assign n318 = n317 ^ n219 ;
  assign n319 = n221 & n318 ;
  assign n320 = n319 ^ n219 ;
  assign n321 = ~n54 & n320 ;
  assign y0 = ~n321 ;
endmodule
