module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 ;
  assign n13 = ~x5 & ~x6 ;
  assign n14 = ~x4 & ~n13 ;
  assign n9 = ~x4 & x5 ;
  assign n10 = x6 & n9 ;
  assign n11 = x2 & x7 ;
  assign n12 = n10 & n11 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = ~x2 & x3 ;
  assign n17 = n16 ^ n12 ;
  assign n18 = n12 ^ x0 ;
  assign n19 = ~n12 & ~n18 ;
  assign n20 = n19 ^ n12 ;
  assign n21 = ~n17 & ~n20 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ n12 ;
  assign n24 = n23 ^ x0 ;
  assign n25 = ~n15 & ~n24 ;
  assign n26 = n25 ^ n14 ;
  assign n27 = x1 & ~n26 ;
  assign y0 = ~n27 ;
endmodule
