module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n17 = x2 ^ x0 ;
  assign n18 = ~x10 & ~x11 ;
  assign n19 = ~x6 & ~x12 ;
  assign n20 = ~x4 & ~x13 ;
  assign n21 = n19 & n20 ;
  assign n22 = ~x3 & ~x15 ;
  assign n23 = x5 & x7 ;
  assign n24 = n22 & n23 ;
  assign n25 = ~x8 & ~x9 ;
  assign n26 = ~x14 & n25 ;
  assign n27 = n24 & n26 ;
  assign n28 = n21 & n27 ;
  assign n29 = n18 & n28 ;
  assign n30 = x1 & ~n29 ;
  assign n31 = ~x2 & n30 ;
  assign n32 = n17 & n31 ;
  assign n33 = n32 ^ n17 ;
  assign y0 = n33 ;
endmodule
