// Benchmark "./pla/newcwp.pla_dbb_orig_2NonExact" written by ABC on Fri Nov 20 10:25:43 2020

module \./pla/newcwp.pla_dbb_orig_2NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = ~x0;
endmodule


