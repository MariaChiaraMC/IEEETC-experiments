module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 ;
  assign n20 = ~x6 & x16 ;
  assign n21 = x7 & x8 ;
  assign n22 = n20 & n21 ;
  assign n23 = x4 ^ x3 ;
  assign n24 = ~x9 & n23 ;
  assign n25 = n24 ^ x3 ;
  assign n26 = n22 & n25 ;
  assign n27 = ~x3 & ~x10 ;
  assign n28 = x1 & n27 ;
  assign n29 = ~x16 & n28 ;
  assign n30 = ~n26 & ~n29 ;
  assign n31 = ~x17 & ~x18 ;
  assign n32 = ~n30 & n31 ;
  assign n33 = ~x7 & x17 ;
  assign n34 = ~x18 & ~n33 ;
  assign n35 = n25 & ~n34 ;
  assign n36 = x7 & ~x17 ;
  assign n37 = x16 ^ x6 ;
  assign n38 = ~n36 & ~n37 ;
  assign n39 = n33 ^ x18 ;
  assign n40 = ~x8 & n39 ;
  assign n41 = n40 ^ x18 ;
  assign n42 = n38 & ~n41 ;
  assign n43 = n35 & n42 ;
  assign n44 = ~n32 & ~n43 ;
  assign n45 = x3 & ~x9 ;
  assign n51 = x8 & x18 ;
  assign n46 = ~x6 & ~x7 ;
  assign n47 = ~x16 & n46 ;
  assign n48 = ~x17 & n47 ;
  assign n52 = n51 ^ n48 ;
  assign n60 = n52 ^ n48 ;
  assign n49 = ~n33 & ~n47 ;
  assign n50 = n49 ^ n48 ;
  assign n53 = n52 ^ n50 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = n54 ^ n48 ;
  assign n56 = n53 ^ n38 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = n55 & n58 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = n61 ^ n55 ;
  assign n63 = ~x8 & ~x18 ;
  assign n64 = n63 ^ n48 ;
  assign n65 = n59 ^ n55 ;
  assign n66 = ~n64 & n65 ;
  assign n67 = n66 ^ n48 ;
  assign n68 = n62 & ~n67 ;
  assign n69 = n68 ^ n48 ;
  assign n70 = n69 ^ n51 ;
  assign n71 = n70 ^ n48 ;
  assign n72 = n45 & n71 ;
  assign n73 = n44 & ~n72 ;
  assign y0 = ~n73 ;
endmodule
