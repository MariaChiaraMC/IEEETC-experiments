module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 ;
  assign n12 = x2 & ~x7 ;
  assign n13 = ~x2 & x7 ;
  assign n14 = ~n12 & ~n13 ;
  assign n9 = x0 & ~x1 ;
  assign n15 = x5 & n9 ;
  assign n16 = n14 & n15 ;
  assign n22 = x2 ^ x0 ;
  assign n23 = n22 ^ x7 ;
  assign n17 = x5 ^ x4 ;
  assign n19 = n17 ^ x5 ;
  assign n18 = n17 ^ x0 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = n20 ^ n19 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n24 ^ n17 ;
  assign n26 = n25 ^ n19 ;
  assign n27 = n26 ^ n17 ;
  assign n28 = n27 ^ n25 ;
  assign n30 = n23 ^ x1 ;
  assign n29 = n17 ^ x7 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = n32 ^ n26 ;
  assign n34 = n33 ^ n25 ;
  assign n35 = ~n28 & ~n34 ;
  assign n36 = n35 ^ n26 ;
  assign n37 = n36 ^ n25 ;
  assign n38 = n32 ^ n25 ;
  assign n39 = n23 ^ n17 ;
  assign n40 = n39 ^ n32 ;
  assign n41 = n40 ^ n25 ;
  assign n42 = ~n38 & n41 ;
  assign n43 = n42 ^ n23 ;
  assign n44 = n43 ^ n17 ;
  assign n45 = n44 ^ n26 ;
  assign n46 = n45 ^ n32 ;
  assign n47 = n46 ^ n25 ;
  assign n48 = n31 ^ n23 ;
  assign n49 = n48 ^ n17 ;
  assign n50 = n49 ^ n26 ;
  assign n51 = n50 ^ n32 ;
  assign n52 = ~n25 & ~n51 ;
  assign n53 = n52 ^ n31 ;
  assign n54 = n53 ^ n23 ;
  assign n55 = n54 ^ n32 ;
  assign n56 = n55 ^ n25 ;
  assign n57 = n47 & n56 ;
  assign n58 = n57 ^ n23 ;
  assign n59 = ~n37 & ~n58 ;
  assign n60 = ~n16 & ~n59 ;
  assign n10 = ~x4 & ~x5 ;
  assign n11 = n9 & n10 ;
  assign n61 = n60 ^ n11 ;
  assign n62 = x3 & ~n61 ;
  assign n63 = n62 ^ n60 ;
  assign y0 = ~n63 ;
endmodule
