module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 ;
  assign n11 = ~x5 & ~x6 ;
  assign n12 = ~x4 & n11 ;
  assign n13 = x3 ^ x2 ;
  assign n14 = ~x7 & ~x9 ;
  assign n15 = n14 ^ x3 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = x7 & x9 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = ~n16 & n18 ;
  assign n20 = n19 ^ n14 ;
  assign n21 = n13 & n20 ;
  assign n22 = n12 & n21 ;
  assign n23 = n22 ^ x1 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = x2 & ~x3 ;
  assign n26 = ~x7 & x9 ;
  assign n27 = n25 & n26 ;
  assign n28 = ~x2 & x3 ;
  assign n29 = n17 & n28 ;
  assign n30 = ~n27 & ~n29 ;
  assign n31 = x4 & x5 ;
  assign n32 = x6 & n31 ;
  assign n33 = ~n30 & n32 ;
  assign n34 = n33 ^ n22 ;
  assign n35 = ~n24 & n34 ;
  assign n36 = n35 ^ n22 ;
  assign n37 = ~x8 & n36 ;
  assign n38 = x8 & x9 ;
  assign n39 = x7 & n38 ;
  assign n40 = x1 & x2 ;
  assign n41 = ~x5 & x6 ;
  assign n42 = x3 & ~x4 ;
  assign n43 = n41 & n42 ;
  assign n44 = n40 & n43 ;
  assign n45 = n39 & n44 ;
  assign n46 = x9 & n42 ;
  assign n47 = ~x7 & n46 ;
  assign n48 = x6 & x8 ;
  assign n49 = ~x1 & ~n48 ;
  assign n50 = x5 & x8 ;
  assign n51 = n50 ^ n41 ;
  assign n52 = x2 & n51 ;
  assign n53 = n52 ^ n41 ;
  assign n54 = n49 & n53 ;
  assign n55 = n40 & n48 ;
  assign n56 = x5 & n55 ;
  assign n57 = ~n54 & ~n56 ;
  assign n58 = n47 & ~n57 ;
  assign n59 = ~x3 & ~x4 ;
  assign n60 = x1 & n59 ;
  assign n61 = ~x5 & ~x8 ;
  assign n62 = ~x6 & x8 ;
  assign n63 = ~x7 & n62 ;
  assign n64 = ~n61 & ~n63 ;
  assign n65 = ~x2 & ~n11 ;
  assign n66 = ~n64 & n65 ;
  assign n67 = n66 ^ x7 ;
  assign n68 = n67 ^ n66 ;
  assign n69 = x2 & n11 ;
  assign n70 = x8 & n69 ;
  assign n71 = n70 ^ n66 ;
  assign n72 = n71 ^ n66 ;
  assign n73 = ~n68 & n72 ;
  assign n74 = n73 ^ n66 ;
  assign n75 = ~x9 & n74 ;
  assign n76 = n75 ^ n66 ;
  assign n77 = n60 & n76 ;
  assign n78 = ~n58 & ~n77 ;
  assign n79 = ~x3 & x4 ;
  assign n80 = ~x2 & n79 ;
  assign n81 = x8 & ~x9 ;
  assign n82 = x5 & ~x6 ;
  assign n83 = n81 & n82 ;
  assign n84 = ~x8 & x9 ;
  assign n85 = n41 & n84 ;
  assign n86 = ~x1 & n85 ;
  assign n87 = ~n83 & ~n86 ;
  assign n88 = n80 & ~n87 ;
  assign n89 = ~x1 & x2 ;
  assign n90 = x6 & x9 ;
  assign n91 = n61 & ~n90 ;
  assign n92 = ~n83 & ~n91 ;
  assign n93 = n59 & ~n92 ;
  assign n94 = n89 & n93 ;
  assign n95 = x3 & x5 ;
  assign n96 = x9 ^ x6 ;
  assign n97 = n96 ^ x6 ;
  assign n102 = x4 & x8 ;
  assign n103 = n40 & n102 ;
  assign n104 = x1 & ~x2 ;
  assign n105 = ~x8 & n104 ;
  assign n106 = ~n103 & ~n105 ;
  assign n107 = n106 ^ x6 ;
  assign n108 = ~x6 & ~n107 ;
  assign n98 = x4 & n89 ;
  assign n99 = x9 ^ x8 ;
  assign n100 = n98 & n99 ;
  assign n111 = n108 ^ n100 ;
  assign n101 = n100 ^ n97 ;
  assign n109 = n108 ^ x6 ;
  assign n110 = ~n101 & ~n109 ;
  assign n112 = n111 ^ n110 ;
  assign n113 = ~n97 & n112 ;
  assign n114 = n113 ^ n108 ;
  assign n115 = n114 ^ n110 ;
  assign n116 = n95 & n115 ;
  assign n117 = ~n94 & ~n116 ;
  assign n118 = ~n88 & n117 ;
  assign n119 = n118 ^ x7 ;
  assign n120 = n119 ^ n118 ;
  assign n200 = ~x1 & ~x2 ;
  assign n190 = x1 & ~x9 ;
  assign n191 = x2 & n82 ;
  assign n192 = ~x2 & n41 ;
  assign n193 = ~n191 & ~n192 ;
  assign n194 = n190 & ~n193 ;
  assign n195 = ~x1 & x5 ;
  assign n196 = n90 & n195 ;
  assign n197 = ~n194 & ~n196 ;
  assign n201 = n200 ^ n197 ;
  assign n202 = n201 ^ n197 ;
  assign n198 = n197 ^ n11 ;
  assign n199 = n198 ^ n197 ;
  assign n203 = n202 ^ n199 ;
  assign n204 = n197 ^ x9 ;
  assign n205 = n204 ^ n197 ;
  assign n206 = n205 ^ n202 ;
  assign n207 = n202 & n206 ;
  assign n208 = n207 ^ n202 ;
  assign n209 = ~n203 & n208 ;
  assign n210 = n209 ^ n207 ;
  assign n211 = n210 ^ n197 ;
  assign n212 = n211 ^ n202 ;
  assign n213 = ~x8 & ~n212 ;
  assign n214 = n213 ^ n197 ;
  assign n152 = n25 & n41 ;
  assign n153 = n81 & n152 ;
  assign n121 = x5 ^ x2 ;
  assign n161 = n121 ^ x6 ;
  assign n154 = x6 ^ x1 ;
  assign n155 = n154 ^ x8 ;
  assign n156 = n155 ^ x5 ;
  assign n162 = n161 ^ n156 ;
  assign n163 = n162 ^ n156 ;
  assign n122 = n121 ^ x8 ;
  assign n157 = n156 ^ n122 ;
  assign n158 = n157 ^ n155 ;
  assign n159 = n158 ^ n121 ;
  assign n160 = n159 ^ n156 ;
  assign n164 = n163 ^ n160 ;
  assign n167 = n159 ^ n121 ;
  assign n165 = n155 ^ n121 ;
  assign n166 = n165 ^ n160 ;
  assign n168 = n167 ^ n166 ;
  assign n169 = n164 & ~n168 ;
  assign n170 = n169 ^ n159 ;
  assign n171 = n170 ^ n165 ;
  assign n172 = n171 ^ n167 ;
  assign n173 = n166 ^ n163 ;
  assign n174 = n170 & n173 ;
  assign n175 = n174 ^ n159 ;
  assign n176 = n175 ^ n160 ;
  assign n177 = n176 ^ n163 ;
  assign n178 = ~n172 & n177 ;
  assign n179 = n178 ^ x3 ;
  assign n180 = n179 ^ n178 ;
  assign n181 = x1 & n69 ;
  assign n182 = x6 & n105 ;
  assign n183 = ~n181 & ~n182 ;
  assign n184 = n183 ^ n178 ;
  assign n185 = ~n180 & ~n184 ;
  assign n186 = n185 ^ n178 ;
  assign n187 = x9 & n186 ;
  assign n188 = ~n153 & ~n187 ;
  assign n215 = n214 ^ n188 ;
  assign n139 = ~x5 & ~n89 ;
  assign n140 = n38 & n139 ;
  assign n123 = n122 ^ x9 ;
  assign n124 = x5 ^ x1 ;
  assign n125 = n124 ^ x8 ;
  assign n126 = n125 ^ n123 ;
  assign n127 = x9 ^ x5 ;
  assign n128 = n127 ^ x9 ;
  assign n129 = n99 ^ x9 ;
  assign n130 = n128 & n129 ;
  assign n131 = n130 ^ x9 ;
  assign n132 = n131 ^ n123 ;
  assign n133 = n126 & n132 ;
  assign n134 = n133 ^ n130 ;
  assign n135 = n134 ^ x9 ;
  assign n136 = n135 ^ n125 ;
  assign n137 = ~n123 & n136 ;
  assign n138 = n137 ^ n123 ;
  assign n141 = n140 ^ n138 ;
  assign n142 = n140 ^ n104 ;
  assign n143 = n140 ^ x6 ;
  assign n144 = n140 & ~n143 ;
  assign n145 = n144 ^ n140 ;
  assign n146 = n142 & n145 ;
  assign n147 = n146 ^ n144 ;
  assign n148 = n147 ^ n140 ;
  assign n149 = n148 ^ x6 ;
  assign n150 = ~n141 & ~n149 ;
  assign n151 = n150 ^ n140 ;
  assign n189 = n188 ^ n151 ;
  assign n216 = n215 ^ n189 ;
  assign n217 = n189 ^ x3 ;
  assign n218 = n217 ^ n189 ;
  assign n219 = ~n216 & n218 ;
  assign n220 = n219 ^ n189 ;
  assign n221 = x4 & ~n220 ;
  assign n222 = n221 ^ n188 ;
  assign n223 = n222 ^ n118 ;
  assign n224 = n120 & n223 ;
  assign n225 = n224 ^ n118 ;
  assign n226 = n78 & n225 ;
  assign n227 = n226 ^ x0 ;
  assign n228 = n227 ^ n226 ;
  assign n229 = ~x2 & ~x3 ;
  assign n230 = n82 & n229 ;
  assign n231 = n230 ^ x7 ;
  assign n232 = n231 ^ n230 ;
  assign n233 = x2 & x3 ;
  assign n234 = n41 & n233 ;
  assign n235 = n234 ^ n230 ;
  assign n236 = ~n232 & n235 ;
  assign n237 = n236 ^ n230 ;
  assign n238 = n84 & n237 ;
  assign n239 = ~x4 & n238 ;
  assign n240 = ~x8 & ~x9 ;
  assign n241 = ~x2 & x7 ;
  assign n242 = n59 & n241 ;
  assign n243 = ~x6 & n242 ;
  assign n244 = n240 & n243 ;
  assign n245 = x7 & ~x9 ;
  assign n246 = n82 & n245 ;
  assign n247 = n59 ^ x4 ;
  assign n248 = n247 ^ n59 ;
  assign n249 = n59 ^ x2 ;
  assign n250 = n249 ^ n59 ;
  assign n251 = n248 & ~n250 ;
  assign n252 = n251 ^ n59 ;
  assign n253 = x8 & n252 ;
  assign n254 = n253 ^ n59 ;
  assign n255 = n246 & n254 ;
  assign n256 = ~x4 & n14 ;
  assign n257 = ~x8 & n256 ;
  assign n258 = ~x7 & ~x8 ;
  assign n259 = x4 & ~n258 ;
  assign n260 = ~n38 & ~n245 ;
  assign n261 = n259 & n260 ;
  assign n262 = ~n257 & ~n261 ;
  assign n263 = n233 & ~n262 ;
  assign n264 = n47 ^ x8 ;
  assign n265 = n264 ^ n47 ;
  assign n266 = x9 ^ x7 ;
  assign n267 = n79 ^ x9 ;
  assign n268 = n267 ^ n79 ;
  assign n269 = n79 ^ n59 ;
  assign n270 = ~n268 & n269 ;
  assign n271 = n270 ^ n79 ;
  assign n272 = n266 & n271 ;
  assign n273 = n272 ^ n47 ;
  assign n274 = n265 & n273 ;
  assign n275 = n274 ^ n47 ;
  assign n276 = ~x2 & n275 ;
  assign n277 = ~n263 & ~n276 ;
  assign n278 = x6 & ~n277 ;
  assign n279 = n79 & n240 ;
  assign n280 = n46 & n62 ;
  assign n281 = ~n279 & ~n280 ;
  assign n282 = x2 & ~n281 ;
  assign n283 = ~x6 & n28 ;
  assign n284 = n240 & n283 ;
  assign n285 = x4 & n284 ;
  assign n286 = ~n282 & ~n285 ;
  assign n287 = ~x7 & ~n286 ;
  assign n288 = ~n278 & ~n287 ;
  assign n289 = n288 ^ x5 ;
  assign n290 = n289 ^ n288 ;
  assign n291 = ~x6 & ~x8 ;
  assign n292 = ~n48 & ~n291 ;
  assign n293 = n25 & ~n292 ;
  assign n294 = ~n283 & ~n293 ;
  assign n295 = n102 & n283 ;
  assign n296 = x9 & n295 ;
  assign n297 = ~n256 & ~n296 ;
  assign n298 = ~n294 & ~n297 ;
  assign n299 = ~x3 & ~n258 ;
  assign n300 = n90 & ~n299 ;
  assign n301 = n79 ^ x4 ;
  assign n302 = ~x2 & ~n301 ;
  assign n303 = n302 ^ x4 ;
  assign n304 = n300 & ~n303 ;
  assign n305 = ~n298 & ~n304 ;
  assign n306 = n305 ^ n288 ;
  assign n307 = ~n290 & n306 ;
  assign n308 = n307 ^ n288 ;
  assign n309 = ~n255 & n308 ;
  assign n310 = ~n244 & n309 ;
  assign n311 = n310 ^ x1 ;
  assign n312 = n311 ^ n310 ;
  assign n322 = ~x5 & ~n81 ;
  assign n323 = ~n50 & n241 ;
  assign n324 = ~n322 & n323 ;
  assign n313 = n26 ^ x6 ;
  assign n314 = n313 ^ n70 ;
  assign n315 = n314 ^ n26 ;
  assign n325 = n324 ^ n315 ;
  assign n329 = n325 ^ n314 ;
  assign n330 = n329 ^ n313 ;
  assign n316 = n315 ^ n314 ;
  assign n317 = n316 ^ n313 ;
  assign n318 = n317 ^ n313 ;
  assign n319 = n314 ^ x2 ;
  assign n320 = n319 ^ n313 ;
  assign n321 = ~n318 & n320 ;
  assign n326 = n325 ^ n321 ;
  assign n327 = n326 ^ n313 ;
  assign n328 = ~n317 & n327 ;
  assign n331 = n330 ^ n328 ;
  assign n332 = n331 ^ n317 ;
  assign n333 = n50 & ~n245 ;
  assign n334 = n333 ^ n313 ;
  assign n335 = n330 ^ n327 ;
  assign n336 = n335 ^ n317 ;
  assign n337 = ~n334 & n336 ;
  assign n338 = n337 ^ n313 ;
  assign n339 = n332 & n338 ;
  assign n340 = n339 ^ n337 ;
  assign n341 = n340 ^ n313 ;
  assign n342 = n341 ^ x6 ;
  assign n343 = n42 & n342 ;
  assign n344 = ~x5 & n81 ;
  assign n345 = ~n84 & ~n344 ;
  assign n346 = n243 & ~n345 ;
  assign n347 = x3 & x4 ;
  assign n348 = n82 & n347 ;
  assign n349 = ~x9 & n258 ;
  assign n350 = ~n39 & ~n349 ;
  assign n351 = n350 ^ x7 ;
  assign n352 = n351 ^ n350 ;
  assign n353 = n350 ^ n240 ;
  assign n354 = n353 ^ n350 ;
  assign n355 = n352 & n354 ;
  assign n356 = n355 ^ n350 ;
  assign n357 = ~x2 & ~n356 ;
  assign n358 = n357 ^ n350 ;
  assign n359 = n348 & ~n358 ;
  assign n362 = n291 ^ n85 ;
  assign n363 = n362 ^ n85 ;
  assign n360 = n85 ^ x5 ;
  assign n361 = n360 ^ n85 ;
  assign n364 = n363 ^ n361 ;
  assign n365 = ~n81 & ~n90 ;
  assign n366 = n365 ^ n85 ;
  assign n367 = n366 ^ n85 ;
  assign n368 = n367 ^ n363 ;
  assign n369 = ~n363 & ~n368 ;
  assign n370 = n369 ^ n363 ;
  assign n371 = ~n364 & ~n370 ;
  assign n372 = n371 ^ n369 ;
  assign n373 = n372 ^ n85 ;
  assign n374 = n373 ^ n363 ;
  assign n375 = x4 & ~n374 ;
  assign n376 = n375 ^ n85 ;
  assign n377 = n229 & n376 ;
  assign n378 = ~x7 & n377 ;
  assign n379 = ~n359 & ~n378 ;
  assign n380 = ~n346 & n379 ;
  assign n381 = ~n343 & n380 ;
  assign n382 = n381 ^ n310 ;
  assign n383 = ~n312 & n382 ;
  assign n384 = n383 ^ n310 ;
  assign n385 = ~n239 & n384 ;
  assign n386 = n385 ^ n226 ;
  assign n387 = n228 & n386 ;
  assign n388 = n387 ^ n226 ;
  assign n389 = ~n45 & n388 ;
  assign n390 = ~n37 & n389 ;
  assign y0 = ~n390 ;
endmodule
