module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n15 = ~x10 & ~x11 ;
  assign n16 = ~x9 & n15 ;
  assign n17 = ~x12 & n16 ;
  assign n18 = x0 & ~n17 ;
  assign n19 = ~x2 & ~x3 ;
  assign n20 = ~n18 & n19 ;
  assign n21 = ~x1 & n20 ;
  assign n22 = x5 & ~n21 ;
  assign n23 = x4 & x7 ;
  assign n24 = ~x5 & ~x8 ;
  assign n25 = n23 & ~n24 ;
  assign n26 = x13 & n25 ;
  assign n27 = ~x6 & n26 ;
  assign n28 = ~n22 & n27 ;
  assign y0 = n28 ;
endmodule
