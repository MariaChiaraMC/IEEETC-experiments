module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 ;
  assign n11 = x5 & ~x8 ;
  assign n12 = n11 ^ x8 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n13 ^ x7 ;
  assign n15 = x0 & ~x1 ;
  assign n16 = ~x2 & ~x3 ;
  assign n17 = n15 & ~n16 ;
  assign n18 = n17 ^ n11 ;
  assign n19 = n18 ^ x9 ;
  assign n20 = x9 & ~n19 ;
  assign n21 = n20 ^ n11 ;
  assign n22 = n21 ^ x9 ;
  assign n23 = n14 & ~n22 ;
  assign n24 = n23 ^ n20 ;
  assign n25 = n24 ^ x9 ;
  assign n26 = ~x7 & n25 ;
  assign n27 = n26 ^ n11 ;
  assign n28 = x6 & n27 ;
  assign n29 = ~x2 & x4 ;
  assign n30 = x3 & n15 ;
  assign n31 = ~x6 & n30 ;
  assign n32 = ~x8 & ~n31 ;
  assign n33 = ~n29 & ~n32 ;
  assign n36 = x3 ^ x0 ;
  assign n37 = n36 ^ x3 ;
  assign n34 = x3 ^ x2 ;
  assign n35 = n34 ^ x3 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = x1 & ~x6 ;
  assign n40 = n39 ^ x3 ;
  assign n41 = n40 ^ x3 ;
  assign n42 = n41 ^ n37 ;
  assign n43 = ~n37 & ~n42 ;
  assign n44 = n43 ^ n37 ;
  assign n45 = n38 & ~n44 ;
  assign n46 = n45 ^ n43 ;
  assign n47 = n46 ^ x3 ;
  assign n48 = n47 ^ n37 ;
  assign n49 = ~x8 & ~n48 ;
  assign n50 = n49 ^ x3 ;
  assign n51 = ~n33 & ~n50 ;
  assign n52 = ~x7 & ~n51 ;
  assign n53 = ~x5 & n52 ;
  assign n54 = ~n28 & ~n53 ;
  assign y0 = ~n54 ;
endmodule
