module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n9 = ~x4 & ~x5 ;
  assign n10 = x6 & x7 ;
  assign n11 = n9 & ~n10 ;
  assign n12 = x2 & ~n11 ;
  assign n13 = x2 & x3 ;
  assign n14 = x1 & ~n13 ;
  assign n15 = x0 & n14 ;
  assign n16 = ~n12 & n15 ;
  assign n17 = n9 ^ x2 ;
  assign n18 = n17 ^ n9 ;
  assign n19 = ~x7 & n9 ;
  assign n20 = ~x6 & n19 ;
  assign n21 = n20 ^ n9 ;
  assign n22 = n18 & n21 ;
  assign n23 = n22 ^ n9 ;
  assign n24 = x3 & ~n23 ;
  assign n25 = n24 ^ x2 ;
  assign n26 = n25 ^ x0 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = x5 & n13 ;
  assign n29 = x4 & n28 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = n27 & n30 ;
  assign n32 = n31 ^ n25 ;
  assign n33 = ~x1 & n32 ;
  assign n34 = ~n16 & ~n33 ;
  assign y0 = ~n34 ;
endmodule
