module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ;
  assign n15 = x11 ^ x10 ;
  assign n21 = n15 ^ x12 ;
  assign n16 = n15 ^ x13 ;
  assign n23 = n21 ^ n16 ;
  assign n19 = x10 ^ x9 ;
  assign n17 = n16 ^ x11 ;
  assign n18 = n17 ^ n15 ;
  assign n20 = n19 ^ n18 ;
  assign n22 = n21 ^ n20 ;
  assign n24 = n23 ^ n22 ;
  assign n27 = n20 ^ n19 ;
  assign n25 = n19 ^ n15 ;
  assign n26 = n25 ^ n22 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = ~n24 & n28 ;
  assign n30 = n29 ^ n20 ;
  assign n31 = n30 ^ n25 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = n26 ^ n23 ;
  assign n34 = n30 & n33 ;
  assign n35 = n34 ^ n20 ;
  assign n36 = n35 ^ n22 ;
  assign n37 = n36 ^ n23 ;
  assign n38 = ~n32 & ~n37 ;
  assign n39 = n38 ^ x9 ;
  assign y0 = ~n39 ;
endmodule
