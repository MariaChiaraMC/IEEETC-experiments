module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 ;
  assign n9 = ~x1 & ~x3 ;
  assign n10 = ~x6 & ~x7 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = ~x2 & x4 ;
  assign n13 = n12 ^ x5 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = x0 & ~x4 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = ~n14 & n16 ;
  assign n18 = n17 ^ n12 ;
  assign n19 = n18 ^ n9 ;
  assign n20 = n11 & n19 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n21 ^ n12 ;
  assign n23 = n22 ^ n10 ;
  assign n24 = n9 & n23 ;
  assign n25 = n24 ^ n9 ;
  assign y0 = n25 ;
endmodule
