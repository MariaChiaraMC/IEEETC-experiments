module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 ;
  output y0 ;
  wire n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 ;
  assign n23 = x1 & ~x2 ;
  assign n24 = ~x0 & n23 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = x0 & ~x1 ;
  assign n28 = ~x2 & ~x3 ;
  assign n29 = n27 & ~n28 ;
  assign n30 = n29 ^ x3 ;
  assign n31 = x5 & n30 ;
  assign n32 = n31 ^ x3 ;
  assign n33 = ~n26 & ~n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n34 ^ x3 ;
  assign n36 = n35 ^ x5 ;
  assign n37 = ~x4 & ~n36 ;
  assign n206 = ~x19 & ~x20 ;
  assign n38 = ~x1 & x2 ;
  assign n39 = ~x6 & ~x7 ;
  assign n40 = ~x13 & ~n39 ;
  assign n41 = x8 & ~x13 ;
  assign n42 = ~x9 & ~n41 ;
  assign n43 = ~n40 & n42 ;
  assign n44 = ~x8 & ~x15 ;
  assign n45 = x9 & ~x12 ;
  assign n46 = ~n44 & n45 ;
  assign n47 = x8 ^ x6 ;
  assign n48 = x7 & ~n47 ;
  assign n49 = n48 ^ x6 ;
  assign n50 = x11 & ~n49 ;
  assign n51 = ~n46 & ~n50 ;
  assign n52 = ~n43 & n51 ;
  assign n53 = x10 & ~n52 ;
  assign n54 = x11 & x16 ;
  assign n55 = x12 & ~n54 ;
  assign n56 = x9 & x11 ;
  assign n57 = n44 & ~n56 ;
  assign n58 = ~x6 & n57 ;
  assign n59 = ~n55 & n58 ;
  assign n60 = x13 & ~n59 ;
  assign n61 = x8 & ~x10 ;
  assign n62 = x16 & ~n61 ;
  assign n63 = ~x8 & ~x11 ;
  assign n64 = n39 & ~n63 ;
  assign n65 = ~n62 & n64 ;
  assign n66 = x12 & ~x13 ;
  assign n67 = n66 ^ x7 ;
  assign n68 = n67 ^ x17 ;
  assign n69 = n56 ^ x6 ;
  assign n70 = ~x7 & n69 ;
  assign n71 = n70 ^ n56 ;
  assign n72 = ~n68 & ~n71 ;
  assign n73 = n72 ^ n70 ;
  assign n74 = n73 ^ n56 ;
  assign n75 = n74 ^ x7 ;
  assign n76 = ~x17 & n75 ;
  assign n77 = ~n65 & n76 ;
  assign n78 = ~n60 & n77 ;
  assign n79 = ~n53 & n78 ;
  assign n80 = n38 & ~n79 ;
  assign n81 = ~x12 & x13 ;
  assign n82 = x10 & ~x12 ;
  assign n83 = n56 & n82 ;
  assign n84 = ~n81 & ~n83 ;
  assign n85 = ~x2 & ~n84 ;
  assign n86 = n23 ^ x0 ;
  assign n87 = n23 ^ x13 ;
  assign n88 = n23 ^ x4 ;
  assign n89 = n23 & n88 ;
  assign n90 = n89 ^ n23 ;
  assign n91 = n87 & n90 ;
  assign n92 = n91 ^ n89 ;
  assign n93 = n92 ^ n23 ;
  assign n94 = n93 ^ x4 ;
  assign n95 = ~n86 & n94 ;
  assign n96 = ~n85 & n95 ;
  assign n97 = x10 & ~x11 ;
  assign n98 = ~x8 & x9 ;
  assign n99 = ~n97 & n98 ;
  assign n100 = x12 ^ x11 ;
  assign n101 = n100 ^ x13 ;
  assign n102 = x13 ^ x12 ;
  assign n103 = n102 ^ n99 ;
  assign n104 = ~n101 & n103 ;
  assign n105 = n104 ^ x12 ;
  assign n106 = x7 & ~x12 ;
  assign n107 = n106 ^ n99 ;
  assign n108 = ~n105 & ~n107 ;
  assign n109 = n108 ^ n106 ;
  assign n110 = ~n99 & n109 ;
  assign n111 = n110 ^ n104 ;
  assign n112 = n111 ^ x12 ;
  assign n113 = ~x1 & ~n112 ;
  assign n114 = n96 & ~n113 ;
  assign n115 = ~n80 & n114 ;
  assign n116 = x5 & ~n115 ;
  assign n117 = x1 & n39 ;
  assign n118 = ~x12 & ~x13 ;
  assign n119 = x9 & n118 ;
  assign n120 = n63 & n119 ;
  assign n121 = n117 & n120 ;
  assign n122 = x2 & ~n121 ;
  assign n123 = ~x4 & ~n122 ;
  assign n124 = ~x0 & n123 ;
  assign n125 = ~x10 & x11 ;
  assign n126 = ~x4 & n117 ;
  assign n127 = n119 & n126 ;
  assign n128 = n125 & n127 ;
  assign n129 = n128 ^ x8 ;
  assign n130 = n129 ^ n128 ;
  assign n131 = ~x9 & n125 ;
  assign n132 = n39 & n118 ;
  assign n133 = n97 & n132 ;
  assign n134 = ~n131 & ~n133 ;
  assign n135 = n27 & ~n134 ;
  assign n136 = ~x9 & n97 ;
  assign n137 = n118 & n126 ;
  assign n138 = n136 & n137 ;
  assign n139 = ~n135 & ~n138 ;
  assign n140 = n139 ^ n128 ;
  assign n141 = ~n130 & ~n140 ;
  assign n142 = n141 ^ n128 ;
  assign n143 = x2 & n142 ;
  assign n144 = ~n124 & ~n143 ;
  assign n145 = ~n116 & n144 ;
  assign n146 = ~x3 & ~n145 ;
  assign n147 = ~x4 & ~n66 ;
  assign n148 = ~n40 & n147 ;
  assign n149 = x5 & ~x8 ;
  assign n150 = n149 ^ x13 ;
  assign n151 = n150 ^ n131 ;
  assign n152 = n151 ^ n149 ;
  assign n153 = n152 ^ n151 ;
  assign n154 = n63 ^ n24 ;
  assign n155 = n154 ^ x9 ;
  assign n157 = x11 & n61 ;
  assign n156 = x2 & x5 ;
  assign n158 = n157 ^ n156 ;
  assign n159 = n63 & ~n158 ;
  assign n160 = n159 ^ n157 ;
  assign n161 = n155 & n160 ;
  assign n162 = n161 ^ n159 ;
  assign n163 = n162 ^ n157 ;
  assign n164 = n163 ^ n63 ;
  assign n165 = x9 & n164 ;
  assign n166 = n165 ^ n151 ;
  assign n167 = n166 ^ n150 ;
  assign n168 = n153 & ~n167 ;
  assign n169 = n168 ^ n165 ;
  assign n170 = ~n136 & ~n165 ;
  assign n171 = n170 ^ n150 ;
  assign n172 = ~n169 & n171 ;
  assign n173 = n172 ^ n170 ;
  assign n174 = n150 & n173 ;
  assign n175 = n174 ^ n168 ;
  assign n176 = n175 ^ x13 ;
  assign n177 = n176 ^ n165 ;
  assign n178 = n148 & n177 ;
  assign n179 = x1 ^ x0 ;
  assign n180 = n179 ^ x3 ;
  assign n181 = x1 & n180 ;
  assign n182 = n180 ^ x2 ;
  assign n183 = x3 & ~x21 ;
  assign n184 = n183 ^ n181 ;
  assign n185 = n182 & n184 ;
  assign n186 = n185 ^ n183 ;
  assign n187 = n181 & n186 ;
  assign n188 = n187 ^ n179 ;
  assign n189 = x4 & n188 ;
  assign n190 = x2 & n39 ;
  assign n191 = n27 & n190 ;
  assign n192 = n157 & n191 ;
  assign n193 = n119 & n192 ;
  assign n194 = ~n189 & ~n193 ;
  assign n195 = n194 ^ x3 ;
  assign n196 = n195 ^ n194 ;
  assign n197 = n194 ^ x1 ;
  assign n198 = n197 ^ x2 ;
  assign n199 = n198 ^ n194 ;
  assign n200 = n196 & ~n199 ;
  assign n201 = n200 ^ n194 ;
  assign n202 = x5 & ~n201 ;
  assign n203 = n202 ^ n194 ;
  assign n204 = ~n178 & n203 ;
  assign n205 = ~n146 & n204 ;
  assign n207 = n206 ^ n205 ;
  assign n208 = n207 ^ n205 ;
  assign n209 = n205 ^ x18 ;
  assign n210 = ~n208 & n209 ;
  assign n211 = n210 ^ n205 ;
  assign n212 = ~n37 & n211 ;
  assign n213 = x14 & ~n212 ;
  assign y0 = n213 ;
endmodule
