module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 ;
  assign n11 = x3 & ~x9 ;
  assign n12 = x4 & ~n11 ;
  assign n13 = ~x5 & ~x9 ;
  assign n14 = ~x1 & x3 ;
  assign n15 = ~n13 & ~n14 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = x7 & x9 ;
  assign n18 = n17 ^ x0 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = n17 ^ x7 ;
  assign n21 = n19 & ~n20 ;
  assign n22 = n21 ^ n17 ;
  assign n23 = n22 ^ n12 ;
  assign n24 = n16 & ~n23 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ n17 ;
  assign n27 = n26 ^ n15 ;
  assign n28 = ~n12 & ~n27 ;
  assign n29 = n28 ^ n12 ;
  assign n30 = x8 & ~n29 ;
  assign n31 = x9 ^ x6 ;
  assign n32 = x9 ^ x5 ;
  assign n33 = n32 ^ x5 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = x3 & ~x4 ;
  assign n36 = ~x1 & ~x5 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = ~n35 & n37 ;
  assign n39 = n38 ^ x5 ;
  assign n40 = n39 ^ n35 ;
  assign n41 = n34 & n40 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = n42 ^ n35 ;
  assign n44 = ~n31 & ~n43 ;
  assign n45 = n30 & n44 ;
  assign n46 = ~x5 & x9 ;
  assign n47 = n35 & n46 ;
  assign n48 = ~x6 & ~x9 ;
  assign n49 = x3 & ~n48 ;
  assign n50 = ~x4 & x9 ;
  assign n51 = x4 & ~x9 ;
  assign n52 = ~n50 & ~n51 ;
  assign n53 = x6 & x9 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = x5 & n54 ;
  assign n56 = ~n49 & n55 ;
  assign n57 = ~n47 & ~n56 ;
  assign n58 = x1 & ~x8 ;
  assign n59 = ~n57 & n58 ;
  assign n60 = x4 ^ x3 ;
  assign n61 = ~x6 & n36 ;
  assign n62 = ~x8 & ~x9 ;
  assign n63 = n61 & n62 ;
  assign n64 = n63 ^ x4 ;
  assign n65 = n64 ^ n63 ;
  assign n66 = n65 ^ n60 ;
  assign n67 = ~x6 & x8 ;
  assign n68 = x9 & ~n67 ;
  assign n69 = ~x1 & x5 ;
  assign n70 = ~n48 & n69 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = ~n68 & ~n71 ;
  assign n73 = n72 ^ n63 ;
  assign n74 = n73 ^ n68 ;
  assign n75 = ~n66 & ~n74 ;
  assign n76 = n75 ^ n72 ;
  assign n77 = n76 ^ n68 ;
  assign n78 = n60 & ~n77 ;
  assign n79 = ~n59 & ~n78 ;
  assign n80 = x0 & n79 ;
  assign n81 = x1 & x3 ;
  assign n82 = x4 & x5 ;
  assign n83 = x6 & ~x9 ;
  assign n84 = x8 & n83 ;
  assign n85 = n82 & n84 ;
  assign n86 = ~x4 & ~x6 ;
  assign n87 = n46 & n86 ;
  assign n88 = ~n85 & ~n87 ;
  assign n89 = n81 & ~n88 ;
  assign n90 = ~x0 & ~n89 ;
  assign n91 = ~x1 & ~x6 ;
  assign n92 = x4 & ~x5 ;
  assign n93 = ~x8 & n92 ;
  assign n94 = ~x4 & ~x9 ;
  assign n95 = x5 & x8 ;
  assign n96 = ~x5 & ~x8 ;
  assign n97 = ~n95 & ~n96 ;
  assign n98 = n94 & n97 ;
  assign n99 = ~n93 & ~n98 ;
  assign n100 = n91 & ~n99 ;
  assign n101 = n100 ^ x3 ;
  assign n102 = n101 ^ n100 ;
  assign n103 = n102 ^ n90 ;
  assign n105 = x1 & x6 ;
  assign n106 = n105 ^ x5 ;
  assign n104 = n91 ^ x8 ;
  assign n107 = n106 ^ n104 ;
  assign n108 = n107 ^ x9 ;
  assign n109 = n105 ^ n91 ;
  assign n110 = n91 & n109 ;
  assign n111 = n110 ^ n104 ;
  assign n112 = n111 ^ n91 ;
  assign n113 = n108 & n112 ;
  assign n114 = n113 ^ n110 ;
  assign n115 = n114 ^ n91 ;
  assign n116 = x9 & n115 ;
  assign n117 = ~n63 & ~n116 ;
  assign n118 = n117 ^ x4 ;
  assign n119 = ~x4 & n118 ;
  assign n120 = n119 ^ n100 ;
  assign n121 = n120 ^ x4 ;
  assign n122 = ~n103 & ~n121 ;
  assign n123 = n122 ^ n119 ;
  assign n124 = n123 ^ x4 ;
  assign n125 = n90 & ~n124 ;
  assign n126 = n125 ^ n90 ;
  assign n127 = ~x7 & ~n126 ;
  assign n128 = ~n80 & n127 ;
  assign n131 = x8 & ~x9 ;
  assign n132 = ~x3 & n131 ;
  assign n133 = ~x6 & n132 ;
  assign n129 = x3 & ~x8 ;
  assign n130 = n53 & n129 ;
  assign n134 = n133 ^ n130 ;
  assign n135 = ~x0 & n134 ;
  assign n136 = n135 ^ n133 ;
  assign n137 = n82 & n136 ;
  assign n138 = x1 & n137 ;
  assign n139 = x4 & x6 ;
  assign n140 = ~x8 & n139 ;
  assign n141 = ~x4 & x8 ;
  assign n142 = ~n140 & ~n141 ;
  assign n143 = x3 & ~n142 ;
  assign n144 = n46 & n143 ;
  assign n145 = ~x5 & x6 ;
  assign n146 = n132 & n145 ;
  assign n147 = n87 ^ x8 ;
  assign n148 = n147 ^ n87 ;
  assign n149 = n148 ^ n146 ;
  assign n150 = n92 ^ n83 ;
  assign n151 = n92 & n150 ;
  assign n152 = n151 ^ n87 ;
  assign n153 = n152 ^ n92 ;
  assign n154 = ~n149 & n153 ;
  assign n155 = n154 ^ n151 ;
  assign n156 = n155 ^ n92 ;
  assign n157 = ~n146 & n156 ;
  assign n158 = n157 ^ n146 ;
  assign n159 = ~n144 & ~n158 ;
  assign n160 = x5 & ~x8 ;
  assign n161 = n160 ^ x9 ;
  assign n162 = n35 ^ x6 ;
  assign n163 = n162 ^ n35 ;
  assign n164 = ~x3 & x4 ;
  assign n165 = n164 ^ n35 ;
  assign n166 = ~n163 & n165 ;
  assign n167 = n166 ^ n35 ;
  assign n168 = n167 ^ n160 ;
  assign n169 = n161 & n168 ;
  assign n170 = n169 ^ n166 ;
  assign n171 = n170 ^ n35 ;
  assign n172 = n171 ^ x9 ;
  assign n173 = n160 & n172 ;
  assign n174 = n173 ^ n160 ;
  assign n175 = ~x1 & ~n174 ;
  assign n176 = n159 & n175 ;
  assign n177 = ~n48 & n164 ;
  assign n178 = ~n132 & ~n177 ;
  assign n179 = x6 & ~n62 ;
  assign n180 = ~n178 & ~n179 ;
  assign n181 = n35 & n84 ;
  assign n182 = ~n180 & ~n181 ;
  assign n183 = ~x5 & ~n182 ;
  assign n184 = n67 & n164 ;
  assign n185 = x1 & ~n184 ;
  assign n186 = ~n183 & n185 ;
  assign n187 = ~n176 & ~n186 ;
  assign n188 = n187 ^ x0 ;
  assign n189 = n188 ^ n187 ;
  assign n190 = n189 ^ x7 ;
  assign n191 = ~x3 & x9 ;
  assign n192 = x8 ^ x6 ;
  assign n193 = x6 ^ x4 ;
  assign n194 = n193 ^ n192 ;
  assign n195 = n69 ^ x8 ;
  assign n196 = n195 ^ n69 ;
  assign n197 = x1 & x5 ;
  assign n198 = n197 ^ n69 ;
  assign n199 = n196 & ~n198 ;
  assign n200 = n199 ^ n69 ;
  assign n201 = n200 ^ n192 ;
  assign n202 = ~n194 & ~n201 ;
  assign n203 = n202 ^ n199 ;
  assign n204 = n203 ^ n69 ;
  assign n205 = n204 ^ n193 ;
  assign n206 = n192 & n205 ;
  assign n207 = n206 ^ n192 ;
  assign n208 = n191 & n207 ;
  assign n209 = ~x8 & ~n11 ;
  assign n210 = n209 ^ n81 ;
  assign n211 = n210 ^ n81 ;
  assign n212 = n81 ^ n36 ;
  assign n213 = n212 ^ n81 ;
  assign n214 = ~n211 & n213 ;
  assign n215 = n214 ^ n81 ;
  assign n216 = ~n131 & n215 ;
  assign n217 = n216 ^ n81 ;
  assign n218 = n139 & n217 ;
  assign n219 = ~n208 & ~n218 ;
  assign n220 = x9 & n160 ;
  assign n221 = ~x6 & n220 ;
  assign n222 = n13 & n67 ;
  assign n223 = ~n221 & ~n222 ;
  assign n224 = n35 & ~n223 ;
  assign n225 = x1 & n224 ;
  assign n226 = n219 & ~n225 ;
  assign n227 = ~n86 & ~n140 ;
  assign n228 = x5 & ~x9 ;
  assign n229 = ~x1 & ~x3 ;
  assign n230 = n228 & n229 ;
  assign n231 = ~n227 & n230 ;
  assign n232 = n231 ^ n226 ;
  assign n233 = n226 & ~n232 ;
  assign n234 = n233 ^ n187 ;
  assign n235 = n234 ^ n226 ;
  assign n236 = n190 & ~n235 ;
  assign n237 = n236 ^ n233 ;
  assign n238 = n237 ^ n226 ;
  assign n239 = x7 & n238 ;
  assign n240 = n239 ^ x7 ;
  assign n241 = ~n138 & ~n240 ;
  assign n242 = ~n128 & n241 ;
  assign n243 = n242 ^ x2 ;
  assign n244 = n243 ^ n242 ;
  assign n245 = n244 ^ n45 ;
  assign n246 = n14 & n50 ;
  assign n247 = ~x9 & n164 ;
  assign n248 = ~n246 & ~n247 ;
  assign n249 = x0 & x7 ;
  assign n250 = n145 & n249 ;
  assign n251 = ~n248 & n250 ;
  assign n252 = x3 & x5 ;
  assign n253 = n83 & ~n252 ;
  assign n254 = ~x0 & ~x1 ;
  assign n255 = ~x4 & ~x7 ;
  assign n256 = n254 & n255 ;
  assign n257 = n253 & n256 ;
  assign n258 = ~x6 & x7 ;
  assign n259 = ~x0 & n258 ;
  assign n260 = n47 & n259 ;
  assign n261 = ~n257 & ~n260 ;
  assign n262 = ~n251 & n261 ;
  assign n263 = n262 ^ x5 ;
  assign n264 = ~x6 & ~x7 ;
  assign n265 = x6 & x7 ;
  assign n266 = ~n264 & ~n265 ;
  assign n267 = x4 & x9 ;
  assign n268 = ~n266 & n267 ;
  assign n269 = n81 & n268 ;
  assign n270 = n229 & n266 ;
  assign n271 = x9 & n270 ;
  assign n272 = ~n86 & n271 ;
  assign n273 = ~n269 & ~n272 ;
  assign n274 = n273 ^ x0 ;
  assign n275 = n274 ^ n273 ;
  assign n276 = n105 & n191 ;
  assign n277 = n255 & n276 ;
  assign n278 = ~x3 & ~x4 ;
  assign n279 = ~x1 & x7 ;
  assign n280 = ~n278 & n279 ;
  assign n281 = n48 ^ x3 ;
  assign n282 = n281 ^ n48 ;
  assign n283 = n52 & ~n86 ;
  assign n284 = n283 ^ n48 ;
  assign n285 = n282 & n284 ;
  assign n286 = n285 ^ n48 ;
  assign n287 = n280 & n286 ;
  assign n288 = ~n277 & ~n287 ;
  assign n289 = n288 ^ n273 ;
  assign n290 = ~n275 & n289 ;
  assign n291 = n290 ^ n273 ;
  assign n292 = n291 ^ n262 ;
  assign n293 = n263 & ~n292 ;
  assign n294 = n293 ^ n290 ;
  assign n295 = n294 ^ n273 ;
  assign n296 = n295 ^ x5 ;
  assign n297 = n262 & ~n296 ;
  assign n298 = n297 ^ n262 ;
  assign n299 = n298 ^ n262 ;
  assign n300 = ~x8 & n299 ;
  assign n301 = ~x1 & x6 ;
  assign n302 = x0 & n301 ;
  assign n303 = n82 & n302 ;
  assign n304 = n17 & n303 ;
  assign n305 = x8 & ~n304 ;
  assign n362 = ~x0 & x5 ;
  assign n363 = n362 ^ x6 ;
  assign n364 = n363 ^ x9 ;
  assign n365 = n364 ^ x9 ;
  assign n366 = n365 ^ n362 ;
  assign n378 = n366 ^ n362 ;
  assign n367 = x9 ^ x4 ;
  assign n368 = n367 ^ x9 ;
  assign n379 = n368 ^ n362 ;
  assign n369 = n368 ^ x9 ;
  assign n380 = n379 ^ n369 ;
  assign n381 = ~n378 & ~n380 ;
  assign n371 = n362 ^ x0 ;
  assign n372 = n371 ^ n362 ;
  assign n373 = n362 ^ n92 ;
  assign n374 = n373 ^ n362 ;
  assign n375 = n372 & ~n374 ;
  assign n382 = n381 ^ n375 ;
  assign n370 = n369 ^ n366 ;
  assign n376 = n375 ^ n362 ;
  assign n377 = ~n370 & n376 ;
  assign n383 = n382 ^ n377 ;
  assign n384 = ~n366 & n383 ;
  assign n385 = n384 ^ n381 ;
  assign n386 = n385 ^ n362 ;
  assign n387 = n386 ^ n362 ;
  assign n388 = x1 & n387 ;
  assign n389 = x7 & ~n388 ;
  assign n390 = ~n303 & n389 ;
  assign n323 = n17 & n61 ;
  assign n324 = n197 ^ x7 ;
  assign n325 = n324 ^ x9 ;
  assign n326 = n197 ^ x6 ;
  assign n327 = n326 ^ x6 ;
  assign n328 = ~n36 & ~n91 ;
  assign n329 = n328 ^ x6 ;
  assign n330 = ~n327 & ~n329 ;
  assign n331 = n330 ^ x6 ;
  assign n332 = n331 ^ n324 ;
  assign n333 = n325 & n332 ;
  assign n334 = n333 ^ n330 ;
  assign n335 = n334 ^ x6 ;
  assign n336 = n335 ^ x9 ;
  assign n337 = ~n324 & n336 ;
  assign n338 = n337 ^ n324 ;
  assign n339 = ~n323 & n338 ;
  assign n340 = ~x4 & ~n339 ;
  assign n306 = n48 & n279 ;
  assign n307 = n228 ^ n46 ;
  assign n308 = n307 ^ x1 ;
  assign n309 = n46 ^ x6 ;
  assign n310 = n46 ^ x7 ;
  assign n311 = n310 ^ n309 ;
  assign n312 = n309 & n311 ;
  assign n313 = n312 ^ n46 ;
  assign n314 = n313 ^ n309 ;
  assign n315 = n308 & n314 ;
  assign n316 = n315 ^ n312 ;
  assign n317 = n316 ^ n309 ;
  assign n318 = x1 & n317 ;
  assign n319 = ~n306 & ~n318 ;
  assign n320 = ~x4 & ~n319 ;
  assign n321 = n36 & n268 ;
  assign n322 = ~n320 & ~n321 ;
  assign n341 = n340 ^ n322 ;
  assign n342 = n341 ^ n322 ;
  assign n343 = n82 ^ x9 ;
  assign n344 = n264 ^ x1 ;
  assign n345 = n344 ^ n264 ;
  assign n346 = n266 ^ n264 ;
  assign n347 = n345 & n346 ;
  assign n348 = n347 ^ n264 ;
  assign n349 = n348 ^ n82 ;
  assign n350 = n343 & n349 ;
  assign n351 = n350 ^ n347 ;
  assign n352 = n351 ^ n264 ;
  assign n353 = n352 ^ x9 ;
  assign n354 = n82 & n353 ;
  assign n355 = n354 ^ n82 ;
  assign n356 = n355 ^ n322 ;
  assign n357 = n356 ^ n322 ;
  assign n358 = ~n342 & ~n357 ;
  assign n359 = n358 ^ n322 ;
  assign n360 = x0 & n359 ;
  assign n361 = n360 ^ n322 ;
  assign n391 = n390 ^ n361 ;
  assign n392 = n391 ^ n361 ;
  assign n401 = ~x9 & n82 ;
  assign n393 = n52 ^ n46 ;
  assign n394 = n393 ^ n46 ;
  assign n395 = n46 ^ x5 ;
  assign n396 = n395 ^ n46 ;
  assign n397 = ~n394 & n396 ;
  assign n398 = n397 ^ n46 ;
  assign n399 = x1 & n398 ;
  assign n400 = n399 ^ n46 ;
  assign n402 = n401 ^ n400 ;
  assign n403 = n402 ^ n400 ;
  assign n404 = n400 ^ x1 ;
  assign n405 = n404 ^ n400 ;
  assign n406 = n403 & ~n405 ;
  assign n407 = n406 ^ n400 ;
  assign n408 = ~x0 & n407 ;
  assign n409 = n408 ^ n400 ;
  assign n410 = x6 & n409 ;
  assign n411 = ~x0 & ~n36 ;
  assign n412 = ~n32 & n411 ;
  assign n413 = n86 & n412 ;
  assign n414 = ~x7 & ~n413 ;
  assign n415 = ~n410 & n414 ;
  assign n416 = n415 ^ n361 ;
  assign n417 = n416 ^ n361 ;
  assign n418 = ~n392 & ~n417 ;
  assign n419 = n418 ^ n361 ;
  assign n420 = x3 & ~n419 ;
  assign n421 = n420 ^ n361 ;
  assign n422 = n305 & n421 ;
  assign n423 = n422 ^ n300 ;
  assign n424 = ~n300 & n423 ;
  assign n425 = n424 ^ n242 ;
  assign n426 = n425 ^ n300 ;
  assign n427 = ~n245 & n426 ;
  assign n428 = n427 ^ n424 ;
  assign n429 = n428 ^ n300 ;
  assign n430 = ~n45 & ~n429 ;
  assign n431 = n430 ^ n45 ;
  assign y0 = n431 ;
endmodule
