module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 ;
  assign n9 = ~x4 & x6 ;
  assign n10 = ~x3 & n9 ;
  assign n11 = ~x2 & ~n10 ;
  assign n12 = x1 & ~n11 ;
  assign n13 = ~x6 & ~x7 ;
  assign n14 = ~x3 & n13 ;
  assign n15 = x3 & ~x4 ;
  assign n16 = ~n14 & ~n15 ;
  assign n17 = x2 & ~n16 ;
  assign n21 = x3 & x4 ;
  assign n22 = x1 & n21 ;
  assign n18 = ~x2 & ~x3 ;
  assign n19 = n18 ^ x7 ;
  assign n20 = n19 ^ n18 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ n19 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n9 & n26 ;
  assign n28 = n27 ^ n22 ;
  assign n29 = ~x4 & ~x6 ;
  assign n30 = n29 ^ n22 ;
  assign n31 = n25 & ~n30 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = n32 ^ n25 ;
  assign n34 = ~n28 & n33 ;
  assign n35 = n24 & n34 ;
  assign n36 = n35 ^ n27 ;
  assign n37 = n36 ^ x7 ;
  assign n38 = x3 ^ x2 ;
  assign n39 = n38 ^ n29 ;
  assign n40 = n39 ^ x3 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = x4 & x6 ;
  assign n43 = n41 ^ n38 ;
  assign n44 = n43 ^ n41 ;
  assign n45 = ~n42 & ~n44 ;
  assign n46 = n45 ^ n39 ;
  assign n47 = n39 ^ n13 ;
  assign n48 = ~n43 & n47 ;
  assign n49 = n48 ^ n41 ;
  assign n50 = n49 ^ n43 ;
  assign n51 = n46 & ~n50 ;
  assign n52 = n41 & n51 ;
  assign n53 = n52 ^ n45 ;
  assign n54 = n53 ^ x2 ;
  assign n56 = n54 ^ n13 ;
  assign n55 = n54 ^ n42 ;
  assign n57 = n56 ^ n55 ;
  assign n58 = n56 ^ x3 ;
  assign n59 = n58 ^ n56 ;
  assign n60 = n57 & n59 ;
  assign n61 = n60 ^ n56 ;
  assign n62 = x1 & ~n61 ;
  assign n63 = n62 ^ n54 ;
  assign n64 = ~n37 & n63 ;
  assign n65 = ~n17 & n64 ;
  assign n66 = n65 ^ x5 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = x4 & ~x7 ;
  assign n69 = ~x2 & ~n68 ;
  assign n70 = x6 & ~n69 ;
  assign n71 = x1 & x4 ;
  assign n72 = ~n70 & ~n71 ;
  assign n73 = ~x3 & ~n72 ;
  assign n75 = x4 ^ x3 ;
  assign n74 = x7 ^ x3 ;
  assign n76 = n75 ^ n74 ;
  assign n77 = n76 ^ n75 ;
  assign n78 = ~x2 & n42 ;
  assign n80 = n78 ^ x3 ;
  assign n79 = n78 ^ x6 ;
  assign n81 = n80 ^ n79 ;
  assign n82 = n81 ^ n75 ;
  assign n83 = n82 ^ n77 ;
  assign n84 = n79 ^ x3 ;
  assign n85 = n84 ^ n77 ;
  assign n86 = ~n79 & n85 ;
  assign n87 = n86 ^ n75 ;
  assign n88 = ~n83 & n87 ;
  assign n89 = n88 ^ n86 ;
  assign n90 = n89 ^ n75 ;
  assign n91 = n90 ^ n79 ;
  assign n92 = ~n77 & ~n91 ;
  assign n93 = n92 ^ n86 ;
  assign n94 = n93 ^ n79 ;
  assign n95 = n94 ^ x6 ;
  assign n96 = ~x1 & n95 ;
  assign n97 = x2 & n21 ;
  assign n98 = ~x6 & n97 ;
  assign n99 = ~n96 & ~n98 ;
  assign n100 = ~n73 & n99 ;
  assign n101 = n100 ^ n65 ;
  assign n102 = ~n67 & n101 ;
  assign n103 = n102 ^ n65 ;
  assign n104 = ~n12 & n103 ;
  assign n105 = ~x0 & ~n104 ;
  assign y0 = n105 ;
endmodule
