// Benchmark "./pla/t2.pla_res_11NonExact" written by ABC on Fri Nov 20 10:31:25 2020

module \./pla/t2.pla_res_11NonExact  ( 
    x0, x1, x2, x3, x4, x5,
    z0  );
  input  x0, x1, x2, x3, x4, x5;
  output z0;
  wire new_n8_, new_n9_, new_n10_, new_n11_, new_n12_, new_n13_, new_n14_,
    new_n15_;
  assign new_n8_ = x3 & x4;
  assign new_n9_ = x5 & new_n8_;
  assign new_n10_ = ~x2 & ~new_n9_;
  assign new_n11_ = x2 & x3;
  assign new_n12_ = ~x4 & ~x5;
  assign new_n13_ = new_n11_ & ~new_n12_;
  assign new_n14_ = ~x0 & x1;
  assign new_n15_ = ~new_n13_ & new_n14_;
  assign z0 = ~new_n10_ & new_n15_;
endmodule


