// Benchmark "./pla/x2dn.pla_dbb_orig_24NonExact" written by ABC on Fri Nov 20 10:30:32 2020

module \./pla/x2dn.pla_dbb_orig_24NonExact  ( 
    x0, x1,
    z0  );
  input  x0, x1;
  output z0;
  assign z0 = ~x0 & ~x1;
endmodule


