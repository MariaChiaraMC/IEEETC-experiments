// Benchmark "./t4.pla" written by ABC on Thu Apr 23 11:00:06 2020

module \./t4.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11,
    z7  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11;
  output z7;
  assign z7 = 1'b1;
endmodule


