module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 ;
  assign n11 = x0 & ~x3 ;
  assign n12 = ~x7 & ~x8 ;
  assign n13 = x8 & ~x9 ;
  assign n14 = ~n12 & ~n13 ;
  assign n15 = x7 & x9 ;
  assign n16 = ~x6 & ~n15 ;
  assign n17 = n14 & n16 ;
  assign n18 = ~x4 & n17 ;
  assign n19 = x6 & ~x9 ;
  assign n20 = ~x8 & n19 ;
  assign n21 = ~x7 & n20 ;
  assign n22 = ~n18 & ~n21 ;
  assign n23 = n11 & ~n22 ;
  assign n24 = ~x0 & ~x4 ;
  assign n25 = x7 & n13 ;
  assign n26 = ~x3 & x6 ;
  assign n27 = n25 & n26 ;
  assign n28 = x3 & x9 ;
  assign n29 = x8 ^ x7 ;
  assign n30 = x8 ^ x6 ;
  assign n31 = ~n29 & ~n30 ;
  assign n32 = n28 & n31 ;
  assign n33 = ~n27 & ~n32 ;
  assign n34 = n24 & ~n33 ;
  assign n35 = x0 & x6 ;
  assign n36 = x7 & x8 ;
  assign n37 = x3 & x4 ;
  assign n38 = n36 & n37 ;
  assign n39 = n35 & n38 ;
  assign n40 = ~n34 & ~n39 ;
  assign n41 = ~n23 & n40 ;
  assign n42 = ~x0 & x4 ;
  assign n43 = x6 & x7 ;
  assign n44 = ~x8 & x9 ;
  assign n45 = n43 & n44 ;
  assign n46 = ~x6 & n25 ;
  assign n47 = ~n45 & ~n46 ;
  assign n48 = n42 & ~n47 ;
  assign n49 = ~x3 & n48 ;
  assign n50 = x5 & ~n49 ;
  assign n51 = n41 & n50 ;
  assign n52 = x0 & x7 ;
  assign n53 = x9 ^ x8 ;
  assign n54 = x4 ^ x3 ;
  assign n55 = x9 ^ x4 ;
  assign n56 = n55 ^ x4 ;
  assign n57 = ~n54 & ~n56 ;
  assign n58 = n57 ^ x4 ;
  assign n59 = ~n53 & ~n58 ;
  assign n60 = n52 & n59 ;
  assign n61 = x4 & ~x7 ;
  assign n62 = ~n13 & n61 ;
  assign n63 = x3 & x8 ;
  assign n64 = n63 ^ x0 ;
  assign n65 = n62 & ~n64 ;
  assign n66 = ~n60 & ~n65 ;
  assign n67 = ~x6 & ~n66 ;
  assign n68 = n13 & n26 ;
  assign n69 = n61 & n68 ;
  assign n70 = ~x5 & ~n69 ;
  assign n71 = ~n67 & n70 ;
  assign n72 = ~x6 & x9 ;
  assign n73 = ~n19 & ~n72 ;
  assign n74 = ~x7 & x8 ;
  assign n75 = ~x0 & n74 ;
  assign n76 = ~x4 & n75 ;
  assign n77 = n76 ^ x3 ;
  assign n78 = n77 ^ n76 ;
  assign n79 = ~x8 & n52 ;
  assign n80 = n79 ^ n76 ;
  assign n81 = ~n78 & n80 ;
  assign n82 = n81 ^ n76 ;
  assign n83 = ~n73 & n82 ;
  assign n84 = n71 & ~n83 ;
  assign n85 = ~n51 & ~n84 ;
  assign n86 = n42 ^ n12 ;
  assign n87 = ~x3 & ~x6 ;
  assign n88 = n87 ^ x9 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = x3 & x6 ;
  assign n91 = n90 ^ n87 ;
  assign n92 = n89 & n91 ;
  assign n93 = n92 ^ n87 ;
  assign n94 = n93 ^ n42 ;
  assign n95 = n86 & n94 ;
  assign n96 = n95 ^ n92 ;
  assign n97 = n96 ^ n87 ;
  assign n98 = n97 ^ n12 ;
  assign n99 = n42 & n98 ;
  assign n100 = n99 ^ n42 ;
  assign n101 = ~n85 & ~n100 ;
  assign n102 = ~x1 & n101 ;
  assign n103 = ~x3 & x5 ;
  assign n104 = n19 & n103 ;
  assign n105 = n76 & n104 ;
  assign n106 = x0 & ~x5 ;
  assign n107 = n74 & n87 ;
  assign n108 = n106 & n107 ;
  assign n109 = x1 & ~n108 ;
  assign n110 = ~x8 & ~x9 ;
  assign n111 = n110 ^ n24 ;
  assign n112 = x5 & x7 ;
  assign n113 = n112 ^ x6 ;
  assign n114 = n113 ^ x6 ;
  assign n115 = n87 ^ x6 ;
  assign n116 = ~n114 & n115 ;
  assign n117 = n116 ^ x6 ;
  assign n118 = n117 ^ n110 ;
  assign n119 = n111 & n118 ;
  assign n120 = n119 ^ n116 ;
  assign n121 = n120 ^ x6 ;
  assign n122 = n121 ^ n24 ;
  assign n123 = n110 & n122 ;
  assign n124 = n123 ^ n110 ;
  assign n125 = n109 & ~n124 ;
  assign n126 = ~n105 & n125 ;
  assign n127 = ~x5 & ~x9 ;
  assign n132 = x6 & ~x8 ;
  assign n133 = n24 & n132 ;
  assign n134 = ~x5 & ~n133 ;
  assign n128 = ~n12 & ~n36 ;
  assign n129 = n42 & ~n128 ;
  assign n130 = n19 & n129 ;
  assign n131 = x5 & ~n130 ;
  assign n135 = n134 ^ n131 ;
  assign n136 = n131 ^ x4 ;
  assign n137 = n136 ^ n135 ;
  assign n141 = ~x6 & ~x7 ;
  assign n142 = n110 & n141 ;
  assign n143 = x8 & x9 ;
  assign n144 = n43 & n143 ;
  assign n145 = ~n142 & ~n144 ;
  assign n146 = x0 & ~n145 ;
  assign n147 = n72 & n128 ;
  assign n148 = ~n52 & n147 ;
  assign n149 = ~n146 & ~n148 ;
  assign n138 = n35 ^ x0 ;
  assign n139 = ~n74 & ~n138 ;
  assign n140 = n139 ^ x0 ;
  assign n150 = n149 ^ n140 ;
  assign n151 = x4 & n150 ;
  assign n152 = n151 ^ n149 ;
  assign n153 = n137 & n152 ;
  assign n154 = n153 ^ n151 ;
  assign n155 = n154 ^ n149 ;
  assign n156 = n155 ^ x4 ;
  assign n157 = n135 & n156 ;
  assign n158 = n157 ^ n134 ;
  assign n159 = ~n127 & ~n158 ;
  assign n160 = n159 ^ x3 ;
  assign n161 = n160 ^ n159 ;
  assign n162 = x0 & x5 ;
  assign n163 = ~x6 & x8 ;
  assign n164 = ~x4 & n163 ;
  assign n165 = ~n20 & ~n164 ;
  assign n166 = n162 & ~n165 ;
  assign n167 = ~x0 & x8 ;
  assign n168 = x9 ^ x6 ;
  assign n169 = x5 ^ x4 ;
  assign n170 = x9 ^ x5 ;
  assign n171 = n170 ^ x5 ;
  assign n172 = n169 & n171 ;
  assign n173 = n172 ^ x5 ;
  assign n174 = n168 & ~n173 ;
  assign n175 = n167 & n174 ;
  assign n176 = ~n166 & ~n175 ;
  assign n177 = x7 & ~n176 ;
  assign n178 = n177 ^ n159 ;
  assign n179 = ~n161 & n178 ;
  assign n180 = n179 ^ n159 ;
  assign n181 = n126 & ~n180 ;
  assign n182 = ~n102 & ~n181 ;
  assign n183 = x3 & ~x6 ;
  assign n184 = n52 & n183 ;
  assign n185 = ~x4 & ~x5 ;
  assign n186 = n184 & n185 ;
  assign n187 = n110 & n186 ;
  assign n188 = ~n182 & ~n187 ;
  assign n189 = ~x2 & ~n188 ;
  assign n190 = n43 & n110 ;
  assign n191 = ~x1 & n162 ;
  assign n192 = n190 & n191 ;
  assign n193 = n37 & n192 ;
  assign n194 = ~x0 & ~x1 ;
  assign n195 = n37 & n194 ;
  assign n196 = n12 & n72 ;
  assign n197 = n195 & n196 ;
  assign n198 = ~x9 & n183 ;
  assign n199 = x1 & x4 ;
  assign n200 = x7 & n167 ;
  assign n201 = n199 & n200 ;
  assign n202 = n198 & n201 ;
  assign n203 = ~n197 & ~n202 ;
  assign n204 = ~x5 & ~n203 ;
  assign n205 = ~x4 & n11 ;
  assign n206 = x8 ^ x1 ;
  assign n207 = n141 ^ n43 ;
  assign n208 = n141 ^ x8 ;
  assign n209 = n208 ^ n141 ;
  assign n210 = n207 & ~n209 ;
  assign n211 = n210 ^ n141 ;
  assign n212 = ~n206 & n211 ;
  assign n213 = n205 & n212 ;
  assign n214 = n127 & n213 ;
  assign n215 = ~n204 & ~n214 ;
  assign n216 = ~n193 & n215 ;
  assign n217 = x1 & x8 ;
  assign n218 = n106 & n217 ;
  assign n219 = x5 & ~x8 ;
  assign n220 = n194 & n219 ;
  assign n221 = ~n218 & ~n220 ;
  assign n222 = ~x3 & ~x7 ;
  assign n223 = x6 & x9 ;
  assign n224 = n222 & n223 ;
  assign n225 = x7 & n198 ;
  assign n226 = ~n224 & ~n225 ;
  assign n227 = ~n221 & ~n226 ;
  assign n228 = x0 & n13 ;
  assign n229 = ~x6 & n44 ;
  assign n230 = ~n228 & ~n229 ;
  assign n231 = ~n87 & ~n90 ;
  assign n232 = ~x7 & n231 ;
  assign n233 = ~n230 & n232 ;
  assign n234 = ~x0 & x7 ;
  assign n235 = n90 & n234 ;
  assign n236 = n53 & n235 ;
  assign n237 = ~n233 & ~n236 ;
  assign n238 = ~x1 & ~x5 ;
  assign n239 = ~n237 & n238 ;
  assign n240 = x1 & n112 ;
  assign n241 = n68 ^ x0 ;
  assign n242 = n241 ^ n68 ;
  assign n243 = ~n143 & ~n223 ;
  assign n244 = n231 & ~n243 ;
  assign n245 = n244 ^ n68 ;
  assign n246 = ~n242 & n245 ;
  assign n247 = n246 ^ n68 ;
  assign n248 = n240 & n247 ;
  assign n249 = ~n239 & ~n248 ;
  assign n250 = ~n227 & n249 ;
  assign n251 = n250 ^ x4 ;
  assign n252 = n251 ^ n250 ;
  assign n253 = n252 ^ x2 ;
  assign n254 = x0 & n190 ;
  assign n255 = ~x0 & ~x6 ;
  assign n256 = ~x7 & n255 ;
  assign n257 = n143 & n256 ;
  assign n258 = ~n254 & ~n257 ;
  assign n259 = n103 & ~n258 ;
  assign n260 = ~x7 & n198 ;
  assign n261 = ~n224 & ~n260 ;
  assign n262 = n162 & ~n261 ;
  assign n264 = n222 & ~n255 ;
  assign n265 = ~n19 & ~n35 ;
  assign n266 = n264 & n265 ;
  assign n267 = ~x9 & ~n87 ;
  assign n268 = n234 & n267 ;
  assign n269 = ~n266 & ~n268 ;
  assign n263 = n15 & n90 ;
  assign n270 = n269 ^ n263 ;
  assign n271 = x5 & ~n270 ;
  assign n272 = n271 ^ n269 ;
  assign n273 = ~n262 & n272 ;
  assign n274 = ~x8 & ~n273 ;
  assign n275 = x9 ^ x7 ;
  assign n276 = n167 & ~n275 ;
  assign n277 = n127 ^ n112 ;
  assign n278 = n277 ^ n127 ;
  assign n279 = n127 ^ x6 ;
  assign n280 = n279 ^ n127 ;
  assign n281 = ~n278 & n280 ;
  assign n282 = n281 ^ n127 ;
  assign n283 = x3 & n282 ;
  assign n284 = n283 ^ n127 ;
  assign n285 = n276 & n284 ;
  assign n286 = ~x0 & x9 ;
  assign n287 = n36 & n103 ;
  assign n288 = ~n73 & n287 ;
  assign n289 = ~n286 & n288 ;
  assign n290 = n44 & n184 ;
  assign n291 = ~x1 & ~n290 ;
  assign n292 = ~n289 & n291 ;
  assign n293 = ~n285 & n292 ;
  assign n294 = ~n274 & n293 ;
  assign n295 = x8 & n286 ;
  assign n296 = x7 & ~n87 ;
  assign n297 = ~n141 & ~n222 ;
  assign n298 = ~n296 & n297 ;
  assign n299 = n295 & n298 ;
  assign n300 = x1 & ~n299 ;
  assign n301 = n267 ^ n219 ;
  assign n302 = n256 ^ x3 ;
  assign n303 = n302 ^ n256 ;
  assign n304 = n256 ^ x7 ;
  assign n305 = ~n303 & n304 ;
  assign n306 = n305 ^ n256 ;
  assign n307 = n306 ^ n219 ;
  assign n308 = n301 & n307 ;
  assign n309 = n308 ^ n305 ;
  assign n310 = n309 ^ n256 ;
  assign n311 = n310 ^ n267 ;
  assign n312 = n219 & n311 ;
  assign n313 = n312 ^ n219 ;
  assign n314 = n300 & ~n313 ;
  assign n315 = ~x0 & n132 ;
  assign n316 = ~n275 & n315 ;
  assign n317 = n17 ^ x6 ;
  assign n318 = n317 ^ n17 ;
  assign n319 = n17 ^ n13 ;
  assign n320 = n319 ^ n17 ;
  assign n321 = ~n318 & n320 ;
  assign n322 = n321 ^ n17 ;
  assign n323 = ~x0 & n322 ;
  assign n324 = n323 ^ n17 ;
  assign n325 = ~n316 & ~n324 ;
  assign n326 = x3 & ~n325 ;
  assign n327 = ~n141 & n286 ;
  assign n328 = n327 ^ n87 ;
  assign n329 = n328 ^ n326 ;
  assign n330 = n74 ^ n25 ;
  assign n331 = ~n87 & ~n330 ;
  assign n332 = n331 ^ n25 ;
  assign n333 = ~n329 & ~n332 ;
  assign n334 = n333 ^ n331 ;
  assign n335 = n334 ^ n25 ;
  assign n336 = n335 ^ n87 ;
  assign n337 = ~n326 & n336 ;
  assign n338 = n337 ^ x5 ;
  assign n339 = n338 ^ n337 ;
  assign n340 = n339 ^ n314 ;
  assign n341 = n13 & n222 ;
  assign n342 = ~n45 & ~n341 ;
  assign n343 = n342 ^ x0 ;
  assign n344 = ~n342 & ~n343 ;
  assign n345 = n344 ^ n337 ;
  assign n346 = n345 ^ n342 ;
  assign n347 = n340 & n346 ;
  assign n348 = n347 ^ n344 ;
  assign n349 = n348 ^ n342 ;
  assign n350 = n314 & ~n349 ;
  assign n351 = n350 ^ n314 ;
  assign n352 = ~n294 & ~n351 ;
  assign n353 = n352 ^ n259 ;
  assign n354 = ~n259 & n353 ;
  assign n355 = n354 ^ n250 ;
  assign n356 = n355 ^ n259 ;
  assign n357 = n253 & ~n356 ;
  assign n358 = n357 ^ n354 ;
  assign n359 = n358 ^ n259 ;
  assign n360 = x2 & ~n359 ;
  assign n361 = n360 ^ x2 ;
  assign n362 = n216 & ~n361 ;
  assign n363 = ~n189 & n362 ;
  assign y0 = ~n363 ;
endmodule
