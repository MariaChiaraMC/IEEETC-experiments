module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 ;
  assign n16 = x12 ^ x11 ;
  assign n17 = ~x0 & ~x10 ;
  assign n19 = x10 & x14 ;
  assign n18 = x0 & ~x1 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = x9 & ~x13 ;
  assign n23 = n22 ^ n18 ;
  assign n24 = ~n21 & ~n23 ;
  assign n25 = n24 ^ n18 ;
  assign n26 = ~n17 & ~n25 ;
  assign n27 = x9 & ~x10 ;
  assign n28 = n27 ^ x13 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = x2 & ~x9 ;
  assign n32 = n17 & ~n31 ;
  assign n33 = x1 & ~n32 ;
  assign n34 = ~x9 & ~x10 ;
  assign n35 = ~x0 & x2 ;
  assign n36 = x4 & x6 ;
  assign n37 = n35 & n36 ;
  assign n38 = ~x5 & n37 ;
  assign n42 = x5 ^ x4 ;
  assign n39 = x4 ^ x2 ;
  assign n43 = n42 ^ n39 ;
  assign n40 = n39 ^ x4 ;
  assign n41 = n40 ^ x4 ;
  assign n44 = n43 ^ n41 ;
  assign n47 = x7 ^ x4 ;
  assign n48 = n47 ^ x4 ;
  assign n45 = x6 ^ x4 ;
  assign n46 = n45 ^ x0 ;
  assign n49 = n48 ^ n46 ;
  assign n50 = ~n40 & n49 ;
  assign n51 = n50 ^ n45 ;
  assign n52 = n51 ^ n46 ;
  assign n53 = n52 ^ n40 ;
  assign n54 = n53 ^ n48 ;
  assign n55 = ~n44 & n54 ;
  assign n56 = n55 ^ n40 ;
  assign n57 = n56 ^ n41 ;
  assign n58 = n53 ^ n41 ;
  assign n59 = n41 & ~n58 ;
  assign n60 = n59 ^ n40 ;
  assign n61 = ~n57 & ~n60 ;
  assign n62 = n61 ^ n45 ;
  assign n63 = n62 ^ n40 ;
  assign n64 = n63 ^ n41 ;
  assign n65 = n64 ^ x4 ;
  assign n66 = n65 ^ n45 ;
  assign n67 = ~n38 & ~n66 ;
  assign n68 = n67 ^ x3 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = ~x4 & n35 ;
  assign n71 = x5 ^ x2 ;
  assign n72 = ~x4 & n71 ;
  assign n73 = n72 ^ x2 ;
  assign n74 = ~n70 & ~n73 ;
  assign n75 = x0 & x2 ;
  assign n76 = x6 & n75 ;
  assign n77 = x5 & n76 ;
  assign n78 = ~n74 & ~n77 ;
  assign n79 = n78 ^ n67 ;
  assign n80 = n69 & n79 ;
  assign n81 = n80 ^ n67 ;
  assign n82 = n34 & n81 ;
  assign n83 = n33 & ~n82 ;
  assign n84 = x6 & x7 ;
  assign n85 = x5 & ~n84 ;
  assign n86 = ~x2 & ~x3 ;
  assign n87 = ~x4 & n86 ;
  assign n88 = ~n85 & n87 ;
  assign n89 = x9 & n17 ;
  assign n90 = ~n88 & n89 ;
  assign n91 = x0 & n86 ;
  assign n92 = n19 & n91 ;
  assign n93 = ~x1 & ~n92 ;
  assign n94 = n36 & n86 ;
  assign n95 = x7 & n94 ;
  assign n96 = n95 ^ n34 ;
  assign n97 = n86 ^ x0 ;
  assign n98 = n97 ^ n86 ;
  assign n99 = x2 & x6 ;
  assign n100 = ~x7 & n99 ;
  assign n101 = x5 & ~n100 ;
  assign n102 = n101 ^ n86 ;
  assign n103 = ~n98 & ~n102 ;
  assign n104 = n103 ^ n86 ;
  assign n105 = n104 ^ n95 ;
  assign n106 = ~n96 & n105 ;
  assign n107 = n106 ^ n103 ;
  assign n108 = n107 ^ n86 ;
  assign n109 = n108 ^ n34 ;
  assign n110 = ~n95 & ~n109 ;
  assign n111 = n110 ^ n95 ;
  assign n112 = n93 & n111 ;
  assign n113 = ~n90 & n112 ;
  assign n114 = n113 ^ n83 ;
  assign n115 = ~n83 & n114 ;
  assign n116 = n115 ^ n27 ;
  assign n117 = n116 ^ n83 ;
  assign n118 = n30 & n117 ;
  assign n119 = n118 ^ n115 ;
  assign n120 = n119 ^ n83 ;
  assign n121 = ~n26 & ~n120 ;
  assign n122 = n121 ^ n26 ;
  assign n123 = n122 ^ x12 ;
  assign n124 = n123 ^ n122 ;
  assign n125 = n124 ^ n16 ;
  assign n126 = n22 ^ x10 ;
  assign n127 = n22 & n126 ;
  assign n128 = n127 ^ n122 ;
  assign n129 = n128 ^ n22 ;
  assign n130 = ~n125 & n129 ;
  assign n131 = n130 ^ n127 ;
  assign n132 = n131 ^ n22 ;
  assign n133 = ~n16 & n132 ;
  assign y0 = n133 ;
endmodule
