module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 ;
  assign n16 = ~x5 & ~x7 ;
  assign n17 = ~x9 & ~x13 ;
  assign n18 = ~x14 & n17 ;
  assign n19 = n16 & n18 ;
  assign n20 = x1 & ~n19 ;
  assign n21 = ~x8 & ~x10 ;
  assign n22 = ~x2 & n21 ;
  assign n23 = ~x6 & ~x11 ;
  assign n24 = ~x4 & ~x12 ;
  assign n25 = n23 & n24 ;
  assign n26 = ~x0 & ~x3 ;
  assign n27 = n25 & n26 ;
  assign n28 = n22 & n27 ;
  assign n29 = ~n20 & n28 ;
  assign n30 = n18 ^ x7 ;
  assign n31 = n30 ^ x5 ;
  assign n32 = n31 ^ n18 ;
  assign n33 = n32 ^ x1 ;
  assign n34 = x13 ^ x9 ;
  assign n35 = x14 & n34 ;
  assign n36 = n35 ^ x5 ;
  assign n37 = ~x5 & ~n36 ;
  assign n38 = n37 ^ n18 ;
  assign n39 = n38 ^ x5 ;
  assign n40 = n33 & ~n39 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n41 ^ x5 ;
  assign n43 = ~x1 & ~n42 ;
  assign n44 = n43 ^ x1 ;
  assign n45 = n29 & n44 ;
  assign y0 = n45 ;
endmodule
