module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 ;
  assign n20 = ~x6 & ~x16 ;
  assign n21 = x8 ^ x7 ;
  assign n22 = ~x10 & x15 ;
  assign n23 = ~x2 & n22 ;
  assign n24 = ~x14 & n23 ;
  assign n25 = n24 ^ x8 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = x14 & ~x15 ;
  assign n28 = n27 ^ x9 ;
  assign n29 = x8 & n28 ;
  assign n30 = n29 ^ x9 ;
  assign n31 = n26 & ~n30 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = n32 ^ x9 ;
  assign n34 = n33 ^ x8 ;
  assign n35 = n21 & ~n34 ;
  assign n36 = n20 & n35 ;
  assign n41 = x8 & x9 ;
  assign n42 = x4 & x7 ;
  assign n43 = ~n41 & n42 ;
  assign n37 = ~x3 & ~x15 ;
  assign n38 = n37 ^ x15 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = n44 ^ n38 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = n39 ^ n38 ;
  assign n46 = n45 ^ n40 ;
  assign n47 = n38 ^ x6 ;
  assign n48 = n47 ^ x16 ;
  assign n49 = n48 ^ n38 ;
  assign n50 = n49 ^ n45 ;
  assign n51 = n45 & ~n50 ;
  assign n52 = n51 ^ n45 ;
  assign n53 = n46 & n52 ;
  assign n54 = n53 ^ n51 ;
  assign n55 = n54 ^ n38 ;
  assign n56 = n55 ^ n45 ;
  assign n57 = ~x14 & n56 ;
  assign n58 = n57 ^ x15 ;
  assign n59 = x18 & ~n58 ;
  assign n60 = ~n36 & ~n59 ;
  assign n61 = n60 ^ x18 ;
  assign n62 = n61 ^ x17 ;
  assign n71 = n62 ^ n61 ;
  assign n63 = x6 & x16 ;
  assign n64 = n35 & n63 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = n65 ^ n61 ;
  assign n67 = n62 ^ n60 ;
  assign n68 = n67 ^ n64 ;
  assign n69 = n68 ^ n66 ;
  assign n70 = ~n66 & n69 ;
  assign n72 = n71 ^ n70 ;
  assign n73 = n72 ^ n66 ;
  assign n74 = x16 ^ x1 ;
  assign n75 = x13 ^ x11 ;
  assign n76 = n75 ^ x11 ;
  assign n77 = ~x11 & x12 ;
  assign n78 = n77 ^ x11 ;
  assign n79 = n76 & n78 ;
  assign n80 = n79 ^ x11 ;
  assign n81 = n80 ^ x16 ;
  assign n82 = ~n74 & ~n81 ;
  assign n83 = n82 ^ n79 ;
  assign n84 = n83 ^ x11 ;
  assign n85 = n84 ^ x1 ;
  assign n86 = ~x16 & n85 ;
  assign n87 = n86 ^ x16 ;
  assign n88 = ~x15 & ~n87 ;
  assign n90 = x7 & x8 ;
  assign n89 = ~x8 & ~x9 ;
  assign n91 = n90 ^ n89 ;
  assign n92 = n91 ^ n90 ;
  assign n93 = n90 ^ x7 ;
  assign n94 = n93 ^ n90 ;
  assign n95 = n92 & ~n94 ;
  assign n96 = n95 ^ n90 ;
  assign n97 = x6 & n96 ;
  assign n98 = n97 ^ n90 ;
  assign n99 = n98 ^ n37 ;
  assign n100 = n99 ^ n37 ;
  assign n101 = n37 ^ n23 ;
  assign n102 = n100 & n101 ;
  assign n103 = n102 ^ n37 ;
  assign n104 = ~x4 & n37 ;
  assign n105 = n104 ^ x16 ;
  assign n106 = n103 & n105 ;
  assign n107 = n106 ^ n104 ;
  assign n108 = x16 & n107 ;
  assign n109 = n108 ^ x16 ;
  assign n110 = ~n88 & ~n109 ;
  assign n111 = ~x14 & ~n110 ;
  assign n112 = ~x6 & n90 ;
  assign n113 = n27 & ~n112 ;
  assign n114 = x16 & n113 ;
  assign n115 = ~n111 & ~n114 ;
  assign n116 = n115 ^ n61 ;
  assign n117 = n70 ^ n66 ;
  assign n118 = n116 & ~n117 ;
  assign n119 = n118 ^ n61 ;
  assign n120 = ~n73 & n119 ;
  assign n121 = n120 ^ n61 ;
  assign n122 = n121 ^ x18 ;
  assign n123 = n122 ^ n61 ;
  assign y0 = ~n123 ;
endmodule
