module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n7 = x2 ^ x1 ;
  assign n8 = x3 ^ x1 ;
  assign n9 = n8 ^ x1 ;
  assign n10 = n9 ^ n7 ;
  assign n11 = n7 & n10 ;
  assign n12 = n11 ^ x1 ;
  assign n13 = n12 ^ n7 ;
  assign n15 = x5 ^ x1 ;
  assign n14 = x2 ^ x0 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = x5 & ~n16 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = n18 ^ x1 ;
  assign n20 = x5 ^ x4 ;
  assign n21 = ~n15 & ~n20 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = n22 ^ n14 ;
  assign n24 = ~n19 & ~n23 ;
  assign n25 = n24 ^ n14 ;
  assign n26 = ~n13 & n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n27 ^ n14 ;
  assign y0 = n28 ;
endmodule
