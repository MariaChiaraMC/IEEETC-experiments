module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 ;
  assign n8 = x3 ^ x2 ;
  assign n9 = n8 ^ x3 ;
  assign n10 = n9 ^ n8 ;
  assign n12 = x3 ^ x0 ;
  assign n11 = x2 ^ x1 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n13 ^ n9 ;
  assign n15 = n14 ^ n9 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = n16 ^ n12 ;
  assign n18 = n17 ^ n10 ;
  assign n19 = ~n10 & n18 ;
  assign n20 = n19 ^ n9 ;
  assign n21 = n17 ^ n8 ;
  assign n26 = x4 & x5 ;
  assign n27 = x6 & n26 ;
  assign n28 = n27 ^ n16 ;
  assign n29 = n16 ^ n8 ;
  assign n30 = n29 ^ n9 ;
  assign n31 = n30 ^ n17 ;
  assign n32 = ~n28 & n31 ;
  assign n22 = ~x4 & ~x5 ;
  assign n23 = n22 ^ n12 ;
  assign n24 = n23 ^ n16 ;
  assign n25 = ~n17 & ~n24 ;
  assign n33 = n32 ^ n25 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = n34 ^ n16 ;
  assign n36 = n35 ^ n9 ;
  assign n37 = n21 & ~n36 ;
  assign n38 = n37 ^ n25 ;
  assign n39 = n38 ^ n16 ;
  assign n40 = n39 ^ n17 ;
  assign n41 = n20 & ~n40 ;
  assign n42 = n41 ^ n25 ;
  assign n43 = n42 ^ n37 ;
  assign n44 = n43 ^ n16 ;
  assign n45 = n44 ^ n17 ;
  assign n46 = n45 ^ n11 ;
  assign y0 = n46 ;
endmodule
