module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 ;
  assign n16 = ~x9 & ~x14 ;
  assign n17 = ~x8 & ~n16 ;
  assign n18 = ~x5 & x6 ;
  assign n19 = x3 ^ x2 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = x4 ^ x3 ;
  assign n22 = ~n20 & n21 ;
  assign n23 = n22 ^ x3 ;
  assign n24 = x1 & ~n23 ;
  assign n25 = n18 & ~n24 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = n25 ^ x3 ;
  assign n28 = n27 ^ x3 ;
  assign n29 = x5 & ~x6 ;
  assign n30 = n29 ^ x3 ;
  assign n31 = ~n28 & n30 ;
  assign n32 = n31 ^ x3 ;
  assign n33 = ~n26 & ~n32 ;
  assign n34 = n33 ^ x4 ;
  assign n35 = ~n17 & ~n34 ;
  assign n36 = ~x1 & ~x8 ;
  assign n37 = ~x3 & ~n36 ;
  assign n38 = n29 & ~n37 ;
  assign n39 = x8 ^ x4 ;
  assign n40 = n39 ^ n16 ;
  assign n41 = n16 ^ x3 ;
  assign n42 = x8 ^ x3 ;
  assign n43 = n41 & n42 ;
  assign n44 = n43 ^ x3 ;
  assign n45 = ~n40 & n44 ;
  assign n46 = n45 ^ x4 ;
  assign n47 = n38 & n46 ;
  assign n48 = ~x2 & n47 ;
  assign n49 = ~n35 & ~n48 ;
  assign n50 = x7 & x13 ;
  assign n51 = ~n49 & n50 ;
  assign y0 = n51 ;
endmodule
