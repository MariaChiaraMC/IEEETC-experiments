module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 ;
  assign n9 = ~x1 & ~x2 ;
  assign n10 = x3 & n9 ;
  assign n11 = ~x0 & n10 ;
  assign n12 = x6 ^ x5 ;
  assign n13 = x7 ^ x6 ;
  assign n14 = x7 ^ x4 ;
  assign n15 = ~x7 & n14 ;
  assign n16 = n15 ^ x7 ;
  assign n17 = ~n13 & ~n16 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n18 ^ x7 ;
  assign n20 = n19 ^ x4 ;
  assign n21 = ~n12 & n20 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = n11 & n22 ;
  assign y0 = ~n23 ;
endmodule
