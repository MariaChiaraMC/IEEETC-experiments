module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 ;
  assign n7 = x3 & ~x5 ;
  assign n8 = n7 ^ x1 ;
  assign n9 = n8 ^ n7 ;
  assign n10 = ~x3 & x5 ;
  assign n11 = n10 ^ n7 ;
  assign n12 = ~n9 & n11 ;
  assign n13 = n12 ^ n7 ;
  assign n14 = ~x0 & n13 ;
  assign n15 = x2 & n14 ;
  assign n16 = x2 & ~x4 ;
  assign n17 = n16 ^ n10 ;
  assign n18 = ~x1 & ~x5 ;
  assign n19 = n18 ^ n10 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = x0 & x1 ;
  assign n22 = ~x4 & ~n21 ;
  assign n23 = n22 ^ n18 ;
  assign n24 = n20 & n23 ;
  assign n25 = n24 ^ n18 ;
  assign n26 = n17 & ~n25 ;
  assign n27 = ~n15 & ~n26 ;
  assign n28 = n7 ^ x2 ;
  assign n29 = n28 ^ x4 ;
  assign n34 = n29 ^ x2 ;
  assign n35 = n34 ^ x4 ;
  assign n36 = n35 ^ x4 ;
  assign n37 = x2 ^ x0 ;
  assign n38 = n37 ^ x4 ;
  assign n39 = ~n36 & n38 ;
  assign n30 = x2 ^ x1 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n31 ^ x4 ;
  assign n33 = n29 & ~n32 ;
  assign n40 = n39 ^ n33 ;
  assign n41 = n40 ^ n29 ;
  assign n42 = n33 ^ x4 ;
  assign n43 = n42 ^ n35 ;
  assign n44 = ~x4 & ~n43 ;
  assign n45 = n44 ^ n33 ;
  assign n46 = n41 & n45 ;
  assign n47 = n46 ^ n39 ;
  assign n48 = n47 ^ n44 ;
  assign n49 = n48 ^ n29 ;
  assign n50 = n49 ^ x4 ;
  assign n51 = n50 ^ n35 ;
  assign n52 = n27 & n51 ;
  assign y0 = n52 ;
endmodule
