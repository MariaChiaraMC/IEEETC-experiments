module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 ;
  assign n10 = x2 & ~x4 ;
  assign n11 = x5 & ~x6 ;
  assign n12 = n11 ^ x5 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = x6 & ~x7 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = n15 ^ n11 ;
  assign n17 = ~n13 & n16 ;
  assign n18 = n17 ^ n11 ;
  assign n19 = x3 & n18 ;
  assign n20 = n19 ^ n11 ;
  assign n21 = n10 & n20 ;
  assign n22 = ~x8 & n21 ;
  assign n23 = ~x2 & ~x3 ;
  assign n24 = n14 & n23 ;
  assign n25 = ~x8 & n24 ;
  assign n26 = ~x2 & x7 ;
  assign n27 = ~x3 & x6 ;
  assign n28 = ~x8 & n27 ;
  assign n29 = ~n26 & ~n28 ;
  assign n30 = x7 & ~x8 ;
  assign n31 = x1 & ~n30 ;
  assign n32 = ~n29 & n31 ;
  assign n33 = ~n25 & ~n32 ;
  assign n34 = ~x5 & ~n33 ;
  assign n35 = x5 & n23 ;
  assign n36 = x3 & ~x5 ;
  assign n37 = x1 & n36 ;
  assign n38 = ~n35 & ~n37 ;
  assign n39 = x6 & x8 ;
  assign n40 = ~x6 & ~x8 ;
  assign n41 = x7 & n40 ;
  assign n42 = ~n39 & ~n41 ;
  assign n43 = ~n38 & ~n42 ;
  assign n44 = ~x5 & ~x6 ;
  assign n45 = x1 & x8 ;
  assign n46 = n44 & n45 ;
  assign n47 = n46 ^ x2 ;
  assign n48 = n47 ^ x3 ;
  assign n49 = n48 ^ n46 ;
  assign n50 = n49 ^ n48 ;
  assign n51 = x6 & x7 ;
  assign n52 = x3 & x8 ;
  assign n53 = n51 & n52 ;
  assign n54 = ~x3 & x7 ;
  assign n55 = n44 & n54 ;
  assign n56 = ~n53 & ~n55 ;
  assign n57 = n56 ^ n48 ;
  assign n58 = n57 ^ n47 ;
  assign n59 = n50 & ~n58 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = x7 & n56 ;
  assign n62 = n61 ^ n47 ;
  assign n63 = n60 & ~n62 ;
  assign n64 = n63 ^ n61 ;
  assign n65 = ~n47 & n64 ;
  assign n66 = n65 ^ n59 ;
  assign n67 = n66 ^ x2 ;
  assign n68 = n67 ^ n56 ;
  assign n69 = ~n43 & ~n68 ;
  assign n70 = ~n34 & n69 ;
  assign n71 = x4 & ~n70 ;
  assign n72 = x4 & n30 ;
  assign n73 = n11 & n72 ;
  assign n74 = n27 & n30 ;
  assign n75 = ~x5 & n74 ;
  assign n76 = ~x5 & x6 ;
  assign n77 = ~x3 & ~n76 ;
  assign n78 = x7 ^ x5 ;
  assign n79 = ~n77 & n78 ;
  assign n80 = n79 ^ x4 ;
  assign n81 = n80 ^ n79 ;
  assign n82 = ~x6 & ~x7 ;
  assign n83 = ~x3 & n82 ;
  assign n84 = n83 ^ n79 ;
  assign n85 = ~n81 & n84 ;
  assign n86 = n85 ^ n79 ;
  assign n87 = x8 & n86 ;
  assign n88 = ~n75 & ~n87 ;
  assign n89 = ~n73 & n88 ;
  assign n107 = x5 & x6 ;
  assign n117 = ~x8 & n107 ;
  assign n118 = n30 ^ x4 ;
  assign n119 = n118 ^ n30 ;
  assign n120 = ~x8 & n82 ;
  assign n121 = x5 & x7 ;
  assign n122 = ~n30 & n121 ;
  assign n123 = ~n120 & ~n122 ;
  assign n124 = n123 ^ n30 ;
  assign n125 = ~n119 & ~n124 ;
  assign n126 = n125 ^ n30 ;
  assign n127 = ~n117 & ~n126 ;
  assign n128 = x3 & ~n127 ;
  assign n90 = ~x4 & ~x5 ;
  assign n91 = ~x3 & ~n82 ;
  assign n92 = n90 & ~n91 ;
  assign n93 = ~n51 & n92 ;
  assign n94 = ~x3 & x4 ;
  assign n95 = n94 ^ x7 ;
  assign n96 = n95 ^ n94 ;
  assign n97 = ~x4 & x5 ;
  assign n98 = n97 ^ n94 ;
  assign n99 = n98 ^ n94 ;
  assign n100 = ~n96 & n99 ;
  assign n101 = n100 ^ n94 ;
  assign n102 = x6 & n101 ;
  assign n103 = n102 ^ n94 ;
  assign n104 = n103 ^ x8 ;
  assign n105 = n104 ^ n103 ;
  assign n106 = n105 ^ n93 ;
  assign n108 = n107 ^ x7 ;
  assign n109 = n107 & n108 ;
  assign n110 = n109 ^ n103 ;
  assign n111 = n110 ^ n107 ;
  assign n112 = n106 & n111 ;
  assign n113 = n112 ^ n109 ;
  assign n114 = n113 ^ n107 ;
  assign n115 = ~n93 & n114 ;
  assign n116 = n115 ^ n93 ;
  assign n129 = n128 ^ n116 ;
  assign n130 = n129 ^ n116 ;
  assign n131 = n14 & n90 ;
  assign n132 = x8 & n131 ;
  assign n133 = n132 ^ n116 ;
  assign n134 = n133 ^ n116 ;
  assign n135 = ~n130 & ~n134 ;
  assign n136 = n135 ^ n116 ;
  assign n137 = ~x2 & ~n136 ;
  assign n138 = n137 ^ n116 ;
  assign n139 = n89 & ~n138 ;
  assign n140 = n139 ^ x1 ;
  assign n141 = n140 ^ n139 ;
  assign n142 = n141 ^ n71 ;
  assign n143 = x6 & ~n10 ;
  assign n144 = n91 & ~n143 ;
  assign n145 = n144 ^ x2 ;
  assign n146 = n145 ^ n144 ;
  assign n147 = ~x4 & n54 ;
  assign n148 = ~n82 & ~n147 ;
  assign n149 = n148 ^ n144 ;
  assign n150 = n149 ^ n144 ;
  assign n151 = ~n146 & ~n150 ;
  assign n152 = n151 ^ n144 ;
  assign n153 = ~x8 & n152 ;
  assign n154 = n153 ^ n144 ;
  assign n155 = ~n53 & ~n154 ;
  assign n156 = ~x5 & n155 ;
  assign n157 = x3 & ~x8 ;
  assign n158 = ~x6 & x7 ;
  assign n159 = ~n157 & ~n158 ;
  assign n160 = x2 & ~n30 ;
  assign n161 = ~n52 & ~n160 ;
  assign n162 = ~n159 & ~n161 ;
  assign n163 = n162 ^ x5 ;
  assign n165 = x8 ^ x3 ;
  assign n164 = x8 ^ x7 ;
  assign n171 = n165 ^ n164 ;
  assign n168 = n165 ^ x6 ;
  assign n172 = n171 ^ n168 ;
  assign n173 = n172 ^ n168 ;
  assign n174 = n165 ^ x8 ;
  assign n175 = n174 ^ n165 ;
  assign n176 = n175 ^ n168 ;
  assign n177 = n173 & n176 ;
  assign n166 = n165 ^ x2 ;
  assign n167 = n166 ^ n164 ;
  assign n169 = n168 ^ n167 ;
  assign n170 = n164 & ~n169 ;
  assign n178 = n177 ^ n170 ;
  assign n179 = n178 ^ n164 ;
  assign n180 = n170 ^ n168 ;
  assign n181 = n180 ^ n172 ;
  assign n182 = n168 & n181 ;
  assign n183 = n182 ^ n170 ;
  assign n184 = n179 & n183 ;
  assign n185 = n184 ^ n177 ;
  assign n186 = n185 ^ n182 ;
  assign n187 = n186 ^ n164 ;
  assign n188 = n187 ^ n168 ;
  assign n189 = n188 ^ n172 ;
  assign n190 = n189 ^ x4 ;
  assign n191 = n190 ^ n189 ;
  assign n192 = x6 ^ x3 ;
  assign n193 = n39 & n192 ;
  assign n194 = n193 ^ n192 ;
  assign n195 = x2 & n194 ;
  assign n196 = ~n120 & ~n195 ;
  assign n197 = n196 ^ n189 ;
  assign n198 = n191 & ~n197 ;
  assign n199 = n198 ^ n189 ;
  assign n200 = n199 ^ n162 ;
  assign n201 = ~n163 & n200 ;
  assign n202 = n201 ^ n198 ;
  assign n203 = n202 ^ n189 ;
  assign n204 = n203 ^ x5 ;
  assign n205 = ~n162 & ~n204 ;
  assign n206 = n205 ^ n162 ;
  assign n207 = n206 ^ n156 ;
  assign n208 = ~n156 & ~n207 ;
  assign n209 = n208 ^ n139 ;
  assign n210 = n209 ^ n156 ;
  assign n211 = ~n142 & n210 ;
  assign n212 = n211 ^ n208 ;
  assign n213 = n212 ^ n156 ;
  assign n214 = ~n71 & ~n213 ;
  assign n215 = n214 ^ n71 ;
  assign n216 = ~n22 & ~n215 ;
  assign n217 = ~x0 & ~n216 ;
  assign n218 = x6 ^ x5 ;
  assign n219 = n218 ^ x8 ;
  assign n220 = x8 ^ x0 ;
  assign n221 = n220 ^ x0 ;
  assign n222 = n221 ^ n219 ;
  assign n223 = x6 ^ x4 ;
  assign n224 = ~x6 & n223 ;
  assign n225 = n224 ^ x0 ;
  assign n226 = n225 ^ x6 ;
  assign n227 = ~n222 & ~n226 ;
  assign n228 = n227 ^ n224 ;
  assign n229 = n228 ^ x6 ;
  assign n230 = n219 & ~n229 ;
  assign n231 = n230 ^ x7 ;
  assign n232 = n231 ^ n230 ;
  assign n233 = n232 ^ n23 ;
  assign n234 = ~x0 & n39 ;
  assign n235 = ~n40 & ~n107 ;
  assign n236 = n235 ^ x4 ;
  assign n237 = n235 ^ x0 ;
  assign n238 = n237 ^ x0 ;
  assign n239 = n44 ^ x0 ;
  assign n240 = n238 & ~n239 ;
  assign n241 = n240 ^ x0 ;
  assign n242 = ~n236 & n241 ;
  assign n243 = n242 ^ n234 ;
  assign n244 = ~n234 & n243 ;
  assign n245 = n244 ^ n230 ;
  assign n246 = n245 ^ n234 ;
  assign n247 = n233 & n246 ;
  assign n248 = n247 ^ n244 ;
  assign n249 = n248 ^ n234 ;
  assign n250 = n23 & ~n249 ;
  assign n251 = n250 ^ n23 ;
  assign n252 = ~x1 & n251 ;
  assign n253 = ~n217 & ~n252 ;
  assign y0 = ~n253 ;
endmodule
