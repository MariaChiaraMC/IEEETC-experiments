module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 ;
  output y0 ;
  wire n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 ;
  assign n14 = ~x3 & x4 ;
  assign n15 = ~x2 & ~n14 ;
  assign n16 = x11 & ~n15 ;
  assign n17 = ~x7 & ~n16 ;
  assign n18 = ~x8 & ~n17 ;
  assign n19 = x10 ^ x9 ;
  assign n66 = n19 ^ x10 ;
  assign n39 = ~x2 & ~x3 ;
  assign n49 = x0 & ~x1 ;
  assign n50 = ~n39 & n49 ;
  assign n51 = x12 & ~n50 ;
  assign n20 = x5 & ~x6 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = ~x1 & ~n21 ;
  assign n23 = n22 ^ x2 ;
  assign n40 = n39 ^ n23 ;
  assign n24 = x6 ^ x4 ;
  assign n25 = x5 & ~n24 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = x3 ^ x1 ;
  assign n28 = x6 ^ x3 ;
  assign n29 = x6 ^ x2 ;
  assign n30 = x6 & n29 ;
  assign n31 = n30 ^ x6 ;
  assign n32 = ~n28 & n31 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ x6 ;
  assign n35 = n34 ^ x2 ;
  assign n36 = ~n27 & n35 ;
  assign n37 = n26 & n36 ;
  assign n38 = n37 ^ n23 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = ~x1 & x5 ;
  assign n43 = n42 ^ n40 ;
  assign n44 = n43 ^ n40 ;
  assign n45 = n41 & ~n44 ;
  assign n46 = n45 ^ n40 ;
  assign n47 = x0 & ~n46 ;
  assign n48 = n47 ^ n23 ;
  assign n52 = n51 ^ n48 ;
  assign n53 = n52 ^ n48 ;
  assign n54 = n48 ^ x10 ;
  assign n55 = n54 ^ n48 ;
  assign n56 = ~n53 & ~n55 ;
  assign n57 = n56 ^ n48 ;
  assign n58 = x8 & n57 ;
  assign n59 = n58 ^ n48 ;
  assign n60 = n59 ^ n19 ;
  assign n61 = n60 ^ x10 ;
  assign n62 = n59 ^ x11 ;
  assign n63 = n62 ^ n59 ;
  assign n64 = n63 ^ n61 ;
  assign n65 = n61 & ~n64 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = n67 ^ n61 ;
  assign n69 = x7 & x10 ;
  assign n70 = n69 ^ x10 ;
  assign n71 = n65 ^ n61 ;
  assign n72 = ~n70 & n71 ;
  assign n73 = n72 ^ x10 ;
  assign n74 = ~n68 & ~n73 ;
  assign n75 = n74 ^ x10 ;
  assign n76 = n75 ^ x10 ;
  assign n77 = ~n18 & n76 ;
  assign y0 = n77 ;
endmodule
