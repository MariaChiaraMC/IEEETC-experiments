module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 ;
  assign n9 = ~x2 & x7 ;
  assign n10 = x0 & n9 ;
  assign n11 = x2 & ~x7 ;
  assign n12 = x0 & x1 ;
  assign n13 = ~n11 & ~n12 ;
  assign n14 = x5 & n13 ;
  assign n15 = ~n10 & n14 ;
  assign n16 = x1 ^ x0 ;
  assign n17 = n16 ^ n11 ;
  assign n18 = n17 ^ x3 ;
  assign n19 = n9 ^ x5 ;
  assign n20 = ~n11 & n19 ;
  assign n21 = n20 ^ x5 ;
  assign n22 = n18 & n21 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n24 ^ n11 ;
  assign n26 = ~x3 & ~n25 ;
  assign n27 = ~n15 & n26 ;
  assign y0 = ~n27 ;
endmodule
