module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 ;
  assign n17 = ~x5 & x6 ;
  assign n18 = x11 ^ x10 ;
  assign n19 = ~x5 & n18 ;
  assign n20 = ~x4 & ~n19 ;
  assign n21 = ~n17 & ~n20 ;
  assign n22 = ~x10 & ~x11 ;
  assign n23 = x6 ^ x5 ;
  assign n24 = x9 ^ x6 ;
  assign n25 = n23 & ~n24 ;
  assign n26 = n25 ^ x6 ;
  assign n27 = n22 & n26 ;
  assign n28 = ~n21 & ~n27 ;
  assign n29 = x7 & ~n28 ;
  assign n30 = x10 & ~x11 ;
  assign n31 = x12 & ~x13 ;
  assign n32 = x14 & ~x15 ;
  assign n33 = ~n31 & ~n32 ;
  assign n34 = n30 & ~n33 ;
  assign n35 = ~x10 & x11 ;
  assign n36 = x12 & x13 ;
  assign n37 = x14 & x15 ;
  assign n38 = ~n36 & ~n37 ;
  assign n39 = n35 & ~n38 ;
  assign n40 = ~n19 & ~n39 ;
  assign n41 = ~n34 & n40 ;
  assign n42 = x6 & ~x7 ;
  assign n43 = ~n41 & n42 ;
  assign n44 = ~n29 & ~n43 ;
  assign n45 = ~x5 & ~x7 ;
  assign n46 = n45 ^ x4 ;
  assign n47 = n46 ^ n43 ;
  assign n48 = ~x9 & n17 ;
  assign n49 = x7 & ~n48 ;
  assign n50 = ~x4 & n49 ;
  assign n51 = n50 ^ n44 ;
  assign n52 = n47 & n51 ;
  assign n53 = n52 ^ n50 ;
  assign n54 = n44 & n53 ;
  assign y0 = ~n54 ;
endmodule
