module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
  assign n10 = ~x4 & x5 ;
  assign n11 = ~x6 & ~n10 ;
  assign n12 = x3 & ~x4 ;
  assign n13 = x2 & n12 ;
  assign n14 = x1 & n13 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n11 & ~n15 ;
  assign n17 = ~x0 & ~x8 ;
  assign n18 = x7 & n17 ;
  assign n19 = ~n16 & n18 ;
  assign n20 = x5 ^ x1 ;
  assign n21 = n20 ^ x6 ;
  assign n22 = x3 ^ x2 ;
  assign n23 = x6 ^ x5 ;
  assign n24 = x4 ^ x3 ;
  assign n25 = n24 ^ x3 ;
  assign n26 = ~n23 & ~n25 ;
  assign n27 = n26 ^ x3 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = ~n22 & n28 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = n21 & ~n30 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = x6 & n32 ;
  assign n34 = n33 ^ x6 ;
  assign n35 = n19 & ~n34 ;
  assign y0 = n35 ;
endmodule
