module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 ;
  assign n17 = ~x8 & ~x9 ;
  assign n18 = x5 & ~n17 ;
  assign n19 = x7 & ~x10 ;
  assign n20 = ~x6 & n19 ;
  assign n21 = ~n18 & n20 ;
  assign n22 = x5 ^ x4 ;
  assign n23 = n22 ^ x7 ;
  assign n24 = n23 ^ x6 ;
  assign n25 = n23 ^ x5 ;
  assign n26 = ~n23 & n25 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = ~n24 & ~n27 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = n30 ^ x5 ;
  assign n32 = x7 & n31 ;
  assign n33 = n32 ^ n23 ;
  assign n34 = ~n21 & ~n33 ;
  assign n35 = x5 & ~x7 ;
  assign n36 = x12 & x13 ;
  assign n37 = n36 ^ x7 ;
  assign n38 = x14 & x15 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n37 & n39 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n35 & n41 ;
  assign n43 = n42 ^ x5 ;
  assign n44 = n43 ^ x6 ;
  assign n45 = x10 ^ x7 ;
  assign n46 = n45 ^ x10 ;
  assign n47 = x9 ^ x8 ;
  assign n48 = ~x4 & n47 ;
  assign n49 = n48 ^ x10 ;
  assign n50 = n46 & ~n49 ;
  assign n51 = n50 ^ x10 ;
  assign n52 = n51 ^ n43 ;
  assign n53 = ~n44 & n52 ;
  assign n54 = n53 ^ n50 ;
  assign n55 = n54 ^ x10 ;
  assign n56 = n55 ^ x6 ;
  assign n57 = ~n43 & ~n56 ;
  assign n58 = n57 ^ n43 ;
  assign n59 = n34 & n58 ;
  assign y0 = ~n59 ;
endmodule
