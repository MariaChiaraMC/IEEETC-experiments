module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 ;
  assign n17 = x11 & x15 ;
  assign n18 = ~x4 & x6 ;
  assign n19 = n17 & n18 ;
  assign n20 = ~x4 & x15 ;
  assign n21 = ~x6 & n20 ;
  assign n22 = ~x4 & ~n17 ;
  assign n24 = x0 & x7 ;
  assign n25 = x8 & x12 ;
  assign n26 = ~n24 & ~n25 ;
  assign n27 = x1 & ~n26 ;
  assign n28 = x9 & x13 ;
  assign n29 = ~n27 & ~n28 ;
  assign n30 = x2 & ~n29 ;
  assign n31 = x10 & x14 ;
  assign n32 = ~n30 & ~n31 ;
  assign n23 = x15 ^ x11 ;
  assign n33 = n32 ^ n23 ;
  assign n34 = ~n22 & ~n33 ;
  assign n35 = ~n21 & ~n34 ;
  assign n36 = n35 ^ x5 ;
  assign n37 = n36 ^ n35 ;
  assign n39 = x3 & x4 ;
  assign n38 = ~n20 & n23 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = ~x6 & n40 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = n42 ^ n35 ;
  assign n44 = ~n37 & ~n43 ;
  assign n45 = n44 ^ n35 ;
  assign n46 = ~n19 & n45 ;
  assign y0 = ~n46 ;
endmodule
