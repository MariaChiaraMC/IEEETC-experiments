module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 ;
  assign n14 = x1 & ~x5 ;
  assign n15 = n14 ^ x1 ;
  assign n16 = n15 ^ x1 ;
  assign n12 = x3 ^ x1 ;
  assign n13 = n12 ^ x1 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = x4 & ~x5 ;
  assign n19 = n18 ^ x1 ;
  assign n20 = n19 ^ x1 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = ~n16 & n21 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = n17 & ~n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n25 ^ x1 ;
  assign n27 = n26 ^ n16 ;
  assign n28 = x2 & ~n27 ;
  assign n29 = n28 ^ x1 ;
  assign n30 = ~x6 & n29 ;
  assign n31 = ~x9 & ~n30 ;
  assign n35 = x0 & ~x7 ;
  assign n36 = ~x10 & n35 ;
  assign n32 = ~x5 & x10 ;
  assign n33 = ~x3 & n32 ;
  assign n34 = ~x4 & n33 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = x1 & n37 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n31 & n39 ;
  assign n41 = ~x3 & x9 ;
  assign n42 = x1 & x6 ;
  assign n43 = x5 ^ x4 ;
  assign n44 = x10 ^ x5 ;
  assign n45 = n43 & n44 ;
  assign n46 = n42 & n45 ;
  assign n47 = n41 & n46 ;
  assign n48 = ~n40 & ~n47 ;
  assign n49 = ~x8 & ~n48 ;
  assign n58 = ~x5 & x9 ;
  assign n64 = x5 & x10 ;
  assign n65 = ~n58 & ~n64 ;
  assign n53 = ~x9 & ~x10 ;
  assign n115 = x3 & ~n53 ;
  assign n116 = n65 & n115 ;
  assign n117 = ~x4 & ~n116 ;
  assign n51 = ~x1 & n35 ;
  assign n52 = ~x8 & ~n51 ;
  assign n54 = x5 & n53 ;
  assign n55 = ~x3 & n54 ;
  assign n56 = ~n52 & n55 ;
  assign n57 = ~x1 & ~x10 ;
  assign n50 = x8 ^ x3 ;
  assign n59 = ~n50 & n58 ;
  assign n60 = ~n57 & n59 ;
  assign n61 = ~n56 & ~n60 ;
  assign n66 = n65 ^ n61 ;
  assign n67 = n66 ^ n61 ;
  assign n62 = n61 ^ n50 ;
  assign n63 = n62 ^ n61 ;
  assign n68 = n67 ^ n63 ;
  assign n69 = ~x1 & n32 ;
  assign n70 = n51 ^ n14 ;
  assign n71 = ~x8 & n70 ;
  assign n72 = n71 ^ n14 ;
  assign n73 = ~n69 & ~n72 ;
  assign n74 = ~x9 & n73 ;
  assign n75 = n74 ^ n61 ;
  assign n76 = n75 ^ n61 ;
  assign n77 = n76 ^ n67 ;
  assign n78 = n67 & ~n77 ;
  assign n79 = n78 ^ n67 ;
  assign n80 = ~n68 & n79 ;
  assign n81 = n80 ^ n78 ;
  assign n82 = n81 ^ n61 ;
  assign n83 = n82 ^ n67 ;
  assign n84 = ~x4 & ~n83 ;
  assign n85 = n84 ^ n61 ;
  assign n86 = n85 ^ x1 ;
  assign n87 = n86 ^ x2 ;
  assign n100 = n87 ^ n86 ;
  assign n89 = ~x5 & ~x10 ;
  assign n90 = x8 & n89 ;
  assign n91 = ~x2 & n90 ;
  assign n92 = ~n64 & ~n91 ;
  assign n93 = x9 ^ x4 ;
  assign n94 = ~n50 & ~n93 ;
  assign n95 = ~n92 & n94 ;
  assign n88 = n87 ^ n85 ;
  assign n96 = n95 ^ n88 ;
  assign n97 = n95 ^ n87 ;
  assign n98 = n97 ^ n86 ;
  assign n99 = n96 & ~n98 ;
  assign n101 = n100 ^ n99 ;
  assign n102 = ~x10 & n18 ;
  assign n103 = n41 & n102 ;
  assign n104 = ~x8 & n103 ;
  assign n105 = n104 ^ n87 ;
  assign n106 = n100 & ~n105 ;
  assign n107 = n106 ^ n104 ;
  assign n108 = n101 & n107 ;
  assign n109 = n108 ^ n99 ;
  assign n110 = n109 ^ n87 ;
  assign n111 = n110 ^ x1 ;
  assign n112 = n111 ^ n86 ;
  assign n118 = n117 ^ n112 ;
  assign n119 = n118 ^ n112 ;
  assign n113 = n112 ^ x1 ;
  assign n114 = n113 ^ n112 ;
  assign n120 = n119 ^ n114 ;
  assign n121 = x4 & ~n32 ;
  assign n122 = n121 ^ n54 ;
  assign n123 = n122 ^ n54 ;
  assign n124 = x4 & ~x9 ;
  assign n125 = n124 ^ n54 ;
  assign n126 = n125 ^ n54 ;
  assign n127 = ~n123 & ~n126 ;
  assign n128 = n127 ^ n54 ;
  assign n129 = x3 & n128 ;
  assign n130 = n129 ^ n54 ;
  assign n131 = x8 & n130 ;
  assign n132 = n131 ^ n112 ;
  assign n133 = n132 ^ n112 ;
  assign n134 = n133 ^ n119 ;
  assign n135 = ~n119 & ~n134 ;
  assign n136 = n135 ^ n119 ;
  assign n137 = ~n120 & ~n136 ;
  assign n138 = n137 ^ n135 ;
  assign n139 = n138 ^ n112 ;
  assign n140 = n139 ^ n119 ;
  assign n141 = x6 & ~n140 ;
  assign n142 = n141 ^ n112 ;
  assign n143 = ~n49 & ~n142 ;
  assign y0 = ~n143 ;
endmodule
