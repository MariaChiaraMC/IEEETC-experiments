// Benchmark "./pla/f51m.pla_7" written by ABC on Mon Apr 20 15:44:01 2020

module \./pla/f51m.pla_7  ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z0  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z0;
  assign z0 = ~x7;
endmodule


