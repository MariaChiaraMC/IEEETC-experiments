module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 ;
  assign n13 = x0 & x5 ;
  assign n14 = ~x11 & n13 ;
  assign n15 = ~x6 & n14 ;
  assign n16 = x1 & n15 ;
  assign n17 = ~x8 & x9 ;
  assign n21 = ~x2 & x3 ;
  assign n22 = x9 & ~n21 ;
  assign n23 = ~x4 & ~n22 ;
  assign n18 = x3 & x4 ;
  assign n19 = ~x2 & ~x7 ;
  assign n20 = ~n18 & n19 ;
  assign n24 = n23 ^ n20 ;
  assign n25 = n24 ^ n20 ;
  assign n26 = x4 & x8 ;
  assign n27 = x3 & ~n26 ;
  assign n28 = n27 ^ x2 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = x4 & x10 ;
  assign n31 = x9 & ~n30 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = ~n29 & n32 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = x7 & n34 ;
  assign n36 = n35 ^ n20 ;
  assign n37 = n36 ^ n20 ;
  assign n38 = ~n25 & n37 ;
  assign n39 = n38 ^ n20 ;
  assign n40 = ~n17 & n39 ;
  assign n41 = n40 ^ n20 ;
  assign n42 = n16 & n41 ;
  assign y0 = n42 ;
endmodule
