module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 ;
  assign n9 = ~x0 & ~x1 ;
  assign n25 = ~x2 & ~x5 ;
  assign n26 = ~x7 & n25 ;
  assign n27 = x3 & ~n26 ;
  assign n10 = x5 ^ x3 ;
  assign n11 = x3 ^ x2 ;
  assign n12 = n11 ^ x5 ;
  assign n13 = n12 ^ x5 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n12 ^ x6 ;
  assign n16 = ~n14 & ~n15 ;
  assign n17 = n16 ^ n12 ;
  assign n18 = ~x7 & n12 ;
  assign n19 = n18 ^ n10 ;
  assign n20 = n17 & n19 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n10 & n21 ;
  assign n23 = n22 ^ n12 ;
  assign n24 = n23 ^ n10 ;
  assign n28 = n27 ^ n24 ;
  assign n29 = n28 ^ x4 ;
  assign n42 = n29 ^ n28 ;
  assign n30 = ~x3 & ~n25 ;
  assign n31 = ~x5 & ~x6 ;
  assign n32 = n31 ^ x2 ;
  assign n33 = ~x7 & ~n32 ;
  assign n34 = n33 ^ x2 ;
  assign n35 = n30 & n34 ;
  assign n36 = n35 ^ n29 ;
  assign n37 = n36 ^ n28 ;
  assign n38 = n29 ^ n24 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n39 ^ n37 ;
  assign n41 = n37 & n40 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = n43 ^ n37 ;
  assign n45 = n28 ^ x6 ;
  assign n46 = n41 ^ n37 ;
  assign n47 = n45 & n46 ;
  assign n48 = n47 ^ n28 ;
  assign n49 = ~n44 & n48 ;
  assign n50 = n49 ^ n28 ;
  assign n51 = n50 ^ n27 ;
  assign n52 = n51 ^ n28 ;
  assign n53 = n9 & ~n52 ;
  assign y0 = n53 ;
endmodule
