module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n11 = x5 ^ x0 ;
  assign n12 = x2 & x3 ;
  assign n13 = x1 & n12 ;
  assign n14 = ~x7 & ~n13 ;
  assign n15 = ~x8 & ~x9 ;
  assign n16 = ~n14 & n15 ;
  assign n17 = ~x6 & n16 ;
  assign n18 = n17 ^ x4 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = x6 & ~x7 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n19 & n21 ;
  assign n23 = n22 ^ n17 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n11 & ~n24 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = n26 ^ n17 ;
  assign n28 = n27 ^ x0 ;
  assign n29 = ~x5 & ~n28 ;
  assign n30 = n29 ^ x5 ;
  assign y0 = ~n30 ;
endmodule
