module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 ;
  assign n7 = x0 & ~x3 ;
  assign n8 = ~x4 & ~n7 ;
  assign n9 = x2 & ~n8 ;
  assign n10 = x5 ^ x2 ;
  assign n15 = n10 ^ x4 ;
  assign n12 = x5 ^ x0 ;
  assign n16 = n15 ^ n12 ;
  assign n11 = n10 ^ x1 ;
  assign n13 = n12 ^ n11 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = n18 ^ n12 ;
  assign n14 = n13 ^ n12 ;
  assign n20 = n19 ^ n14 ;
  assign n21 = n20 ^ n10 ;
  assign n24 = n19 ^ n10 ;
  assign n22 = n17 ^ n13 ;
  assign n23 = n22 ^ n19 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = ~n21 & ~n26 ;
  assign n28 = n27 ^ n19 ;
  assign n29 = n28 ^ n21 ;
  assign n30 = n12 ^ x3 ;
  assign n31 = n30 ^ n10 ;
  assign n32 = n31 ^ n19 ;
  assign n33 = n32 ^ n24 ;
  assign n34 = n22 ^ n17 ;
  assign n39 = n34 ^ n24 ;
  assign n40 = n39 ^ n21 ;
  assign n41 = ~n24 & n40 ;
  assign n35 = n34 ^ n19 ;
  assign n36 = n35 ^ n21 ;
  assign n37 = n35 ^ n24 ;
  assign n38 = n36 & n37 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = n42 ^ n22 ;
  assign n44 = n43 ^ n31 ;
  assign n45 = n44 ^ n19 ;
  assign n46 = n45 ^ n24 ;
  assign n47 = n46 ^ n21 ;
  assign n48 = ~n33 & n47 ;
  assign n49 = n48 ^ n38 ;
  assign n50 = n49 ^ n31 ;
  assign n51 = n50 ^ n24 ;
  assign n52 = n51 ^ n21 ;
  assign n53 = n29 & ~n52 ;
  assign n54 = n53 ^ n38 ;
  assign n55 = n54 ^ n17 ;
  assign n56 = n55 ^ n22 ;
  assign n57 = n56 ^ n19 ;
  assign n58 = n57 ^ n21 ;
  assign n59 = n58 ^ x5 ;
  assign n60 = n59 ^ n13 ;
  assign n61 = ~n9 & ~n60 ;
  assign y0 = ~n61 ;
endmodule
