module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 ;
  assign n22 = ~x0 & ~x1 ;
  assign n23 = ~x4 & ~n22 ;
  assign n24 = ~x0 & ~x2 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = ~x2 & ~x3 ;
  assign n28 = ~x1 & ~n27 ;
  assign n29 = n28 ^ x3 ;
  assign n30 = x5 & n29 ;
  assign n31 = n30 ^ x3 ;
  assign n32 = n26 & ~n31 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ x3 ;
  assign n35 = n34 ^ x5 ;
  assign n36 = n23 & ~n35 ;
  assign n37 = ~x19 & ~x20 ;
  assign n38 = n37 ^ x18 ;
  assign n39 = n38 ^ x18 ;
  assign n40 = ~x3 & n24 ;
  assign n41 = ~x6 & ~x7 ;
  assign n42 = x12 & ~x13 ;
  assign n43 = n41 & ~n42 ;
  assign n44 = ~x13 & ~n43 ;
  assign n45 = ~x9 & ~x10 ;
  assign n46 = ~x8 & ~x11 ;
  assign n47 = ~n45 & n46 ;
  assign n48 = ~x13 & n47 ;
  assign n49 = n48 ^ x5 ;
  assign n50 = n49 ^ n44 ;
  assign n56 = ~x10 & x11 ;
  assign n57 = ~x8 & ~x9 ;
  assign n58 = n56 & n57 ;
  assign n51 = ~x9 & ~n22 ;
  assign n52 = ~x1 & x3 ;
  assign n53 = ~x2 & n52 ;
  assign n54 = ~n24 & ~n53 ;
  assign n55 = ~n51 & ~n54 ;
  assign n59 = n58 ^ n55 ;
  assign n60 = n48 & ~n59 ;
  assign n61 = n60 ^ n58 ;
  assign n62 = ~n50 & n61 ;
  assign n63 = n62 ^ n60 ;
  assign n64 = n63 ^ n58 ;
  assign n65 = n64 ^ n48 ;
  assign n66 = ~n44 & n65 ;
  assign n67 = ~n40 & ~n66 ;
  assign n68 = ~x12 & ~x13 ;
  assign n69 = x9 & n68 ;
  assign n80 = n41 & n56 ;
  assign n81 = ~n24 & ~n52 ;
  assign n82 = n80 & ~n81 ;
  assign n70 = x8 ^ x5 ;
  assign n72 = n70 ^ x2 ;
  assign n71 = n70 ^ x8 ;
  assign n73 = n72 ^ n71 ;
  assign n83 = n82 ^ n73 ;
  assign n87 = n83 ^ n72 ;
  assign n88 = n87 ^ n70 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = n74 ^ n70 ;
  assign n76 = n75 ^ n70 ;
  assign n77 = n72 ^ n53 ;
  assign n78 = n77 ^ n70 ;
  assign n79 = ~n76 & ~n78 ;
  assign n84 = n83 ^ n79 ;
  assign n85 = n84 ^ n70 ;
  assign n86 = ~n75 & ~n85 ;
  assign n89 = n88 ^ n86 ;
  assign n90 = n89 ^ n75 ;
  assign n91 = x10 & ~x11 ;
  assign n92 = n91 ^ n70 ;
  assign n93 = n88 ^ n85 ;
  assign n94 = n93 ^ n75 ;
  assign n95 = ~n92 & ~n94 ;
  assign n96 = n95 ^ n70 ;
  assign n97 = n90 & n96 ;
  assign n98 = n97 ^ n95 ;
  assign n99 = n98 ^ n70 ;
  assign n100 = n99 ^ x8 ;
  assign n101 = n69 & n100 ;
  assign n102 = n67 & ~n101 ;
  assign n103 = ~x4 & ~n102 ;
  assign n104 = x2 & n58 ;
  assign n105 = ~x4 & ~n104 ;
  assign n106 = x0 & ~n105 ;
  assign n107 = x11 & ~x12 ;
  assign n108 = ~x8 & x9 ;
  assign n109 = n107 & n108 ;
  assign n110 = x5 & n109 ;
  assign n111 = ~n106 & ~n110 ;
  assign n112 = ~x1 & ~n111 ;
  assign n113 = ~x11 & n108 ;
  assign n114 = ~x10 & n113 ;
  assign n115 = ~x15 & x16 ;
  assign n116 = n115 ^ x12 ;
  assign n117 = x2 & n116 ;
  assign n118 = n117 ^ x12 ;
  assign n119 = ~n114 & n118 ;
  assign n120 = x13 & ~n119 ;
  assign n121 = x11 ^ x10 ;
  assign n122 = x16 ^ x8 ;
  assign n123 = n122 ^ x17 ;
  assign n124 = n121 & ~n123 ;
  assign n125 = n124 ^ n121 ;
  assign n126 = x16 ^ x11 ;
  assign n127 = n126 ^ n124 ;
  assign n128 = n122 & ~n127 ;
  assign n129 = n128 ^ n122 ;
  assign n130 = n129 ^ x17 ;
  assign n131 = n125 & ~n130 ;
  assign n132 = n43 & n131 ;
  assign n133 = x2 & ~n132 ;
  assign n134 = x10 & n107 ;
  assign n135 = ~x2 & ~n134 ;
  assign n136 = x9 & ~n135 ;
  assign n137 = x0 & ~x13 ;
  assign n138 = x1 & ~n137 ;
  assign n139 = ~n136 & ~n138 ;
  assign n140 = x4 & n139 ;
  assign n141 = ~n133 & n140 ;
  assign n142 = ~n120 & n141 ;
  assign n143 = x5 & ~n142 ;
  assign n144 = ~n22 & ~n27 ;
  assign n145 = ~x4 & n68 ;
  assign n148 = n47 ^ n41 ;
  assign n157 = n148 ^ n47 ;
  assign n146 = x8 & x9 ;
  assign n147 = n146 ^ n47 ;
  assign n149 = n148 ^ n147 ;
  assign n150 = n149 ^ n148 ;
  assign n151 = n150 ^ n47 ;
  assign n152 = n149 ^ x11 ;
  assign n153 = n152 ^ x10 ;
  assign n154 = n153 ^ n149 ;
  assign n155 = n154 ^ n151 ;
  assign n156 = n151 & n155 ;
  assign n158 = n157 ^ n156 ;
  assign n159 = n158 ^ n151 ;
  assign n160 = n47 ^ x10 ;
  assign n161 = n156 ^ n151 ;
  assign n162 = ~n160 & n161 ;
  assign n163 = n162 ^ n47 ;
  assign n164 = n159 & ~n163 ;
  assign n165 = n164 ^ n47 ;
  assign n166 = n165 ^ n41 ;
  assign n167 = n166 ^ n47 ;
  assign n168 = n145 & n167 ;
  assign n169 = n144 & n168 ;
  assign n170 = ~n143 & ~n169 ;
  assign n171 = ~n112 & n170 ;
  assign n172 = ~x3 & ~n171 ;
  assign n173 = ~x0 & x4 ;
  assign n174 = ~x5 & ~n173 ;
  assign n175 = x1 & x2 ;
  assign n176 = ~n174 & n175 ;
  assign n177 = n53 ^ x5 ;
  assign n178 = n177 ^ n53 ;
  assign n179 = x3 & x4 ;
  assign n180 = n144 & n179 ;
  assign n181 = n180 ^ n53 ;
  assign n182 = ~n178 & n181 ;
  assign n183 = n182 ^ n53 ;
  assign n184 = ~n176 & ~n183 ;
  assign n185 = ~n172 & n184 ;
  assign n186 = ~n103 & n185 ;
  assign n187 = n186 ^ x18 ;
  assign n188 = n39 & n187 ;
  assign n189 = n188 ^ x18 ;
  assign n190 = x14 & n189 ;
  assign n191 = ~n36 & n190 ;
  assign y0 = ~n191 ;
endmodule
