module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 ;
  assign n20 = ~x11 & ~x14 ;
  assign n21 = x3 & ~x5 ;
  assign n22 = ~x10 & n21 ;
  assign n23 = x1 & ~x12 ;
  assign n24 = ~n22 & n23 ;
  assign n25 = n20 & n24 ;
  assign n26 = ~x18 & ~n25 ;
  assign n27 = ~x16 & ~x17 ;
  assign n28 = ~x0 & n27 ;
  assign n29 = ~n26 & n28 ;
  assign n30 = ~x6 & ~x7 ;
  assign n31 = x8 & x9 ;
  assign n32 = n30 & ~n31 ;
  assign n33 = x4 & n32 ;
  assign n34 = ~x14 & x18 ;
  assign n35 = ~x3 & n34 ;
  assign n36 = ~x15 & n35 ;
  assign n37 = ~n33 & n36 ;
  assign n38 = n29 & ~n37 ;
  assign n39 = x15 ^ x14 ;
  assign n40 = ~x8 & n30 ;
  assign n41 = n40 ^ x15 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = n42 ^ n39 ;
  assign n44 = ~x10 & n32 ;
  assign n45 = ~x2 & n44 ;
  assign n46 = n45 ^ x18 ;
  assign n47 = ~n45 & ~n46 ;
  assign n48 = n47 ^ n40 ;
  assign n49 = n48 ^ n45 ;
  assign n50 = n43 & ~n49 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = n51 ^ n45 ;
  assign n53 = n39 & ~n52 ;
  assign n54 = n53 ^ x15 ;
  assign n55 = n38 & ~n54 ;
  assign y0 = n55 ;
endmodule
