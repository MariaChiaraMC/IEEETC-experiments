module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 ;
  assign n20 = ~x0 & ~x14 ;
  assign n21 = x4 & ~x9 ;
  assign n22 = x16 & ~x18 ;
  assign n23 = x7 & x8 ;
  assign n24 = n22 & n23 ;
  assign n25 = ~x6 & n24 ;
  assign n26 = ~x8 & x18 ;
  assign n27 = ~x7 & n26 ;
  assign n28 = x16 ^ x6 ;
  assign n29 = n27 & ~n28 ;
  assign n30 = ~n25 & ~n29 ;
  assign n31 = n21 & ~n30 ;
  assign n32 = x1 & ~x16 ;
  assign n33 = x3 & ~x5 ;
  assign n34 = ~x10 & n33 ;
  assign n35 = x11 & x12 ;
  assign n36 = x13 & n35 ;
  assign n37 = ~n34 & ~n36 ;
  assign n38 = n32 & n37 ;
  assign n39 = ~x18 & n38 ;
  assign n40 = ~x15 & ~n39 ;
  assign n41 = ~n31 & n40 ;
  assign n42 = x6 & x16 ;
  assign n43 = ~x18 & ~n42 ;
  assign n44 = x7 & ~n43 ;
  assign n46 = n22 & ~n23 ;
  assign n45 = ~x16 & x18 ;
  assign n47 = n46 ^ n45 ;
  assign n48 = n45 ^ x6 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = x8 ^ x6 ;
  assign n51 = x9 ^ x6 ;
  assign n52 = n51 ^ n50 ;
  assign n53 = n50 & n52 ;
  assign n54 = n53 ^ x6 ;
  assign n55 = n54 ^ n50 ;
  assign n56 = n49 & n55 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n57 ^ n50 ;
  assign n59 = n47 & n58 ;
  assign n60 = n59 ^ n46 ;
  assign n61 = x15 & ~n60 ;
  assign n62 = ~n44 & n61 ;
  assign n63 = ~n41 & ~n62 ;
  assign n64 = x18 ^ x16 ;
  assign n65 = x3 ^ x2 ;
  assign n66 = n65 ^ x3 ;
  assign n67 = x10 ^ x3 ;
  assign n68 = n67 ^ x3 ;
  assign n69 = ~n66 & ~n68 ;
  assign n70 = n69 ^ x3 ;
  assign n71 = x15 & ~n70 ;
  assign n72 = n71 ^ x3 ;
  assign n73 = n64 & n72 ;
  assign n74 = ~x17 & ~n73 ;
  assign n75 = ~n63 & n74 ;
  assign n76 = x8 & ~x18 ;
  assign n77 = ~x7 & n76 ;
  assign n78 = x7 & n26 ;
  assign n79 = ~n77 & ~n78 ;
  assign n80 = ~x15 & ~n28 ;
  assign n81 = n21 & n80 ;
  assign n82 = ~n79 & n81 ;
  assign n83 = x18 ^ x8 ;
  assign n84 = x8 ^ x7 ;
  assign n85 = n84 ^ x9 ;
  assign n86 = n85 ^ n84 ;
  assign n87 = n84 ^ x18 ;
  assign n88 = ~n86 & n87 ;
  assign n89 = n88 ^ n84 ;
  assign n90 = ~n83 & n89 ;
  assign n91 = n90 ^ n84 ;
  assign n92 = x16 & x18 ;
  assign n93 = n28 & ~n92 ;
  assign n94 = n91 & ~n93 ;
  assign n95 = x15 & ~n94 ;
  assign n96 = x17 & ~n95 ;
  assign n97 = ~n82 & n96 ;
  assign n98 = ~n75 & ~n97 ;
  assign n99 = n92 ^ n72 ;
  assign n100 = n92 ^ x17 ;
  assign n101 = n100 ^ x17 ;
  assign n102 = n101 ^ n99 ;
  assign n103 = x8 & x9 ;
  assign n104 = x6 & ~n103 ;
  assign n105 = n104 ^ x15 ;
  assign n106 = x15 & ~n105 ;
  assign n107 = n106 ^ x17 ;
  assign n108 = n107 ^ x15 ;
  assign n109 = n102 & ~n108 ;
  assign n110 = n109 ^ n106 ;
  assign n111 = n110 ^ x15 ;
  assign n112 = n99 & n111 ;
  assign n113 = n112 ^ n72 ;
  assign n114 = ~n98 & ~n113 ;
  assign n115 = n20 & ~n114 ;
  assign y0 = n115 ;
endmodule
