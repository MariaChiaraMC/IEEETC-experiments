module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;
  assign n9 = x3 ^ x2 ;
  assign n10 = n9 ^ x0 ;
  assign n11 = n10 ^ x4 ;
  assign n13 = x4 ^ x3 ;
  assign n16 = n11 & n13 ;
  assign n7 = x4 ^ x0 ;
  assign n8 = n7 ^ x0 ;
  assign n12 = n11 ^ x0 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n8 & ~n14 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n13 ^ x5 ;
  assign n19 = n15 & n18 ;
  assign n20 = n17 & n19 ;
  assign n21 = n20 ^ n15 ;
  assign n22 = n21 ^ n16 ;
  assign n23 = n22 ^ n9 ;
  assign n24 = x1 & ~n23 ;
  assign n25 = x0 & x4 ;
  assign n26 = x2 & ~x3 ;
  assign n27 = n25 & n26 ;
  assign n28 = x5 & n27 ;
  assign n29 = x3 ^ x0 ;
  assign n30 = x4 ^ x2 ;
  assign n31 = n30 ^ x2 ;
  assign n32 = x2 ^ x1 ;
  assign n33 = ~n31 & n32 ;
  assign n34 = n33 ^ x2 ;
  assign n35 = n34 ^ x3 ;
  assign n36 = n29 & ~n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ x2 ;
  assign n39 = n38 ^ x0 ;
  assign n40 = x3 & ~n39 ;
  assign n41 = n40 ^ x3 ;
  assign n42 = ~n28 & ~n41 ;
  assign n43 = ~n24 & n42 ;
  assign y0 = ~n43 ;
endmodule
