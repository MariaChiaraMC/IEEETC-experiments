module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n17 = ~x7 & ~x10 ;
  assign n18 = ~x2 & ~x14 ;
  assign n19 = ~x4 & ~x6 ;
  assign n20 = n18 & n19 ;
  assign n21 = x5 & ~x11 ;
  assign n22 = ~x9 & ~x12 ;
  assign n23 = n21 & n22 ;
  assign n24 = ~x3 & ~x15 ;
  assign n25 = ~x8 & ~x13 ;
  assign n26 = n24 & n25 ;
  assign n27 = n23 & n26 ;
  assign n28 = n20 & n27 ;
  assign n29 = n17 & n28 ;
  assign n30 = x1 & ~n29 ;
  assign y0 = ~n30 ;
endmodule
