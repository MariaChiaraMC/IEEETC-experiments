// Benchmark "./newcond.pla" written by ABC on Thu Apr 23 10:59:57 2020

module \./newcond.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10,
    z1  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10;
  output z1;
  assign z1 = 1'b1;
endmodule


