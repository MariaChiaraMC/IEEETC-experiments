module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 ;
  assign n11 = x4 & ~x5 ;
  assign n12 = x3 & x6 ;
  assign n13 = x2 & ~x9 ;
  assign n14 = n12 & n13 ;
  assign n15 = ~x3 & x7 ;
  assign n16 = ~x2 & ~x8 ;
  assign n17 = n15 & n16 ;
  assign n18 = ~x8 & ~x9 ;
  assign n19 = ~x3 & x8 ;
  assign n20 = x3 & x9 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = n21 ^ x0 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = x2 & ~x3 ;
  assign n25 = ~x2 & x3 ;
  assign n26 = ~n24 & ~n25 ;
  assign n27 = n26 ^ n21 ;
  assign n28 = n23 & n27 ;
  assign n29 = n28 ^ n21 ;
  assign n30 = ~n18 & ~n29 ;
  assign n31 = x1 & ~n30 ;
  assign n32 = ~n17 & ~n31 ;
  assign n33 = ~n14 & n32 ;
  assign n34 = n11 & ~n33 ;
  assign n35 = ~x2 & ~x7 ;
  assign n36 = n19 & n35 ;
  assign n37 = x2 & ~x6 ;
  assign n38 = n20 & n37 ;
  assign n39 = ~n36 & ~n38 ;
  assign n40 = x0 & ~n39 ;
  assign n41 = ~n34 & ~n40 ;
  assign n42 = x0 & x8 ;
  assign n43 = x9 & n42 ;
  assign n44 = ~n35 & ~n37 ;
  assign n45 = ~x0 & ~x5 ;
  assign n46 = ~n44 & n45 ;
  assign n47 = n46 ^ n21 ;
  assign n48 = n11 & ~n21 ;
  assign n49 = ~n47 & n48 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = ~n43 & n50 ;
  assign n52 = n51 ^ x1 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = ~x7 & n24 ;
  assign n55 = x0 & n54 ;
  assign n56 = x9 & n55 ;
  assign n59 = ~x6 & n25 ;
  assign n57 = ~x6 & ~x7 ;
  assign n58 = ~x4 & ~n57 ;
  assign n60 = n59 ^ n58 ;
  assign n61 = n58 ^ n54 ;
  assign n62 = n61 ^ n54 ;
  assign n63 = n54 ^ n42 ;
  assign n64 = ~n62 & ~n63 ;
  assign n65 = n64 ^ n54 ;
  assign n66 = n60 & n65 ;
  assign n67 = n66 ^ n59 ;
  assign n86 = ~n12 & ~n15 ;
  assign n68 = ~n26 & n46 ;
  assign n69 = x3 ^ x2 ;
  assign n70 = n69 ^ x0 ;
  assign n71 = x9 ^ x8 ;
  assign n72 = x8 ^ x3 ;
  assign n73 = n72 ^ x8 ;
  assign n74 = n71 & ~n73 ;
  assign n75 = n74 ^ x8 ;
  assign n76 = n75 ^ n69 ;
  assign n77 = n70 & ~n76 ;
  assign n78 = n77 ^ n74 ;
  assign n79 = n78 ^ x8 ;
  assign n80 = n79 ^ x0 ;
  assign n81 = n69 & ~n80 ;
  assign n82 = n81 ^ n69 ;
  assign n83 = n82 ^ x0 ;
  assign n84 = n11 & ~n83 ;
  assign n85 = ~n68 & ~n84 ;
  assign n87 = n86 ^ n85 ;
  assign n88 = n87 ^ n85 ;
  assign n89 = ~n11 & ~n45 ;
  assign n90 = n89 ^ n85 ;
  assign n91 = n88 & ~n90 ;
  assign n92 = n91 ^ n85 ;
  assign n93 = ~n67 & n92 ;
  assign n94 = ~n56 & n93 ;
  assign n95 = n94 ^ n51 ;
  assign n96 = ~n53 & n95 ;
  assign n97 = n96 ^ n51 ;
  assign n98 = n41 & n97 ;
  assign y0 = ~n98 ;
endmodule
