module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 ;
  assign n9 = ~x0 & ~x1 ;
  assign n10 = x4 ^ x3 ;
  assign n11 = n10 ^ x5 ;
  assign n15 = n11 ^ x5 ;
  assign n16 = n15 ^ x6 ;
  assign n17 = n16 ^ n11 ;
  assign n12 = x5 ^ x4 ;
  assign n20 = n12 ^ x6 ;
  assign n21 = n20 ^ x7 ;
  assign n28 = n21 ^ n11 ;
  assign n29 = n28 ^ n17 ;
  assign n30 = n17 & n29 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n13 ^ n11 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = n16 ^ x7 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ n11 ;
  assign n24 = n23 ^ n18 ;
  assign n25 = n18 & n24 ;
  assign n35 = n30 ^ n25 ;
  assign n26 = n25 ^ n13 ;
  assign n27 = n26 ^ n18 ;
  assign n31 = n30 ^ n13 ;
  assign n32 = n31 ^ n17 ;
  assign n33 = n32 ^ x2 ;
  assign n34 = n27 & n33 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = x2 & n36 ;
  assign n38 = n37 ^ n30 ;
  assign n39 = n38 ^ n25 ;
  assign n40 = n39 ^ n34 ;
  assign n41 = n40 ^ x2 ;
  assign n42 = n41 ^ x3 ;
  assign n43 = n42 ^ x2 ;
  assign n44 = n9 & ~n43 ;
  assign y0 = n44 ;
endmodule
