// Benchmark "./bcd.div3.pla" written by ABC on Thu Apr 23 10:59:48 2020

module \./bcd.div3.pla  ( 
    x0, x1, x2, x3,
    z2  );
  input  x0, x1, x2, x3;
  output z2;
  assign z2 = 1'b1;
endmodule


