module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n9 = ~x4 & x5 ;
  assign n10 = n9 ^ x3 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = ~x4 & x6 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = n13 ^ n9 ;
  assign n15 = n11 & n14 ;
  assign n16 = n15 ^ n9 ;
  assign n17 = x0 & ~n16 ;
  assign n18 = n17 ^ n9 ;
  assign n19 = x2 ^ x1 ;
  assign n28 = n19 ^ x1 ;
  assign n20 = x1 & ~x5 ;
  assign n21 = x7 & ~n20 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ x1 ;
  assign n24 = n21 ^ n12 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n23 & n26 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = x1 ^ x0 ;
  assign n32 = n27 ^ n23 ;
  assign n33 = ~n31 & n32 ;
  assign n34 = n33 ^ x1 ;
  assign n35 = n30 & n34 ;
  assign n36 = n35 ^ x1 ;
  assign n37 = n36 ^ x1 ;
  assign n38 = ~n18 & n37 ;
  assign y0 = ~n38 ;
endmodule
