module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 ;
  assign n10 = x4 ^ x2 ;
  assign n11 = n10 ^ x4 ;
  assign n12 = n11 ^ x1 ;
  assign n8 = x4 ^ x3 ;
  assign n9 = n8 ^ x1 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = n12 ^ x1 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n12 ^ x5 ;
  assign n18 = ~n12 & n17 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = n19 ^ n12 ;
  assign n21 = ~n16 & ~n20 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = n22 ^ n12 ;
  assign n24 = ~n14 & ~n23 ;
  assign n25 = n24 ^ n18 ;
  assign n26 = n25 ^ n12 ;
  assign n27 = n26 ^ n10 ;
  assign n28 = x6 & ~n27 ;
  assign n29 = ~x5 & ~x6 ;
  assign n30 = ~x1 & x4 ;
  assign n31 = n29 & n30 ;
  assign n32 = ~x0 & ~n31 ;
  assign n33 = x6 ^ x3 ;
  assign n34 = n33 ^ x6 ;
  assign n35 = n33 ^ x5 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = n37 ^ n33 ;
  assign n44 = n38 ^ n33 ;
  assign n45 = n44 ^ n34 ;
  assign n39 = ~x4 & ~x6 ;
  assign n40 = n39 ^ n33 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n41 ^ n33 ;
  assign n43 = n42 ^ n34 ;
  assign n46 = n45 ^ n43 ;
  assign n47 = ~n34 & n46 ;
  assign n48 = n47 ^ n38 ;
  assign n49 = n48 ^ n45 ;
  assign n50 = ~x2 & ~x4 ;
  assign n54 = n50 ^ n33 ;
  assign n51 = n50 ^ x2 ;
  assign n52 = n45 ^ n38 ;
  assign n53 = n51 & ~n52 ;
  assign n55 = n54 ^ n53 ;
  assign n56 = n55 ^ n51 ;
  assign n57 = n56 ^ n34 ;
  assign n58 = ~n48 & ~n57 ;
  assign n59 = n58 ^ n38 ;
  assign n60 = n59 ^ n34 ;
  assign n61 = n60 ^ n45 ;
  assign n62 = ~n49 & n61 ;
  assign n63 = n62 ^ n38 ;
  assign n64 = n63 ^ n34 ;
  assign n65 = n64 ^ n45 ;
  assign n66 = n65 ^ x6 ;
  assign n67 = x1 & ~n66 ;
  assign n68 = n32 & ~n67 ;
  assign n69 = ~n28 & n68 ;
  assign n70 = x5 ^ x4 ;
  assign n71 = x5 ^ x1 ;
  assign n72 = n71 ^ x1 ;
  assign n73 = x3 & x6 ;
  assign n74 = n73 ^ x1 ;
  assign n75 = n72 & n74 ;
  assign n76 = n75 ^ x1 ;
  assign n77 = ~n70 & n76 ;
  assign n78 = x2 & n77 ;
  assign n79 = x3 & ~x5 ;
  assign n80 = x6 ^ x5 ;
  assign n81 = ~n50 & ~n80 ;
  assign n82 = ~n79 & ~n81 ;
  assign n83 = ~x1 & ~n82 ;
  assign n84 = x5 & x6 ;
  assign n85 = n84 ^ x5 ;
  assign n86 = ~x3 & ~n85 ;
  assign n87 = n86 ^ x5 ;
  assign n88 = n87 ^ x4 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = n89 ^ x1 ;
  assign n91 = n29 ^ x6 ;
  assign n92 = ~x3 & n91 ;
  assign n93 = n92 ^ x6 ;
  assign n94 = n93 ^ x2 ;
  assign n95 = ~x2 & ~n94 ;
  assign n96 = n95 ^ n87 ;
  assign n97 = n96 ^ x2 ;
  assign n98 = n90 & n97 ;
  assign n99 = n98 ^ n95 ;
  assign n100 = n99 ^ x2 ;
  assign n101 = x1 & ~n100 ;
  assign n102 = n101 ^ x1 ;
  assign n103 = ~n83 & ~n102 ;
  assign n104 = ~x2 & ~x3 ;
  assign n105 = n104 ^ n31 ;
  assign n106 = n105 ^ n31 ;
  assign n107 = n84 ^ n31 ;
  assign n108 = n106 & n107 ;
  assign n109 = n108 ^ n31 ;
  assign n110 = x0 & ~n109 ;
  assign n111 = ~n103 & n110 ;
  assign n112 = ~n78 & n111 ;
  assign n113 = ~n69 & ~n112 ;
  assign y0 = n113 ;
endmodule
