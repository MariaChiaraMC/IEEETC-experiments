module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 ;
  assign n9 = ~x6 & x7 ;
  assign n10 = ~x2 & n9 ;
  assign n11 = x0 & ~x7 ;
  assign n12 = x2 & ~n9 ;
  assign n13 = ~n11 & n12 ;
  assign n14 = ~n10 & ~n13 ;
  assign n15 = ~x3 & x4 ;
  assign n16 = ~x0 & x6 ;
  assign n17 = x1 & ~n16 ;
  assign n18 = ~x5 & n17 ;
  assign n19 = n15 & n18 ;
  assign n20 = ~n14 & n19 ;
  assign n21 = x3 ^ x0 ;
  assign n22 = x5 ^ x2 ;
  assign n23 = x7 ^ x6 ;
  assign n24 = x6 ^ x5 ;
  assign n25 = n23 & n24 ;
  assign n26 = n22 & n25 ;
  assign n27 = n26 ^ x3 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = n28 ^ n21 ;
  assign n30 = x5 & x6 ;
  assign n31 = x7 ^ x2 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = n30 & ~n32 ;
  assign n34 = n33 ^ n26 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n29 & n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ n30 ;
  assign n39 = ~n21 & n38 ;
  assign n40 = ~x4 & n39 ;
  assign n41 = ~x1 & n40 ;
  assign n42 = ~n20 & ~n41 ;
  assign y0 = ~n42 ;
endmodule
