module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 ;
  assign n22 = ~x0 & ~x5 ;
  assign n23 = ~x6 & n22 ;
  assign n67 = x7 & ~x8 ;
  assign n68 = x9 & n67 ;
  assign n69 = n23 & n68 ;
  assign n53 = x6 & x7 ;
  assign n11 = x8 & x9 ;
  assign n14 = ~x0 & x5 ;
  assign n70 = n11 & n14 ;
  assign n71 = n53 & n70 ;
  assign n72 = ~x8 & ~x9 ;
  assign n73 = n23 & n72 ;
  assign n74 = ~n71 & ~n73 ;
  assign n75 = x5 & ~x7 ;
  assign n45 = ~x6 & x8 ;
  assign n76 = x9 & n45 ;
  assign n77 = n76 ^ x0 ;
  assign n78 = n77 ^ n76 ;
  assign n79 = n78 ^ n75 ;
  assign n42 = ~x6 & ~x8 ;
  assign n25 = x6 & ~x9 ;
  assign n80 = n42 ^ n25 ;
  assign n81 = ~n42 & n80 ;
  assign n82 = n81 ^ n76 ;
  assign n83 = n82 ^ n42 ;
  assign n84 = n79 & n83 ;
  assign n85 = n84 ^ n81 ;
  assign n86 = n85 ^ n42 ;
  assign n87 = n75 & ~n86 ;
  assign n88 = n87 ^ n75 ;
  assign n89 = n74 & ~n88 ;
  assign n90 = n89 ^ x2 ;
  assign n91 = n90 ^ n89 ;
  assign n92 = n91 ^ n69 ;
  assign n93 = ~x7 & x8 ;
  assign n94 = n25 & n93 ;
  assign n95 = x0 & ~n94 ;
  assign n96 = ~x5 & x8 ;
  assign n97 = ~x6 & x7 ;
  assign n98 = ~n25 & ~n97 ;
  assign n99 = n96 & ~n98 ;
  assign n55 = ~x8 & x9 ;
  assign n100 = n55 & n75 ;
  assign n101 = ~n99 & ~n100 ;
  assign n102 = ~x0 & n101 ;
  assign n103 = n102 ^ n95 ;
  assign n104 = ~n95 & n103 ;
  assign n105 = n104 ^ n89 ;
  assign n106 = n105 ^ n95 ;
  assign n107 = n92 & n106 ;
  assign n108 = n107 ^ n104 ;
  assign n109 = n108 ^ n95 ;
  assign n110 = ~n69 & ~n109 ;
  assign n111 = n110 ^ n69 ;
  assign n112 = ~x1 & n111 ;
  assign n12 = x7 & n11 ;
  assign n13 = ~x2 & n12 ;
  assign n15 = x0 & ~x5 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = ~x6 & n16 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n13 & n18 ;
  assign n31 = x0 & x9 ;
  assign n32 = x5 & n31 ;
  assign n43 = x5 & n42 ;
  assign n44 = x6 & ~x8 ;
  assign n46 = ~n44 & ~n45 ;
  assign n47 = n31 & ~n46 ;
  assign n48 = ~n43 & ~n47 ;
  assign n49 = ~n32 & ~n48 ;
  assign n50 = ~x7 & n49 ;
  assign n20 = x8 & ~x9 ;
  assign n21 = ~x7 & n20 ;
  assign n24 = n21 & n23 ;
  assign n26 = ~x0 & n25 ;
  assign n27 = n26 ^ x7 ;
  assign n28 = n27 ^ x5 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = n29 ^ x8 ;
  assign n33 = n32 ^ x8 ;
  assign n34 = ~x6 & n33 ;
  assign n35 = n34 ^ n26 ;
  assign n36 = n30 & n35 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = x8 & n37 ;
  assign n39 = n38 ^ n34 ;
  assign n40 = n39 ^ n36 ;
  assign n41 = ~n24 & ~n40 ;
  assign n51 = n50 ^ n41 ;
  assign n52 = n51 ^ n41 ;
  assign n54 = x5 & n20 ;
  assign n56 = n22 & n55 ;
  assign n57 = ~n54 & ~n56 ;
  assign n58 = n53 & ~n57 ;
  assign n59 = n58 ^ n41 ;
  assign n60 = n59 ^ n41 ;
  assign n61 = ~n52 & ~n60 ;
  assign n62 = n61 ^ n41 ;
  assign n63 = x2 & n62 ;
  assign n64 = n63 ^ n41 ;
  assign n65 = ~x1 & ~n64 ;
  assign n66 = ~n19 & ~n65 ;
  assign n113 = n112 ^ n66 ;
  assign n114 = n113 ^ x4 ;
  assign n122 = n114 ^ n113 ;
  assign n115 = ~x2 & x4 ;
  assign n116 = n115 ^ n114 ;
  assign n117 = n116 ^ n113 ;
  assign n118 = n114 ^ n66 ;
  assign n119 = n118 ^ n115 ;
  assign n120 = n119 ^ n117 ;
  assign n121 = n117 & n120 ;
  assign n123 = n122 ^ n121 ;
  assign n124 = n123 ^ n117 ;
  assign n125 = ~x7 & ~x9 ;
  assign n126 = x0 & n42 ;
  assign n127 = n125 & n126 ;
  assign n128 = n127 ^ n113 ;
  assign n129 = n121 ^ n117 ;
  assign n130 = ~n128 & n129 ;
  assign n131 = n130 ^ n113 ;
  assign n132 = ~n124 & ~n131 ;
  assign n133 = n132 ^ n113 ;
  assign n134 = n133 ^ n112 ;
  assign n135 = n134 ^ n113 ;
  assign n136 = ~x3 & n135 ;
  assign n137 = x3 & ~x4 ;
  assign n138 = ~x0 & n137 ;
  assign n139 = x5 & n97 ;
  assign n140 = n138 & n139 ;
  assign n141 = n72 ^ n55 ;
  assign n142 = ~x2 & n141 ;
  assign n143 = n142 ^ n72 ;
  assign n144 = n140 & n143 ;
  assign n145 = n144 ^ n136 ;
  assign n146 = x2 & x7 ;
  assign n147 = n137 & n146 ;
  assign n148 = n55 & n147 ;
  assign n149 = x4 & ~x7 ;
  assign n150 = ~x3 & ~n149 ;
  assign n151 = ~x2 & n150 ;
  assign n152 = ~x7 & x9 ;
  assign n153 = n152 ^ x8 ;
  assign n154 = n151 & n153 ;
  assign n155 = ~n148 & ~n154 ;
  assign n156 = n15 & ~n155 ;
  assign n157 = x4 & ~x5 ;
  assign n165 = x2 ^ x0 ;
  assign n160 = x7 ^ x3 ;
  assign n161 = n160 ^ x9 ;
  assign n158 = x8 ^ x7 ;
  assign n159 = n158 ^ x9 ;
  assign n162 = n161 ^ n159 ;
  assign n163 = n162 ^ x7 ;
  assign n164 = n163 ^ x7 ;
  assign n166 = n165 ^ n164 ;
  assign n167 = ~n158 & ~n161 ;
  assign n168 = n167 ^ n163 ;
  assign n169 = n166 & ~n168 ;
  assign n170 = n169 ^ n165 ;
  assign n171 = n170 ^ n166 ;
  assign n172 = x7 ^ x2 ;
  assign n173 = n172 ^ n161 ;
  assign n174 = n173 ^ x7 ;
  assign n175 = n174 ^ n165 ;
  assign n176 = n168 ^ n165 ;
  assign n177 = n176 ^ n166 ;
  assign n178 = ~n175 & n177 ;
  assign n179 = n178 ^ n163 ;
  assign n180 = n179 ^ n165 ;
  assign n181 = n180 ^ n166 ;
  assign n182 = ~n171 & n181 ;
  assign n183 = n182 ^ n178 ;
  assign n184 = n183 ^ n163 ;
  assign n185 = n184 ^ n165 ;
  assign n186 = n185 ^ n166 ;
  assign n187 = n157 & n186 ;
  assign n188 = ~x0 & ~x7 ;
  assign n189 = x3 & n55 ;
  assign n190 = ~x3 & x8 ;
  assign n191 = ~n189 & ~n190 ;
  assign n192 = n188 & ~n191 ;
  assign n193 = x0 & ~x3 ;
  assign n194 = n12 & n193 ;
  assign n195 = ~n192 & ~n194 ;
  assign n196 = n115 & ~n195 ;
  assign n197 = ~n187 & ~n196 ;
  assign n198 = ~x4 & n21 ;
  assign n199 = ~n68 & ~n198 ;
  assign n200 = n193 & ~n199 ;
  assign n201 = n12 ^ x4 ;
  assign n202 = x0 & x3 ;
  assign n203 = n202 ^ n12 ;
  assign n204 = n203 ^ n202 ;
  assign n205 = n72 & n188 ;
  assign n206 = n205 ^ n202 ;
  assign n207 = ~n204 & ~n206 ;
  assign n208 = n207 ^ n202 ;
  assign n209 = ~n201 & n208 ;
  assign n210 = n209 ^ x4 ;
  assign n211 = ~n137 & ~n210 ;
  assign n212 = ~n200 & ~n211 ;
  assign n213 = n212 ^ x2 ;
  assign n214 = n213 ^ n212 ;
  assign n215 = n214 ^ x5 ;
  assign n216 = ~x4 & x8 ;
  assign n217 = x0 & n216 ;
  assign n218 = n152 ^ x7 ;
  assign n219 = ~x3 & n218 ;
  assign n220 = n219 ^ x7 ;
  assign n221 = n217 & n220 ;
  assign n222 = ~x3 & x4 ;
  assign n223 = x0 & n67 ;
  assign n224 = ~n93 & ~n223 ;
  assign n225 = n222 & ~n224 ;
  assign n226 = ~x9 & n225 ;
  assign n227 = ~n221 & ~n226 ;
  assign n228 = ~x0 & ~x9 ;
  assign n229 = n67 & n137 ;
  assign n230 = x4 & n190 ;
  assign n231 = ~n229 & ~n230 ;
  assign n232 = n228 & ~n231 ;
  assign n233 = n232 ^ n227 ;
  assign n234 = n227 & ~n233 ;
  assign n235 = n234 ^ n212 ;
  assign n236 = n235 ^ n227 ;
  assign n237 = ~n215 & n236 ;
  assign n238 = n237 ^ n234 ;
  assign n239 = n238 ^ n227 ;
  assign n240 = x5 & n239 ;
  assign n241 = n240 ^ x5 ;
  assign n242 = n197 & ~n241 ;
  assign n243 = ~n156 & n242 ;
  assign n244 = x6 & ~n243 ;
  assign n295 = x7 & n20 ;
  assign n296 = n22 & n295 ;
  assign n245 = ~x5 & ~x8 ;
  assign n297 = x0 & n245 ;
  assign n298 = n297 ^ n125 ;
  assign n299 = ~x6 & n14 ;
  assign n300 = n299 ^ n297 ;
  assign n301 = n300 ^ n299 ;
  assign n302 = x9 & n97 ;
  assign n303 = n302 ^ n299 ;
  assign n304 = n301 & ~n303 ;
  assign n305 = n304 ^ n299 ;
  assign n306 = n298 & ~n305 ;
  assign n307 = n306 ^ n125 ;
  assign n308 = ~n296 & ~n307 ;
  assign n309 = n222 & ~n308 ;
  assign n310 = ~x4 & ~x5 ;
  assign n277 = x3 & ~x9 ;
  assign n311 = n67 & n277 ;
  assign n312 = n310 & n311 ;
  assign n313 = ~x5 & x7 ;
  assign n314 = x8 & ~n313 ;
  assign n315 = n137 & ~n245 ;
  assign n316 = ~n314 & n315 ;
  assign n317 = n75 & n190 ;
  assign n318 = ~n316 & ~n317 ;
  assign n319 = x9 & ~n318 ;
  assign n320 = ~n312 & ~n319 ;
  assign n321 = x0 & ~x6 ;
  assign n322 = ~n320 & n321 ;
  assign n323 = ~n309 & ~n322 ;
  assign n324 = n149 & n202 ;
  assign n325 = n45 ^ n20 ;
  assign n326 = n20 ^ x5 ;
  assign n327 = n326 ^ n20 ;
  assign n328 = n327 ^ n324 ;
  assign n329 = n325 & ~n328 ;
  assign n330 = n329 ^ n45 ;
  assign n331 = n324 & n330 ;
  assign n332 = n323 & ~n331 ;
  assign n246 = n245 ^ x3 ;
  assign n247 = n246 ^ x4 ;
  assign n256 = n247 ^ n245 ;
  assign n248 = n245 ^ x4 ;
  assign n249 = n248 ^ n247 ;
  assign n250 = n249 ^ n247 ;
  assign n251 = n250 ^ n245 ;
  assign n252 = n249 ^ x0 ;
  assign n253 = n252 ^ n249 ;
  assign n254 = n253 ^ n251 ;
  assign n255 = ~n251 & ~n254 ;
  assign n257 = n256 ^ n255 ;
  assign n258 = n257 ^ n251 ;
  assign n259 = n245 ^ x5 ;
  assign n260 = n255 ^ n251 ;
  assign n261 = n259 & ~n260 ;
  assign n262 = n261 ^ n245 ;
  assign n263 = ~n258 & n262 ;
  assign n264 = n263 ^ n245 ;
  assign n265 = n264 ^ n245 ;
  assign n266 = n125 & n265 ;
  assign n267 = x8 ^ x5 ;
  assign n268 = x4 ^ x3 ;
  assign n269 = x8 ^ x4 ;
  assign n270 = n269 ^ x4 ;
  assign n271 = ~n268 & ~n270 ;
  assign n272 = n271 ^ x4 ;
  assign n273 = ~n267 & ~n272 ;
  assign n274 = x7 ^ x4 ;
  assign n275 = n31 & n274 ;
  assign n276 = n273 & n275 ;
  assign n278 = ~x0 & n277 ;
  assign n279 = n278 ^ x7 ;
  assign n280 = n96 ^ x4 ;
  assign n281 = n280 ^ n96 ;
  assign n282 = n96 ^ x5 ;
  assign n283 = n281 & n282 ;
  assign n284 = n283 ^ n96 ;
  assign n285 = n284 ^ n278 ;
  assign n286 = n279 & n285 ;
  assign n287 = n286 ^ n283 ;
  assign n288 = n287 ^ n96 ;
  assign n289 = n288 ^ x7 ;
  assign n290 = n278 & n289 ;
  assign n291 = n290 ^ n278 ;
  assign n292 = ~n276 & ~n291 ;
  assign n293 = ~n266 & n292 ;
  assign n294 = ~x6 & ~n293 ;
  assign n333 = n332 ^ n294 ;
  assign n334 = ~x2 & ~n333 ;
  assign n335 = n334 ^ n332 ;
  assign n336 = ~n244 & n335 ;
  assign n337 = n336 ^ x1 ;
  assign n338 = n337 ^ n336 ;
  assign n339 = n71 & n137 ;
  assign n340 = x9 ^ x3 ;
  assign n341 = x3 ^ x0 ;
  assign n342 = ~n340 & n341 ;
  assign n343 = n342 ^ x0 ;
  assign n344 = n93 & n343 ;
  assign n345 = ~x5 & ~n344 ;
  assign n346 = n55 & n188 ;
  assign n347 = ~x5 & ~x7 ;
  assign n348 = ~n311 & ~n347 ;
  assign n349 = ~n346 & n348 ;
  assign n350 = ~x6 & ~n349 ;
  assign n351 = ~n345 & n350 ;
  assign n352 = x8 & n75 ;
  assign n353 = n22 & n67 ;
  assign n354 = ~n352 & ~n353 ;
  assign n355 = x3 & n25 ;
  assign n356 = ~n354 & n355 ;
  assign n357 = ~n351 & ~n356 ;
  assign n358 = n115 & ~n357 ;
  assign n359 = ~n339 & ~n358 ;
  assign n360 = n321 & n352 ;
  assign n361 = n14 ^ x8 ;
  assign n362 = n361 ^ n14 ;
  assign n363 = n16 ^ n14 ;
  assign n364 = n362 & n363 ;
  assign n365 = n364 ^ n14 ;
  assign n366 = x7 & n365 ;
  assign n367 = n366 ^ n14 ;
  assign n368 = n367 ^ x7 ;
  assign n369 = n368 ^ x6 ;
  assign n376 = n369 ^ n368 ;
  assign n370 = n369 ^ n43 ;
  assign n371 = n370 ^ n368 ;
  assign n372 = n369 ^ n367 ;
  assign n373 = n372 ^ n43 ;
  assign n374 = n373 ^ n371 ;
  assign n375 = ~n371 & ~n374 ;
  assign n377 = n376 ^ n375 ;
  assign n378 = n377 ^ n371 ;
  assign n379 = n368 ^ n22 ;
  assign n380 = n375 ^ n371 ;
  assign n381 = ~n379 & ~n380 ;
  assign n382 = n381 ^ n368 ;
  assign n383 = ~n378 & n382 ;
  assign n384 = n383 ^ n368 ;
  assign n385 = n384 ^ x7 ;
  assign n386 = n385 ^ n368 ;
  assign n387 = ~n360 & ~n386 ;
  assign n388 = ~x9 & n137 ;
  assign n389 = ~n387 & n388 ;
  assign n390 = n53 ^ x6 ;
  assign n391 = n390 ^ n53 ;
  assign n392 = n53 ^ x4 ;
  assign n393 = n392 ^ n53 ;
  assign n394 = ~n391 & n393 ;
  assign n395 = n394 ^ n53 ;
  assign n396 = x8 & n395 ;
  assign n397 = n396 ^ n53 ;
  assign n398 = n32 & n397 ;
  assign n399 = n12 & n23 ;
  assign n400 = ~n398 & ~n399 ;
  assign n401 = x3 & ~n400 ;
  assign n402 = x0 & x5 ;
  assign n403 = ~x4 & n402 ;
  assign n404 = n97 & n403 ;
  assign n405 = n11 & n404 ;
  assign n406 = ~n401 & ~n405 ;
  assign n407 = ~n389 & n406 ;
  assign n408 = n407 ^ x2 ;
  assign n409 = n408 ^ n407 ;
  assign n410 = n409 ^ n359 ;
  assign n411 = x3 & ~x7 ;
  assign n412 = ~x4 & n55 ;
  assign n413 = ~n25 & ~n412 ;
  assign n414 = n402 & ~n413 ;
  assign n415 = ~n44 & n414 ;
  assign n416 = n11 & n310 ;
  assign n417 = x6 & n416 ;
  assign n418 = ~n415 & ~n417 ;
  assign n419 = n418 ^ n411 ;
  assign n420 = n411 & ~n419 ;
  assign n421 = n420 ^ n407 ;
  assign n422 = n421 ^ n411 ;
  assign n423 = ~n410 & ~n422 ;
  assign n424 = n423 ^ n420 ;
  assign n425 = n424 ^ n411 ;
  assign n426 = n359 & n425 ;
  assign n427 = n426 ^ n359 ;
  assign n428 = n427 ^ n336 ;
  assign n429 = ~n338 & n428 ;
  assign n430 = n429 ^ n336 ;
  assign n431 = n430 ^ n136 ;
  assign n432 = n145 & ~n431 ;
  assign n433 = n432 ^ n429 ;
  assign n434 = n433 ^ n336 ;
  assign n435 = n434 ^ n144 ;
  assign n436 = ~n136 & ~n435 ;
  assign n437 = n436 ^ n136 ;
  assign y0 = n437 ;
endmodule
