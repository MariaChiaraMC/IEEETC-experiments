module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n13 = ~x2 & x4 ;
  assign n14 = ~x0 & ~n13 ;
  assign n15 = x1 & ~x4 ;
  assign n16 = x2 & ~x3 ;
  assign n17 = ~n15 & n16 ;
  assign n18 = x6 & ~x7 ;
  assign n19 = ~x5 & ~x8 ;
  assign n20 = n18 & n19 ;
  assign n21 = x10 ^ x9 ;
  assign n22 = n21 ^ x11 ;
  assign n23 = x10 & x11 ;
  assign n24 = n22 & n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n20 & n25 ;
  assign n27 = ~n17 & n26 ;
  assign n28 = n14 & ~n27 ;
  assign y0 = ~n28 ;
endmodule
