module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 ;
  assign n8 = ~x0 & x1 ;
  assign n9 = ~x3 & n8 ;
  assign n10 = ~x4 & n9 ;
  assign n14 = ~x0 & x3 ;
  assign n18 = ~x4 & ~x5 ;
  assign n19 = ~n14 & ~n18 ;
  assign n20 = x1 ^ x0 ;
  assign n21 = n19 & ~n20 ;
  assign n22 = ~x2 & ~n21 ;
  assign n11 = x5 & x6 ;
  assign n12 = x1 & n11 ;
  assign n13 = x1 & x4 ;
  assign n15 = ~n13 & n14 ;
  assign n16 = ~n12 & n15 ;
  assign n17 = x2 & ~n16 ;
  assign n23 = n22 ^ n17 ;
  assign n24 = n17 ^ x3 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = ~x5 & ~x6 ;
  assign n33 = x4 & ~n26 ;
  assign n34 = ~x1 & ~n33 ;
  assign n35 = n11 & n13 ;
  assign n36 = ~x0 & ~n35 ;
  assign n37 = ~n34 & n36 ;
  assign n27 = n26 ^ x4 ;
  assign n28 = x4 ^ x1 ;
  assign n29 = n27 & n28 ;
  assign n30 = n29 ^ x1 ;
  assign n31 = x0 & ~n30 ;
  assign n32 = ~n8 & ~n31 ;
  assign n38 = n37 ^ n32 ;
  assign n39 = x3 & n38 ;
  assign n40 = n39 ^ n32 ;
  assign n41 = n25 & n40 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = n42 ^ n32 ;
  assign n44 = n43 ^ x3 ;
  assign n45 = n23 & n44 ;
  assign n46 = n45 ^ n22 ;
  assign n47 = ~n10 & n46 ;
  assign y0 = ~n47 ;
endmodule
