module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;
  assign n29 = ~x0 & x2 ;
  assign n7 = ~x3 & x5 ;
  assign n8 = n7 ^ x0 ;
  assign n9 = x3 ^ x1 ;
  assign n10 = n9 ^ x3 ;
  assign n11 = x5 ^ x3 ;
  assign n12 = ~n10 & ~n11 ;
  assign n13 = n12 ^ x3 ;
  assign n14 = ~x2 & ~n13 ;
  assign n15 = n14 ^ n7 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n16 ^ n8 ;
  assign n18 = x2 ^ x1 ;
  assign n19 = x2 & n18 ;
  assign n20 = n19 ^ n14 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = n17 & n21 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n23 ^ x2 ;
  assign n25 = n8 & n24 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = n30 ^ n25 ;
  assign n26 = ~x1 & ~x5 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = n27 ^ n25 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = n25 ^ x3 ;
  assign n34 = n33 ^ n25 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = n31 & ~n35 ;
  assign n37 = n36 ^ n31 ;
  assign n38 = n32 & n37 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n39 ^ n25 ;
  assign n41 = n40 ^ n31 ;
  assign n42 = ~x4 & n41 ;
  assign n43 = n42 ^ n25 ;
  assign y0 = n43 ;
endmodule
