module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n20 = ~x12 & x15 ;
  assign n21 = ~x5 & n20 ;
  assign n22 = ~x2 & x7 ;
  assign n23 = ~x3 & ~n22 ;
  assign n24 = n21 & n23 ;
  assign n25 = x13 & x17 ;
  assign n26 = x9 & x11 ;
  assign n27 = ~x6 & n26 ;
  assign n28 = n25 & n27 ;
  assign n29 = n24 & n28 ;
  assign n30 = ~x4 & x18 ;
  assign n31 = ~x1 & x8 ;
  assign n32 = ~x10 & x16 ;
  assign n33 = x0 & x14 ;
  assign n34 = n32 & n33 ;
  assign n35 = n31 & n34 ;
  assign n36 = n30 & n35 ;
  assign n37 = n29 & n36 ;
  assign y0 = n37 ;
endmodule
