module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n11 = ~x6 & ~x7 ;
  assign n12 = ~x5 & n11 ;
  assign n13 = ~x0 & ~x1 ;
  assign n14 = ~x2 & ~x3 ;
  assign n15 = n13 & n14 ;
  assign n16 = n15 ^ x4 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = x2 & x3 ;
  assign n20 = x9 ^ x1 ;
  assign n19 = x8 ^ x1 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = x1 ^ x0 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = ~n20 & ~n23 ;
  assign n25 = n24 ^ n20 ;
  assign n26 = n21 & ~n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n27 ^ x1 ;
  assign n29 = n28 ^ n20 ;
  assign n30 = n18 & ~n29 ;
  assign n31 = n30 ^ n15 ;
  assign n32 = ~n17 & n31 ;
  assign n33 = n32 ^ n15 ;
  assign n34 = n12 & n33 ;
  assign y0 = n34 ;
endmodule
