module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 ;
  assign n8 = ~x0 & ~x1 ;
  assign n9 = x3 & ~x6 ;
  assign n10 = n9 ^ x2 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = ~x5 & x6 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = n13 ^ n9 ;
  assign n15 = n11 & n14 ;
  assign n16 = n15 ^ n9 ;
  assign n17 = x4 & n16 ;
  assign n18 = n17 ^ n9 ;
  assign n19 = ~n8 & n18 ;
  assign n20 = ~x4 & ~x6 ;
  assign n21 = x2 & x3 ;
  assign n22 = x5 & ~n21 ;
  assign n23 = n20 & ~n22 ;
  assign n24 = ~n19 & ~n23 ;
  assign n26 = x1 & n21 ;
  assign n27 = x5 & ~n26 ;
  assign n25 = x6 ^ x4 ;
  assign n28 = n27 ^ n25 ;
  assign n37 = n28 ^ n27 ;
  assign n29 = n28 ^ x6 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = ~x2 & ~x3 ;
  assign n32 = ~n12 & ~n31 ;
  assign n33 = n32 ^ x6 ;
  assign n34 = n33 ^ x6 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n30 & ~n35 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = n38 ^ n30 ;
  assign n40 = n27 ^ x3 ;
  assign n41 = n36 ^ n30 ;
  assign n42 = ~n40 & n41 ;
  assign n43 = n42 ^ n27 ;
  assign n44 = n39 & ~n43 ;
  assign n45 = n44 ^ n27 ;
  assign n46 = n45 ^ n25 ;
  assign n47 = n46 ^ n27 ;
  assign n48 = n24 & ~n47 ;
  assign y0 = ~n48 ;
endmodule
