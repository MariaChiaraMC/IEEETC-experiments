module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 ;
  assign n9 = x1 & x5 ;
  assign n10 = ~x3 & ~x7 ;
  assign n11 = n9 & ~n10 ;
  assign n12 = x6 & n11 ;
  assign n13 = x4 & ~n12 ;
  assign n14 = x6 ^ x5 ;
  assign n15 = n14 ^ x2 ;
  assign n16 = x1 & x3 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = x6 ^ x2 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = x7 ^ x2 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = n19 & ~n21 ;
  assign n23 = n22 ^ x2 ;
  assign n24 = n23 ^ n15 ;
  assign n25 = ~n17 & ~n24 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = n26 ^ x2 ;
  assign n28 = n27 ^ n16 ;
  assign n29 = ~n15 & n28 ;
  assign n30 = n29 ^ n15 ;
  assign n31 = ~n13 & n30 ;
  assign n32 = ~x0 & ~n31 ;
  assign n33 = x2 & x6 ;
  assign n34 = x3 & x7 ;
  assign n35 = n33 & n34 ;
  assign n36 = ~x1 & ~n35 ;
  assign n37 = ~x7 & ~n33 ;
  assign n38 = n37 ^ x5 ;
  assign n39 = x6 ^ x0 ;
  assign n40 = n39 ^ x0 ;
  assign n41 = x2 & ~x3 ;
  assign n42 = n41 ^ x0 ;
  assign n43 = ~n40 & ~n42 ;
  assign n44 = n43 ^ x0 ;
  assign n45 = n44 ^ n37 ;
  assign n46 = ~n38 & n45 ;
  assign n47 = n46 ^ n43 ;
  assign n48 = n47 ^ x0 ;
  assign n49 = n48 ^ x5 ;
  assign n50 = ~n37 & ~n49 ;
  assign n51 = n50 ^ n37 ;
  assign n52 = ~n36 & ~n51 ;
  assign n53 = x2 & n11 ;
  assign n54 = x0 & ~n53 ;
  assign n55 = ~x4 & ~n54 ;
  assign n56 = ~n52 & n55 ;
  assign n58 = ~x1 & ~x5 ;
  assign n57 = ~n9 & ~n34 ;
  assign n59 = n58 ^ n57 ;
  assign n60 = n59 ^ x4 ;
  assign n61 = ~x2 & ~x6 ;
  assign n62 = n61 ^ n33 ;
  assign n63 = ~n58 & n62 ;
  assign n64 = n63 ^ n33 ;
  assign n65 = n60 & n64 ;
  assign n66 = n65 ^ n63 ;
  assign n67 = n66 ^ n33 ;
  assign n68 = n67 ^ n58 ;
  assign n69 = x4 & ~n68 ;
  assign n70 = ~n56 & ~n69 ;
  assign n71 = ~n32 & ~n70 ;
  assign y0 = ~n71 ;
endmodule
