// Benchmark "./dk48.pla" written by ABC on Thu Apr 23 10:59:50 2020

module \./dk48.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    z3  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14;
  output z3;
  assign z3 = 1'b1;
endmodule


