module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 ;
  assign n9 = x0 & ~x7 ;
  assign n10 = x6 ^ x4 ;
  assign n11 = x1 & ~n10 ;
  assign n12 = n11 ^ x2 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = ~x1 & ~x4 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = n13 & n15 ;
  assign n17 = n16 ^ n11 ;
  assign n18 = n9 & n17 ;
  assign n19 = n18 ^ x5 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = x1 & x4 ;
  assign n22 = x2 & n21 ;
  assign n23 = x0 & x6 ;
  assign n24 = n23 ^ x6 ;
  assign n25 = x7 & ~n24 ;
  assign n26 = n25 ^ x6 ;
  assign n27 = n22 & ~n26 ;
  assign n28 = x4 ^ x1 ;
  assign n29 = n23 & n28 ;
  assign n30 = n29 ^ x7 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = ~x6 & n14 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n31 & n33 ;
  assign n35 = n34 ^ n29 ;
  assign n36 = ~x2 & n35 ;
  assign n37 = ~n27 & ~n36 ;
  assign n38 = n37 ^ n18 ;
  assign n39 = n20 & ~n38 ;
  assign n40 = n39 ^ n18 ;
  assign n41 = x3 & n40 ;
  assign n68 = x3 & ~x4 ;
  assign n69 = x1 & ~x5 ;
  assign n70 = n10 & n69 ;
  assign n71 = x2 & ~n70 ;
  assign n72 = ~n68 & ~n71 ;
  assign n44 = ~x1 & ~x3 ;
  assign n73 = ~x4 & x5 ;
  assign n74 = n44 & n73 ;
  assign n75 = x6 & n74 ;
  assign n76 = ~n72 & ~n75 ;
  assign n46 = x1 & x3 ;
  assign n56 = ~x4 & ~x7 ;
  assign n57 = n46 & n56 ;
  assign n43 = x4 & ~x6 ;
  assign n45 = n44 ^ n43 ;
  assign n47 = x7 & ~n46 ;
  assign n48 = n47 ^ n43 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = ~x6 & ~x7 ;
  assign n51 = ~x4 & ~n50 ;
  assign n52 = n51 ^ n47 ;
  assign n53 = ~n49 & n52 ;
  assign n54 = n53 ^ n47 ;
  assign n55 = n45 & ~n54 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = n58 ^ n55 ;
  assign n60 = n55 ^ x6 ;
  assign n61 = n60 ^ n55 ;
  assign n62 = n59 & n61 ;
  assign n63 = n62 ^ n55 ;
  assign n64 = ~x5 & n63 ;
  assign n65 = n64 ^ n55 ;
  assign n66 = n65 ^ x2 ;
  assign n42 = x7 ^ x2 ;
  assign n67 = n66 ^ n42 ;
  assign n77 = n76 ^ n67 ;
  assign n78 = n77 ^ n67 ;
  assign n79 = n67 ^ n66 ;
  assign n80 = n79 ^ x2 ;
  assign n81 = ~n78 & n80 ;
  assign n82 = n81 ^ n66 ;
  assign n83 = x5 & ~x6 ;
  assign n84 = ~x5 & x6 ;
  assign n85 = x4 & ~n84 ;
  assign n86 = ~n83 & n85 ;
  assign n87 = x3 ^ x1 ;
  assign n88 = x5 ^ x3 ;
  assign n89 = n87 & n88 ;
  assign n90 = n89 ^ x1 ;
  assign n91 = n86 & ~n90 ;
  assign n92 = ~n66 & n91 ;
  assign n93 = n92 ^ x2 ;
  assign n94 = ~n82 & ~n93 ;
  assign n95 = n94 ^ n92 ;
  assign n96 = ~x2 & n95 ;
  assign n97 = n96 ^ n81 ;
  assign n98 = n97 ^ n65 ;
  assign n99 = n98 ^ n66 ;
  assign n100 = n99 ^ x0 ;
  assign n101 = n100 ^ n99 ;
  assign n102 = ~x2 & n84 ;
  assign n103 = ~n83 & ~n102 ;
  assign n104 = x7 & n44 ;
  assign n105 = x4 & n104 ;
  assign n106 = ~n103 & n105 ;
  assign n107 = x2 & ~x3 ;
  assign n108 = x5 ^ x4 ;
  assign n109 = n108 ^ x1 ;
  assign n116 = n109 ^ x5 ;
  assign n111 = n109 ^ x6 ;
  assign n117 = n116 ^ n111 ;
  assign n118 = n117 ^ n111 ;
  assign n110 = n109 ^ x7 ;
  assign n112 = n111 ^ n110 ;
  assign n113 = n112 ^ n109 ;
  assign n114 = n113 ^ n108 ;
  assign n115 = n114 ^ n111 ;
  assign n119 = n118 ^ n115 ;
  assign n122 = n114 ^ n108 ;
  assign n120 = n109 ^ n108 ;
  assign n121 = n120 ^ n115 ;
  assign n123 = n122 ^ n121 ;
  assign n124 = n119 & ~n123 ;
  assign n125 = n124 ^ n114 ;
  assign n126 = n125 ^ n120 ;
  assign n127 = n126 ^ n122 ;
  assign n128 = n121 ^ n118 ;
  assign n129 = n125 & ~n128 ;
  assign n130 = n129 ^ n114 ;
  assign n131 = n130 ^ n115 ;
  assign n132 = n131 ^ n118 ;
  assign n133 = ~n127 & n132 ;
  assign n134 = n107 & n133 ;
  assign n135 = ~n106 & ~n134 ;
  assign n136 = n135 ^ n99 ;
  assign n137 = n101 & n136 ;
  assign n138 = n137 ^ n99 ;
  assign n139 = ~n41 & n138 ;
  assign y0 = ~n139 ;
endmodule
