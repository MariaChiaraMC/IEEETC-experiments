module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 ;
  output y0 ;
  wire n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 ;
  assign n28 = x24 & x25 ;
  assign n29 = x19 & x21 ;
  assign n30 = x3 & x26 ;
  assign n31 = x4 & x22 ;
  assign n32 = n30 & n31 ;
  assign n33 = x18 & x23 ;
  assign n34 = n32 & n33 ;
  assign n35 = n29 & n34 ;
  assign n36 = x0 & x17 ;
  assign n37 = x20 & n36 ;
  assign n38 = x2 & x5 ;
  assign n39 = n37 & n38 ;
  assign n40 = x1 & n39 ;
  assign n41 = n35 & n40 ;
  assign n42 = x6 & n41 ;
  assign n43 = ~x17 & ~x19 ;
  assign n44 = ~x18 & n43 ;
  assign n45 = ~x2 & ~x26 ;
  assign n46 = ~x1 & n45 ;
  assign n47 = n44 & n46 ;
  assign n48 = ~x0 & ~x20 ;
  assign n49 = ~x3 & ~x22 ;
  assign n50 = n48 & n49 ;
  assign n51 = ~x5 & ~x21 ;
  assign n52 = ~x4 & ~x23 ;
  assign n53 = n51 & n52 ;
  assign n54 = n50 & n53 ;
  assign n55 = n47 & n54 ;
  assign n56 = x14 & n55 ;
  assign n57 = ~n42 & ~n56 ;
  assign n58 = x9 ^ x8 ;
  assign n59 = x9 & ~n58 ;
  assign n60 = x7 & n59 ;
  assign n61 = n60 ^ n58 ;
  assign n62 = ~n57 & ~n61 ;
  assign n63 = x15 & n55 ;
  assign n64 = x10 & n41 ;
  assign n65 = ~n63 & ~n64 ;
  assign n66 = ~x11 & ~x12 ;
  assign n67 = ~n65 & n66 ;
  assign n68 = n67 ^ x7 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = n69 ^ n62 ;
  assign n71 = ~x8 & ~x9 ;
  assign n72 = x16 & n55 ;
  assign n73 = x13 & n41 ;
  assign n74 = ~n72 & ~n73 ;
  assign n75 = n74 ^ n71 ;
  assign n76 = ~n71 & n75 ;
  assign n77 = n76 ^ n67 ;
  assign n78 = n77 ^ n71 ;
  assign n79 = ~n70 & ~n78 ;
  assign n80 = n79 ^ n76 ;
  assign n81 = n80 ^ n71 ;
  assign n82 = ~n62 & ~n81 ;
  assign n83 = n82 ^ n62 ;
  assign n84 = ~n28 & n83 ;
  assign y0 = n84 ;
endmodule
