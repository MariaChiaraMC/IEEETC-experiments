module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 ;
  assign n11 = ~x1 & ~x2 ;
  assign n29 = ~x6 & ~x9 ;
  assign n30 = ~x0 & ~x3 ;
  assign n31 = ~x5 & n30 ;
  assign n32 = ~n29 & n31 ;
  assign n12 = ~x5 & ~x6 ;
  assign n13 = ~x9 & ~n12 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = n14 ^ n13 ;
  assign n17 = x6 ^ x0 ;
  assign n18 = n17 ^ n13 ;
  assign n16 = x6 ^ x3 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n19 ^ n15 ;
  assign n21 = n15 & ~n20 ;
  assign n22 = n21 ^ n14 ;
  assign n23 = n22 ^ n15 ;
  assign n24 = x3 & n18 ;
  assign n25 = n24 ^ n14 ;
  assign n26 = ~n23 & ~n25 ;
  assign n27 = n26 ^ n14 ;
  assign n28 = n27 ^ n13 ;
  assign n33 = n32 ^ n28 ;
  assign n34 = ~x4 & ~n33 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = ~x8 & n35 ;
  assign n37 = ~x4 & x9 ;
  assign n38 = ~x5 & ~n37 ;
  assign n39 = x8 ^ x6 ;
  assign n40 = ~n38 & ~n39 ;
  assign n42 = ~x3 & ~x4 ;
  assign n41 = x0 & ~x9 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = n43 ^ n41 ;
  assign n45 = n41 ^ x0 ;
  assign n46 = ~n44 & ~n45 ;
  assign n47 = n46 ^ n41 ;
  assign n48 = x3 & x5 ;
  assign n49 = ~n41 & n48 ;
  assign n50 = n49 ^ n40 ;
  assign n51 = ~n47 & n50 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = n40 & n52 ;
  assign n54 = n53 ^ n40 ;
  assign n55 = ~n36 & ~n54 ;
  assign n56 = n11 & ~n55 ;
  assign n57 = ~x0 & x3 ;
  assign n58 = x2 & ~x3 ;
  assign n59 = ~n57 & ~n58 ;
  assign n60 = x5 & x6 ;
  assign n61 = n60 ^ x8 ;
  assign n62 = ~n30 & ~n60 ;
  assign n63 = ~n61 & n62 ;
  assign n64 = n63 ^ n61 ;
  assign n65 = ~n59 & ~n64 ;
  assign n67 = ~x6 & ~x8 ;
  assign n66 = x6 & x8 ;
  assign n68 = n67 ^ n66 ;
  assign n69 = x0 & n68 ;
  assign n70 = n69 ^ n67 ;
  assign n71 = n48 & n70 ;
  assign n72 = x0 & ~x8 ;
  assign n73 = ~n60 & n72 ;
  assign n74 = n73 ^ x5 ;
  assign n75 = n74 ^ x2 ;
  assign n98 = ~x3 & ~x9 ;
  assign n76 = ~n41 & ~n67 ;
  assign n77 = n76 ^ x9 ;
  assign n78 = n77 ^ x3 ;
  assign n86 = n78 ^ n77 ;
  assign n79 = x3 & ~x8 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n78 ^ n76 ;
  assign n83 = n82 ^ n79 ;
  assign n84 = n83 ^ n81 ;
  assign n85 = ~n81 & ~n84 ;
  assign n87 = n86 ^ n85 ;
  assign n88 = n87 ^ n81 ;
  assign n89 = ~x0 & x8 ;
  assign n90 = n89 ^ n77 ;
  assign n91 = n85 ^ n81 ;
  assign n92 = n90 & ~n91 ;
  assign n93 = n92 ^ n77 ;
  assign n94 = ~n88 & ~n93 ;
  assign n95 = n94 ^ n77 ;
  assign n96 = n95 ^ x9 ;
  assign n97 = n96 ^ n77 ;
  assign n99 = n98 ^ n97 ;
  assign n100 = ~x5 & n99 ;
  assign n101 = n100 ^ n98 ;
  assign n102 = ~n75 & ~n101 ;
  assign n103 = n102 ^ n100 ;
  assign n104 = n103 ^ n98 ;
  assign n105 = n104 ^ x5 ;
  assign n106 = x2 & n105 ;
  assign n107 = ~n71 & ~n106 ;
  assign n108 = n107 ^ x1 ;
  assign n109 = n108 ^ n107 ;
  assign n110 = ~x0 & ~x8 ;
  assign n111 = ~x2 & n110 ;
  assign n112 = x0 & x8 ;
  assign n113 = n112 ^ x9 ;
  assign n114 = n113 ^ x2 ;
  assign n115 = n114 ^ n113 ;
  assign n116 = n115 ^ x3 ;
  assign n117 = x9 & ~n72 ;
  assign n118 = n113 ^ n112 ;
  assign n119 = n118 ^ n117 ;
  assign n120 = ~n117 & ~n119 ;
  assign n121 = n120 ^ n113 ;
  assign n122 = n121 ^ n117 ;
  assign n123 = ~n116 & n122 ;
  assign n124 = n123 ^ n120 ;
  assign n125 = n124 ^ n117 ;
  assign n126 = x3 & ~n125 ;
  assign n127 = ~n111 & ~n126 ;
  assign n128 = ~x6 & ~n127 ;
  assign n129 = x0 & n66 ;
  assign n130 = ~n58 & n129 ;
  assign n131 = x5 & ~n130 ;
  assign n132 = ~n128 & n131 ;
  assign n133 = n132 ^ x3 ;
  assign n134 = ~x5 & ~n79 ;
  assign n135 = n134 ^ n133 ;
  assign n136 = n135 ^ n132 ;
  assign n137 = n136 ^ n135 ;
  assign n138 = x0 & ~x6 ;
  assign n139 = n138 ^ x2 ;
  assign n140 = n139 ^ x8 ;
  assign n141 = n140 ^ n138 ;
  assign n142 = n141 ^ n140 ;
  assign n143 = n13 & n89 ;
  assign n144 = n143 ^ n140 ;
  assign n145 = n144 ^ n139 ;
  assign n146 = n142 & n145 ;
  assign n147 = n146 ^ n143 ;
  assign n148 = ~x9 & ~n143 ;
  assign n149 = n148 ^ n139 ;
  assign n150 = ~n147 & n149 ;
  assign n151 = n150 ^ n148 ;
  assign n152 = n139 & n151 ;
  assign n153 = n152 ^ n146 ;
  assign n154 = n153 ^ x2 ;
  assign n155 = n154 ^ n143 ;
  assign n156 = n155 ^ n135 ;
  assign n157 = n156 ^ n133 ;
  assign n158 = ~n137 & n157 ;
  assign n159 = n158 ^ n155 ;
  assign n160 = x2 ^ x0 ;
  assign n161 = n160 ^ x8 ;
  assign n162 = x8 ^ x2 ;
  assign n163 = n162 ^ x8 ;
  assign n164 = n163 ^ n161 ;
  assign n165 = x9 ^ x6 ;
  assign n166 = x6 & n165 ;
  assign n167 = n166 ^ x8 ;
  assign n168 = n167 ^ x6 ;
  assign n169 = ~n164 & ~n168 ;
  assign n170 = n169 ^ n166 ;
  assign n171 = n170 ^ x6 ;
  assign n172 = ~n161 & n171 ;
  assign n173 = ~n155 & ~n172 ;
  assign n174 = n173 ^ n133 ;
  assign n175 = ~n159 & ~n174 ;
  assign n176 = n175 ^ n173 ;
  assign n177 = ~n133 & n176 ;
  assign n178 = n177 ^ n158 ;
  assign n179 = n178 ^ x3 ;
  assign n180 = n179 ^ n155 ;
  assign n181 = n180 ^ n107 ;
  assign n182 = n109 & ~n181 ;
  assign n183 = n182 ^ n107 ;
  assign n184 = ~n65 & n183 ;
  assign n185 = ~x4 & ~n184 ;
  assign n186 = ~n56 & ~n185 ;
  assign n187 = ~x7 & ~n186 ;
  assign n188 = ~x9 & n11 ;
  assign n189 = ~n89 & n188 ;
  assign n190 = x2 ^ x1 ;
  assign n191 = x7 & n190 ;
  assign n193 = ~n89 & n117 ;
  assign n194 = ~n41 & ~n193 ;
  assign n192 = ~x9 & n89 ;
  assign n195 = n194 ^ n192 ;
  assign n196 = n194 ^ x1 ;
  assign n197 = n196 ^ n194 ;
  assign n198 = n197 ^ n191 ;
  assign n199 = ~n195 & ~n198 ;
  assign n200 = n199 ^ n192 ;
  assign n201 = n191 & n200 ;
  assign n202 = ~n189 & ~n201 ;
  assign n203 = n12 & n42 ;
  assign n204 = ~n202 & n203 ;
  assign n205 = ~n187 & ~n204 ;
  assign y0 = ~n205 ;
endmodule
