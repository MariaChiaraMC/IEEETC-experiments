module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 ;
  assign n9 = x5 ^ x4 ;
  assign n10 = ~x1 & n9 ;
  assign n11 = n10 ^ x4 ;
  assign n15 = n11 ^ x6 ;
  assign n14 = n11 ^ x7 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n15 ^ x1 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n16 & n18 ;
  assign n20 = n19 ^ n15 ;
  assign n21 = x0 & ~n20 ;
  assign n12 = x2 & ~x3 ;
  assign n13 = n12 ^ n11 ;
  assign n22 = n21 ^ n13 ;
  assign y0 = ~n22 ;
endmodule
