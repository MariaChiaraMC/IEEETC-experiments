module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n15 = x11 ^ x9 ;
  assign n20 = n15 ^ x9 ;
  assign n17 = x13 ^ x9 ;
  assign n16 = n15 ^ x12 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = n18 ^ x9 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = n16 ^ n15 ;
  assign n23 = n22 ^ x9 ;
  assign n24 = n23 ^ x9 ;
  assign n25 = n18 & ~n24 ;
  assign n26 = n25 ^ n18 ;
  assign n27 = ~n23 & n26 ;
  assign n28 = n27 ^ x9 ;
  assign n29 = n21 & n28 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = n30 ^ x9 ;
  assign n32 = n31 ^ n20 ;
  assign y0 = n32 ;
endmodule
