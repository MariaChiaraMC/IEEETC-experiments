module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 ;
  assign n15 = x7 ^ x5 ;
  assign n16 = n15 ^ x5 ;
  assign n17 = x5 ^ x1 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = n16 & n18 ;
  assign n20 = n19 ^ x5 ;
  assign n21 = ~x2 & n20 ;
  assign n22 = n21 ^ x5 ;
  assign n23 = x0 & n22 ;
  assign n24 = ~x3 & ~x4 ;
  assign n25 = ~x2 & x6 ;
  assign n26 = n24 & n25 ;
  assign n27 = x2 & x5 ;
  assign n28 = n27 ^ x1 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = ~x0 & x7 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = ~n29 & n31 ;
  assign n33 = n32 ^ n27 ;
  assign n34 = ~n26 & ~n33 ;
  assign n35 = ~n23 & n34 ;
  assign n36 = ~x10 & ~x13 ;
  assign n37 = ~x8 & ~x11 ;
  assign n38 = ~x12 & n37 ;
  assign n39 = ~x9 & n38 ;
  assign n40 = n36 & n39 ;
  assign n41 = ~n35 & n40 ;
  assign y0 = n41 ;
endmodule
