module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 ;
  assign n22 = x19 & x20 ;
  assign n23 = ~x4 & n22 ;
  assign n24 = n23 ^ x18 ;
  assign n25 = ~x0 & n24 ;
  assign y0 = n25 ;
endmodule
