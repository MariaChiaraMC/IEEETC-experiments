module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 ;
  assign n20 = ~x14 & x15 ;
  assign n21 = x17 ^ x16 ;
  assign n22 = n21 ^ x8 ;
  assign n23 = n22 ^ x7 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n24 ^ x17 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = x6 & n26 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = x7 ^ x6 ;
  assign n30 = n29 ^ n21 ;
  assign n31 = ~n25 & ~n30 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = n32 ^ n25 ;
  assign n34 = n28 & n33 ;
  assign n35 = ~n24 & n34 ;
  assign n36 = n35 ^ n27 ;
  assign n37 = n36 ^ x16 ;
  assign n38 = n20 & n37 ;
  assign n39 = ~x16 & ~x17 ;
  assign n40 = x14 & ~x15 ;
  assign n41 = ~x8 & n40 ;
  assign n42 = ~x10 & x15 ;
  assign n43 = ~x2 & n42 ;
  assign n44 = ~x3 & ~x15 ;
  assign n45 = ~x14 & ~n44 ;
  assign n46 = ~n43 & n45 ;
  assign n47 = ~x8 & n20 ;
  assign n48 = x9 & n47 ;
  assign n49 = ~n46 & ~n48 ;
  assign n50 = ~n41 & n49 ;
  assign n51 = ~n39 & ~n50 ;
  assign n55 = ~x11 & ~x12 ;
  assign n56 = x1 & ~x13 ;
  assign n57 = ~n55 & n56 ;
  assign n52 = ~x7 & x16 ;
  assign n53 = x6 & x16 ;
  assign n54 = ~n52 & ~n53 ;
  assign n58 = n57 ^ n54 ;
  assign n59 = n58 ^ x14 ;
  assign n60 = n59 ^ n58 ;
  assign n62 = x7 & x8 ;
  assign n61 = ~x8 & ~x9 ;
  assign n63 = n62 ^ n61 ;
  assign n64 = n63 ^ n62 ;
  assign n65 = n62 ^ x7 ;
  assign n66 = n65 ^ n62 ;
  assign n67 = n64 & ~n66 ;
  assign n68 = n67 ^ n62 ;
  assign n69 = x6 & n68 ;
  assign n70 = n69 ^ n62 ;
  assign n71 = x4 & n70 ;
  assign n72 = n71 ^ n58 ;
  assign n73 = n72 ^ n54 ;
  assign n74 = n60 ^ x16 ;
  assign n75 = n74 ^ n60 ;
  assign n76 = n73 & n75 ;
  assign n77 = n76 ^ n58 ;
  assign n78 = n58 ^ n54 ;
  assign n79 = n74 & n78 ;
  assign n80 = n79 ^ n60 ;
  assign n81 = n80 ^ n74 ;
  assign n82 = ~n77 & n81 ;
  assign n83 = n60 & n82 ;
  assign n84 = n83 ^ n76 ;
  assign n85 = n84 ^ n57 ;
  assign n86 = n85 ^ x17 ;
  assign n87 = n86 ^ n85 ;
  assign n88 = n87 ^ x15 ;
  assign n89 = ~x7 & ~x14 ;
  assign n90 = ~n61 & ~n89 ;
  assign n91 = ~x7 & ~x8 ;
  assign n92 = x4 & ~n91 ;
  assign n93 = x16 ^ x6 ;
  assign n94 = n92 & ~n93 ;
  assign n95 = ~n90 & n94 ;
  assign n96 = ~x7 & ~n93 ;
  assign n97 = x14 & ~n96 ;
  assign n98 = n97 ^ n95 ;
  assign n99 = ~n95 & n98 ;
  assign n100 = n99 ^ n85 ;
  assign n101 = n100 ^ n95 ;
  assign n102 = ~n88 & n101 ;
  assign n103 = n102 ^ n99 ;
  assign n104 = n103 ^ n95 ;
  assign n105 = ~x15 & ~n104 ;
  assign n106 = n105 ^ x15 ;
  assign n107 = ~n51 & n106 ;
  assign n108 = ~n38 & n107 ;
  assign n109 = n108 ^ x18 ;
  assign n110 = n109 ^ n108 ;
  assign n112 = n40 ^ x8 ;
  assign n120 = n112 ^ n40 ;
  assign n111 = n40 ^ x14 ;
  assign n113 = n112 ^ n111 ;
  assign n114 = n113 ^ n112 ;
  assign n115 = n114 ^ n40 ;
  assign n116 = n113 ^ n43 ;
  assign n117 = n116 ^ n113 ;
  assign n118 = n117 ^ n115 ;
  assign n119 = ~n115 & ~n118 ;
  assign n121 = n120 ^ n119 ;
  assign n122 = n121 ^ n115 ;
  assign n123 = n40 ^ x9 ;
  assign n124 = n119 ^ n115 ;
  assign n125 = n123 & ~n124 ;
  assign n126 = n125 ^ n40 ;
  assign n127 = n122 & ~n126 ;
  assign n128 = n127 ^ n40 ;
  assign n129 = n128 ^ x8 ;
  assign n130 = n129 ^ n40 ;
  assign n131 = x7 & ~x17 ;
  assign n132 = ~x7 & x17 ;
  assign n133 = ~n131 & ~n132 ;
  assign n134 = ~n93 & n133 ;
  assign n135 = ~n130 & n134 ;
  assign n136 = n135 ^ n108 ;
  assign n137 = n110 & ~n136 ;
  assign n138 = n137 ^ n108 ;
  assign n139 = ~x0 & ~n138 ;
  assign y0 = n139 ;
endmodule
