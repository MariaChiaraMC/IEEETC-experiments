module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 ;
  assign n33 = ~x2 & ~x3 ;
  assign n34 = ~x6 & ~x7 ;
  assign n35 = ~x10 & ~x11 ;
  assign n36 = ~x14 & ~x15 ;
  assign n37 = ~x18 & ~x19 ;
  assign n38 = ~x22 & ~x23 ;
  assign n39 = ~x26 & ~x27 ;
  assign n40 = ~x30 & ~x31 ;
  assign n41 = ~x28 & ~x29 ;
  assign n42 = ~n40 & n41 ;
  assign n43 = n39 & ~n42 ;
  assign n44 = ~x24 & ~x25 ;
  assign n45 = ~n43 & n44 ;
  assign n46 = n38 & ~n45 ;
  assign n47 = ~x20 & ~x21 ;
  assign n48 = ~n46 & n47 ;
  assign n49 = n37 & ~n48 ;
  assign n50 = ~x16 & ~x17 ;
  assign n51 = ~n49 & n50 ;
  assign n52 = n36 & ~n51 ;
  assign n53 = ~x12 & ~x13 ;
  assign n54 = ~n52 & n53 ;
  assign n55 = n35 & ~n54 ;
  assign n56 = ~x8 & ~x9 ;
  assign n57 = ~n55 & n56 ;
  assign n58 = n34 & ~n57 ;
  assign n59 = ~x4 & ~x5 ;
  assign n60 = ~n58 & n59 ;
  assign n61 = n33 & ~n60 ;
  assign y0 = ~n61 ;
endmodule
