module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 ;
  assign n10 = ~x1 & ~x3 ;
  assign n11 = x4 & x8 ;
  assign n12 = x6 & x8 ;
  assign n13 = ~n11 & ~n12 ;
  assign n14 = n10 & ~n13 ;
  assign n15 = ~x5 & n14 ;
  assign n16 = x5 & x6 ;
  assign n17 = ~x4 & n16 ;
  assign n18 = x5 & n11 ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = n19 ^ x1 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = x6 & ~x8 ;
  assign n23 = ~x5 & n22 ;
  assign n24 = n23 ^ n19 ;
  assign n25 = ~n21 & ~n24 ;
  assign n26 = n25 ^ n19 ;
  assign n27 = x3 & ~n26 ;
  assign n28 = ~n15 & ~n27 ;
  assign n29 = x7 & ~n28 ;
  assign n30 = x1 & ~x4 ;
  assign n31 = n23 & n30 ;
  assign n32 = ~x3 & n31 ;
  assign n33 = ~n29 & ~n32 ;
  assign n34 = ~x1 & x4 ;
  assign n35 = ~x8 & n34 ;
  assign n36 = n16 & n35 ;
  assign n37 = x1 & x6 ;
  assign n38 = x8 & n37 ;
  assign n39 = ~x5 & ~x8 ;
  assign n40 = n34 ^ x4 ;
  assign n41 = n34 ^ x6 ;
  assign n42 = n41 ^ n34 ;
  assign n43 = ~n40 & n42 ;
  assign n44 = n43 ^ n34 ;
  assign n45 = n39 & n44 ;
  assign n46 = ~n38 & ~n45 ;
  assign n47 = ~x3 & ~n46 ;
  assign n48 = ~n36 & ~n47 ;
  assign n49 = x5 & ~x6 ;
  assign n50 = x3 & n49 ;
  assign n51 = n50 ^ n30 ;
  assign n52 = n51 ^ n50 ;
  assign n53 = n52 ^ x8 ;
  assign n54 = n37 ^ n17 ;
  assign n55 = ~n17 & n54 ;
  assign n56 = n55 ^ n50 ;
  assign n57 = n56 ^ n17 ;
  assign n58 = ~n53 & n57 ;
  assign n59 = n58 ^ n55 ;
  assign n60 = n59 ^ n17 ;
  assign n61 = x8 & ~n60 ;
  assign n62 = n61 ^ x8 ;
  assign n63 = n48 & ~n62 ;
  assign n64 = ~x7 & ~n63 ;
  assign n65 = n64 ^ n33 ;
  assign n66 = ~x7 & ~x8 ;
  assign n67 = ~n10 & ~n37 ;
  assign n68 = n66 & ~n67 ;
  assign n94 = x7 & x8 ;
  assign n95 = ~x4 & ~n94 ;
  assign n69 = x8 ^ x3 ;
  assign n75 = n69 ^ x5 ;
  assign n76 = n75 ^ x1 ;
  assign n77 = n76 ^ x1 ;
  assign n78 = n69 ^ x8 ;
  assign n79 = n78 ^ n69 ;
  assign n80 = n79 ^ x1 ;
  assign n81 = ~n77 & ~n80 ;
  assign n70 = n69 ^ x7 ;
  assign n71 = n70 ^ n69 ;
  assign n72 = n71 ^ x5 ;
  assign n73 = n72 ^ x1 ;
  assign n74 = ~x5 & n73 ;
  assign n82 = n81 ^ n74 ;
  assign n83 = n82 ^ x5 ;
  assign n84 = n74 ^ x1 ;
  assign n85 = n84 ^ n76 ;
  assign n86 = ~x1 & ~n85 ;
  assign n87 = n86 ^ n74 ;
  assign n88 = ~n83 & n87 ;
  assign n89 = n88 ^ n81 ;
  assign n90 = n89 ^ n86 ;
  assign n91 = n90 ^ x5 ;
  assign n92 = n91 ^ x1 ;
  assign n93 = n92 ^ n76 ;
  assign n96 = n95 ^ n93 ;
  assign n97 = n96 ^ x6 ;
  assign n104 = n97 ^ n96 ;
  assign n98 = n97 ^ x4 ;
  assign n99 = n98 ^ n96 ;
  assign n100 = n97 ^ n93 ;
  assign n101 = n100 ^ x4 ;
  assign n102 = n101 ^ n99 ;
  assign n103 = n99 & n102 ;
  assign n105 = n104 ^ n103 ;
  assign n106 = n105 ^ n99 ;
  assign n107 = n96 ^ x5 ;
  assign n108 = n103 ^ n99 ;
  assign n109 = n107 & n108 ;
  assign n110 = n109 ^ n96 ;
  assign n111 = ~n106 & ~n110 ;
  assign n112 = n111 ^ n96 ;
  assign n113 = n112 ^ n95 ;
  assign n114 = n113 ^ n96 ;
  assign n115 = ~n68 & n114 ;
  assign n116 = ~x6 & n66 ;
  assign n117 = x3 & ~x5 ;
  assign n118 = ~x7 & n117 ;
  assign n119 = ~n116 & ~n118 ;
  assign n120 = x1 & ~n119 ;
  assign n121 = ~x5 & x6 ;
  assign n122 = ~x7 & x8 ;
  assign n123 = n121 & n122 ;
  assign n124 = x8 ^ x7 ;
  assign n125 = n124 ^ n49 ;
  assign n126 = x8 ^ x1 ;
  assign n127 = n49 ^ x1 ;
  assign n128 = ~n126 & n127 ;
  assign n129 = n128 ^ x1 ;
  assign n130 = n125 & n129 ;
  assign n131 = n130 ^ n49 ;
  assign n132 = ~x3 & ~n131 ;
  assign n133 = ~n123 & n132 ;
  assign n138 = x7 ^ x1 ;
  assign n134 = n16 ^ x1 ;
  assign n135 = n134 ^ n22 ;
  assign n136 = n135 ^ x7 ;
  assign n137 = n136 ^ n134 ;
  assign n139 = n138 ^ n137 ;
  assign n140 = n134 ^ x3 ;
  assign n141 = ~n139 & ~n140 ;
  assign n142 = n141 ^ n134 ;
  assign n143 = n142 ^ n136 ;
  assign n144 = n143 ^ x3 ;
  assign n145 = n138 ^ x1 ;
  assign n146 = ~x3 & ~n145 ;
  assign n147 = n146 ^ n134 ;
  assign n148 = n147 ^ n136 ;
  assign n149 = n148 ^ x1 ;
  assign n150 = n149 ^ x3 ;
  assign n151 = n134 ^ n39 ;
  assign n152 = n151 ^ n138 ;
  assign n153 = n152 ^ x3 ;
  assign n154 = n151 & n153 ;
  assign n155 = n154 ^ n136 ;
  assign n156 = n155 ^ x3 ;
  assign n157 = ~n150 & ~n156 ;
  assign n158 = n157 ^ n136 ;
  assign n159 = ~n144 & n158 ;
  assign n160 = n159 ^ n146 ;
  assign n161 = n160 ^ n141 ;
  assign n162 = n161 ^ n134 ;
  assign n163 = n162 ^ n136 ;
  assign n164 = n163 ^ x1 ;
  assign n165 = n164 ^ n138 ;
  assign n166 = n165 ^ x3 ;
  assign n167 = ~n133 & ~n166 ;
  assign n168 = x4 & ~n167 ;
  assign n169 = ~n120 & n168 ;
  assign n170 = ~n115 & ~n169 ;
  assign n171 = n94 & n117 ;
  assign n172 = ~x6 & n171 ;
  assign n173 = ~n170 & ~n172 ;
  assign n174 = n173 ^ x2 ;
  assign n175 = n174 ^ n173 ;
  assign n176 = x1 & x7 ;
  assign n177 = ~n34 & ~n176 ;
  assign n178 = ~n95 & n177 ;
  assign n179 = x3 & ~n66 ;
  assign n180 = ~n94 & n179 ;
  assign n181 = ~n178 & ~n180 ;
  assign n182 = n121 & ~n181 ;
  assign n183 = ~x4 & ~x5 ;
  assign n184 = x7 & ~x8 ;
  assign n185 = ~x6 & n184 ;
  assign n186 = n183 & n185 ;
  assign n187 = ~n182 & ~n186 ;
  assign n188 = x4 & x5 ;
  assign n189 = x7 & ~n188 ;
  assign n190 = n38 & ~n189 ;
  assign n191 = n190 ^ n187 ;
  assign n192 = ~x4 & x8 ;
  assign n193 = n49 & ~n192 ;
  assign n194 = ~n94 & n193 ;
  assign n195 = ~x1 & n194 ;
  assign n196 = x7 & n49 ;
  assign n197 = ~x4 & n196 ;
  assign n198 = x5 ^ x4 ;
  assign n199 = n66 ^ x5 ;
  assign n200 = n199 ^ n66 ;
  assign n201 = n122 ^ n66 ;
  assign n202 = ~n200 & n201 ;
  assign n203 = n202 ^ n66 ;
  assign n204 = ~n198 & n203 ;
  assign n205 = ~n197 & ~n204 ;
  assign n206 = ~n195 & n205 ;
  assign n207 = n206 ^ x3 ;
  assign n208 = n207 ^ n206 ;
  assign n209 = n49 & n192 ;
  assign n210 = x4 ^ x1 ;
  assign n211 = n210 ^ x4 ;
  assign n212 = n183 ^ x4 ;
  assign n213 = n211 & ~n212 ;
  assign n214 = n213 ^ x4 ;
  assign n215 = ~x8 & n214 ;
  assign n216 = n215 ^ x1 ;
  assign n219 = n216 ^ n30 ;
  assign n220 = n219 ^ n216 ;
  assign n217 = n216 ^ n121 ;
  assign n218 = n217 ^ n216 ;
  assign n221 = n220 ^ n218 ;
  assign n222 = n216 ^ n188 ;
  assign n223 = n222 ^ n216 ;
  assign n224 = n223 ^ n220 ;
  assign n225 = ~n220 & n224 ;
  assign n226 = n225 ^ n220 ;
  assign n227 = n221 & ~n226 ;
  assign n228 = n227 ^ n225 ;
  assign n229 = n228 ^ n216 ;
  assign n230 = n229 ^ n220 ;
  assign n231 = x7 & ~n230 ;
  assign n232 = n231 ^ n216 ;
  assign n233 = ~n209 & ~n232 ;
  assign n234 = n233 ^ n206 ;
  assign n235 = ~n208 & n234 ;
  assign n236 = n235 ^ n206 ;
  assign n237 = n236 ^ n187 ;
  assign n238 = ~n191 & n237 ;
  assign n239 = n238 ^ n235 ;
  assign n240 = n239 ^ n206 ;
  assign n241 = n240 ^ n190 ;
  assign n242 = n187 & ~n241 ;
  assign n243 = n242 ^ n187 ;
  assign n244 = n243 ^ n173 ;
  assign n245 = ~n175 & n244 ;
  assign n246 = n245 ^ n173 ;
  assign n247 = n246 ^ n33 ;
  assign n248 = ~n65 & n247 ;
  assign n249 = n248 ^ n245 ;
  assign n250 = n249 ^ n173 ;
  assign n251 = n250 ^ n64 ;
  assign n252 = n33 & ~n251 ;
  assign n253 = n252 ^ n33 ;
  assign n254 = ~x0 & ~n253 ;
  assign n255 = x4 & x6 ;
  assign n256 = ~x7 & n255 ;
  assign n257 = n121 & n184 ;
  assign n258 = x6 ^ x4 ;
  assign n259 = n66 & n258 ;
  assign n260 = n259 ^ x4 ;
  assign n261 = ~n257 & ~n260 ;
  assign n262 = x0 & ~n261 ;
  assign n263 = ~n256 & n262 ;
  assign n264 = n122 & n255 ;
  assign n265 = x5 & n264 ;
  assign n266 = ~n197 & ~n265 ;
  assign n267 = ~n263 & n266 ;
  assign n268 = ~x2 & n10 ;
  assign n269 = ~n267 & n268 ;
  assign n270 = ~n254 & ~n269 ;
  assign y0 = ~n270 ;
endmodule
