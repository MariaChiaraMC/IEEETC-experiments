module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 ;
  assign n8 = ~x0 & x2 ;
  assign n9 = x5 & x6 ;
  assign n10 = x4 & n9 ;
  assign n11 = n8 & n10 ;
  assign n12 = ~x3 & n11 ;
  assign n52 = ~x3 & ~x4 ;
  assign n53 = ~n9 & ~n52 ;
  assign n54 = x0 & ~n53 ;
  assign n55 = ~x4 & ~x6 ;
  assign n56 = x3 & ~x5 ;
  assign n57 = ~x6 & ~n56 ;
  assign n58 = ~x5 & n57 ;
  assign n59 = n58 ^ n56 ;
  assign n60 = ~n55 & n59 ;
  assign n61 = ~n54 & ~n60 ;
  assign n62 = x6 ^ x0 ;
  assign n30 = x3 ^ x0 ;
  assign n63 = ~x5 & n55 ;
  assign n64 = n63 ^ x0 ;
  assign n65 = ~x0 & n64 ;
  assign n66 = n65 ^ x0 ;
  assign n67 = n30 & ~n66 ;
  assign n68 = n67 ^ n65 ;
  assign n69 = n68 ^ x0 ;
  assign n70 = n69 ^ n63 ;
  assign n71 = ~n62 & n70 ;
  assign n72 = n71 ^ n63 ;
  assign n73 = x2 & n72 ;
  assign n74 = ~n61 & ~n73 ;
  assign n75 = ~x4 & n8 ;
  assign n76 = ~n57 & n75 ;
  assign n37 = x3 & x4 ;
  assign n77 = x5 & ~n37 ;
  assign n78 = x0 & x2 ;
  assign n79 = ~n59 & n78 ;
  assign n80 = ~n77 & n79 ;
  assign n81 = ~n76 & ~n80 ;
  assign n82 = ~n74 & n81 ;
  assign n13 = x4 ^ x3 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = n14 ^ x5 ;
  assign n16 = x5 ^ x4 ;
  assign n17 = n14 ^ x0 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = ~x5 & ~n18 ;
  assign n20 = n19 ^ x5 ;
  assign n21 = n16 & ~n20 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ x5 ;
  assign n24 = n23 ^ n17 ;
  assign n25 = ~n15 & ~n24 ;
  assign n26 = n25 ^ n14 ;
  assign n27 = ~x6 & ~n26 ;
  assign n28 = ~x0 & ~x2 ;
  assign n29 = ~x4 & ~n28 ;
  assign n31 = ~x2 & n30 ;
  assign n32 = n31 ^ x0 ;
  assign n33 = x6 & ~n32 ;
  assign n34 = ~n29 & n33 ;
  assign n35 = ~x5 & n34 ;
  assign n36 = x0 & x6 ;
  assign n38 = ~x4 & x5 ;
  assign n39 = x2 & n38 ;
  assign n40 = ~n37 & ~n39 ;
  assign n41 = n36 & ~n40 ;
  assign n42 = x3 & ~x4 ;
  assign n43 = n28 ^ x5 ;
  assign n44 = n43 ^ n28 ;
  assign n45 = n28 ^ x0 ;
  assign n46 = ~n44 & n45 ;
  assign n47 = n46 ^ n28 ;
  assign n48 = n42 & n47 ;
  assign n49 = ~n41 & ~n48 ;
  assign n50 = ~n35 & n49 ;
  assign n51 = ~n27 & n50 ;
  assign n83 = n82 ^ n51 ;
  assign n84 = x1 & n83 ;
  assign n85 = n84 ^ n82 ;
  assign n86 = ~n12 & n85 ;
  assign y0 = ~n86 ;
endmodule
