module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 ;
  assign n9 = x1 & ~x2 ;
  assign n10 = ~x4 & ~x7 ;
  assign n11 = ~x5 & ~x6 ;
  assign n12 = ~x0 & n11 ;
  assign n13 = n10 & n12 ;
  assign n14 = n9 & n13 ;
  assign n15 = ~x4 & x7 ;
  assign n16 = ~x0 & x2 ;
  assign n17 = x5 & x6 ;
  assign n18 = n17 ^ n11 ;
  assign n19 = x1 & n18 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n16 & n20 ;
  assign n22 = ~x5 & x6 ;
  assign n23 = n9 & n22 ;
  assign n24 = ~n21 & ~n23 ;
  assign n25 = n15 & n24 ;
  assign n42 = x1 ^ x0 ;
  assign n43 = x4 ^ x1 ;
  assign n44 = ~n42 & ~n43 ;
  assign n45 = x2 & n18 ;
  assign n46 = n45 ^ n17 ;
  assign n47 = n44 & n46 ;
  assign n26 = x0 & x1 ;
  assign n27 = ~x5 & ~n26 ;
  assign n28 = n16 ^ x1 ;
  assign n29 = ~x6 & ~n28 ;
  assign n30 = n29 ^ x1 ;
  assign n31 = n27 & n30 ;
  assign n32 = x0 & x5 ;
  assign n33 = x1 & x6 ;
  assign n34 = n33 ^ x2 ;
  assign n35 = n34 ^ n33 ;
  assign n36 = n33 ^ x1 ;
  assign n37 = ~n35 & ~n36 ;
  assign n38 = n37 ^ n33 ;
  assign n39 = n32 & n38 ;
  assign n40 = x4 & ~n39 ;
  assign n41 = ~n31 & n40 ;
  assign n48 = n47 ^ n41 ;
  assign n49 = n48 ^ n41 ;
  assign n50 = x4 & ~x6 ;
  assign n51 = x1 & x2 ;
  assign n52 = ~x0 & x5 ;
  assign n53 = n51 & n52 ;
  assign n54 = ~n50 & n53 ;
  assign n55 = n54 ^ n41 ;
  assign n56 = n55 ^ n41 ;
  assign n57 = ~n49 & ~n56 ;
  assign n58 = n57 ^ n41 ;
  assign n59 = ~x7 & n58 ;
  assign n60 = n59 ^ n41 ;
  assign n61 = ~n25 & ~n60 ;
  assign n62 = n61 ^ x3 ;
  assign n63 = n62 ^ n61 ;
  assign n64 = x4 & ~x7 ;
  assign n65 = n11 & n64 ;
  assign n66 = n15 & n17 ;
  assign n67 = ~n65 & ~n66 ;
  assign n68 = n26 & ~n67 ;
  assign n69 = ~x1 & ~x4 ;
  assign n70 = x0 & n69 ;
  assign n71 = n22 & n70 ;
  assign n72 = ~x7 & n71 ;
  assign n73 = ~n68 & ~n72 ;
  assign n74 = ~x1 & n17 ;
  assign n75 = x7 & n74 ;
  assign n76 = ~x0 & n75 ;
  assign n77 = ~n13 & ~n76 ;
  assign n78 = ~n10 & ~n50 ;
  assign n79 = n52 & ~n78 ;
  assign n80 = x1 & n79 ;
  assign n81 = ~x2 & ~n80 ;
  assign n82 = n77 & n81 ;
  assign n83 = n73 & n82 ;
  assign n84 = x7 ^ x4 ;
  assign n85 = x6 ^ x5 ;
  assign n86 = n85 ^ n84 ;
  assign n87 = x7 ^ x6 ;
  assign n88 = n87 ^ x6 ;
  assign n89 = x6 ^ x0 ;
  assign n90 = n89 ^ x6 ;
  assign n91 = n88 & ~n90 ;
  assign n92 = n91 ^ x6 ;
  assign n93 = n92 ^ n84 ;
  assign n94 = n86 & n93 ;
  assign n95 = n94 ^ n91 ;
  assign n96 = n95 ^ x6 ;
  assign n97 = n96 ^ n85 ;
  assign n98 = n84 & n97 ;
  assign n99 = n98 ^ n84 ;
  assign n100 = x1 & n99 ;
  assign n101 = n17 ^ x7 ;
  assign n102 = n101 ^ n17 ;
  assign n103 = n18 & n102 ;
  assign n104 = n103 ^ n17 ;
  assign n105 = n70 & n104 ;
  assign n106 = x2 & ~n105 ;
  assign n107 = ~n100 & n106 ;
  assign n108 = ~n83 & ~n107 ;
  assign n109 = n108 ^ n61 ;
  assign n110 = ~n63 & n109 ;
  assign n111 = n110 ^ n61 ;
  assign n112 = ~n14 & ~n111 ;
  assign y0 = ~n112 ;
endmodule
