module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;
  assign n16 = x7 & x8 ;
  assign n17 = ~x2 & ~x9 ;
  assign n18 = ~x4 & ~x6 ;
  assign n19 = n17 & n18 ;
  assign n20 = ~x1 & ~x12 ;
  assign n21 = ~x0 & n20 ;
  assign n22 = n19 & n21 ;
  assign n23 = ~n16 & n22 ;
  assign n24 = ~x11 & ~x14 ;
  assign n25 = x10 & ~n24 ;
  assign n26 = ~x7 & ~x8 ;
  assign n27 = x5 & ~n26 ;
  assign n28 = ~n25 & ~n27 ;
  assign n29 = ~x13 & n28 ;
  assign n30 = n23 & n29 ;
  assign n32 = ~x5 & n26 ;
  assign n31 = ~x10 & ~x11 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = n31 ^ x14 ;
  assign n35 = n31 ^ x3 ;
  assign n36 = n31 & ~n35 ;
  assign n37 = n36 ^ n31 ;
  assign n38 = ~n34 & n37 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n39 ^ n31 ;
  assign n41 = n40 ^ x3 ;
  assign n42 = n33 & ~n41 ;
  assign n43 = n30 & n42 ;
  assign y0 = n43 ;
endmodule
