module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 ;
  assign n9 = x2 & x4 ;
  assign n10 = x1 & ~n9 ;
  assign n11 = x0 & n10 ;
  assign n12 = ~x0 & ~x5 ;
  assign n13 = ~x1 & x7 ;
  assign n14 = n13 ^ x4 ;
  assign n15 = n14 ^ x4 ;
  assign n16 = x4 ^ x2 ;
  assign n17 = n16 ^ x4 ;
  assign n18 = n15 & ~n17 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = ~x6 & n19 ;
  assign n21 = n20 ^ x4 ;
  assign n22 = n12 & n21 ;
  assign n23 = ~x4 & ~x5 ;
  assign n24 = x6 & x7 ;
  assign n25 = x1 & ~n24 ;
  assign n26 = x6 ^ x2 ;
  assign n27 = ~n25 & n26 ;
  assign n28 = n23 & ~n27 ;
  assign n30 = ~x7 & n23 ;
  assign n29 = x1 & n9 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = ~x1 & x2 ;
  assign n34 = n33 ^ n29 ;
  assign n35 = n34 ^ n29 ;
  assign n36 = ~n32 & ~n35 ;
  assign n37 = n36 ^ n29 ;
  assign n38 = x0 & ~n37 ;
  assign n39 = n38 ^ n29 ;
  assign n40 = ~n28 & ~n39 ;
  assign n41 = ~n22 & n40 ;
  assign n42 = n41 ^ x3 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = x1 ^ x0 ;
  assign n46 = n44 ^ x2 ;
  assign n45 = n44 ^ x4 ;
  assign n47 = n46 ^ n45 ;
  assign n48 = n47 ^ x1 ;
  assign n49 = n46 ^ x1 ;
  assign n50 = n49 ^ n44 ;
  assign n52 = n50 ^ n44 ;
  assign n51 = n50 ^ x1 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = ~n48 & ~n53 ;
  assign n55 = n54 ^ n50 ;
  assign n56 = n55 ^ n52 ;
  assign n57 = n44 ^ x6 ;
  assign n58 = n57 ^ x1 ;
  assign n59 = n58 ^ n50 ;
  assign n60 = n59 ^ n52 ;
  assign n61 = n58 ^ n47 ;
  assign n62 = n61 ^ n52 ;
  assign n63 = ~n60 & n62 ;
  assign n64 = n63 ^ n50 ;
  assign n65 = n64 ^ x1 ;
  assign n66 = n65 ^ n58 ;
  assign n67 = n66 ^ n52 ;
  assign n68 = n58 ^ n51 ;
  assign n69 = n68 ^ n52 ;
  assign n70 = ~x7 & ~n69 ;
  assign n71 = n70 ^ x7 ;
  assign n72 = n71 ^ x1 ;
  assign n73 = n72 ^ n58 ;
  assign n74 = n73 ^ n52 ;
  assign n75 = ~n67 & n74 ;
  assign n76 = n75 ^ x1 ;
  assign n77 = n76 ^ n52 ;
  assign n78 = ~n56 & ~n77 ;
  assign n79 = n78 ^ n75 ;
  assign n80 = n79 ^ x1 ;
  assign n81 = n80 ^ n52 ;
  assign n82 = n81 ^ x0 ;
  assign n83 = n82 ^ n41 ;
  assign n84 = ~n43 & n83 ;
  assign n85 = n84 ^ n41 ;
  assign n86 = ~n11 & n85 ;
  assign n87 = ~x6 & ~x7 ;
  assign n88 = ~x3 & n87 ;
  assign n89 = ~x2 & x4 ;
  assign n90 = x1 & n89 ;
  assign n91 = ~n88 & n90 ;
  assign n92 = ~x2 & ~x4 ;
  assign n93 = ~x4 & ~x6 ;
  assign n94 = ~n92 & ~n93 ;
  assign n95 = ~x1 & x3 ;
  assign n96 = ~n24 & n95 ;
  assign n97 = ~n94 & n96 ;
  assign n98 = x6 & ~x7 ;
  assign n99 = x4 & n26 ;
  assign n100 = ~n98 & n99 ;
  assign n101 = ~n97 & ~n100 ;
  assign n102 = ~x0 & ~n101 ;
  assign n103 = ~n91 & ~n102 ;
  assign n104 = x1 & n92 ;
  assign n105 = x6 ^ x4 ;
  assign n106 = n105 ^ x7 ;
  assign n107 = n106 ^ n105 ;
  assign n108 = n105 ^ x6 ;
  assign n109 = n108 ^ n105 ;
  assign n110 = n107 & ~n109 ;
  assign n111 = n110 ^ n105 ;
  assign n112 = ~x2 & ~n105 ;
  assign n113 = n112 ^ x1 ;
  assign n114 = ~n111 & ~n113 ;
  assign n115 = n114 ^ n112 ;
  assign n116 = ~x1 & n115 ;
  assign n117 = n116 ^ x1 ;
  assign n118 = n117 ^ x0 ;
  assign n119 = n118 ^ n117 ;
  assign n120 = n119 ^ n104 ;
  assign n121 = x2 & ~x4 ;
  assign n122 = x2 & ~x6 ;
  assign n123 = ~x7 & n122 ;
  assign n124 = n123 ^ n121 ;
  assign n125 = ~n121 & n124 ;
  assign n126 = n125 ^ n117 ;
  assign n127 = n126 ^ n121 ;
  assign n128 = ~n120 & n127 ;
  assign n129 = n128 ^ n125 ;
  assign n130 = n129 ^ n121 ;
  assign n131 = ~n104 & ~n130 ;
  assign n132 = n131 ^ n104 ;
  assign n133 = n132 ^ x3 ;
  assign n134 = n133 ^ n132 ;
  assign n135 = n134 ^ n103 ;
  assign n136 = n123 ^ x4 ;
  assign n137 = ~x4 & ~n136 ;
  assign n138 = n137 ^ n132 ;
  assign n139 = n138 ^ x4 ;
  assign n140 = n135 & ~n139 ;
  assign n141 = n140 ^ n137 ;
  assign n142 = n141 ^ x4 ;
  assign n143 = n103 & ~n142 ;
  assign n144 = n143 ^ n103 ;
  assign n145 = n144 ^ x5 ;
  assign n146 = n145 ^ n144 ;
  assign n147 = n146 ^ n86 ;
  assign n148 = x4 & x6 ;
  assign n149 = n13 & n148 ;
  assign n150 = ~x4 & n122 ;
  assign n151 = ~x3 & n150 ;
  assign n152 = ~n149 & ~n151 ;
  assign n153 = n152 ^ x0 ;
  assign n154 = ~n152 & n153 ;
  assign n155 = n154 ^ n144 ;
  assign n156 = n155 ^ n152 ;
  assign n157 = ~n147 & n156 ;
  assign n158 = n157 ^ n154 ;
  assign n159 = n158 ^ n152 ;
  assign n160 = n86 & ~n159 ;
  assign n161 = n160 ^ n86 ;
  assign y0 = ~n161 ;
endmodule
