module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 ;
  assign n16 = ~x3 & x4 ;
  assign n17 = ~x2 & ~n16 ;
  assign n18 = n17 ^ x13 ;
  assign n19 = n18 ^ n17 ;
  assign n30 = x6 ^ x4 ;
  assign n31 = x5 & ~n30 ;
  assign n32 = n31 ^ x4 ;
  assign n33 = x3 ^ x1 ;
  assign n34 = x6 ^ x3 ;
  assign n20 = x6 ^ x2 ;
  assign n35 = x6 & n20 ;
  assign n36 = n35 ^ x6 ;
  assign n37 = ~n34 & n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = n38 ^ x6 ;
  assign n40 = n39 ^ x2 ;
  assign n41 = ~n33 & n40 ;
  assign n42 = n32 & n41 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = x5 ^ x2 ;
  assign n23 = n22 ^ x2 ;
  assign n24 = ~n21 & n23 ;
  assign n25 = n24 ^ x2 ;
  assign n26 = ~x1 & ~n25 ;
  assign n27 = n26 ^ x2 ;
  assign n43 = n42 ^ n27 ;
  assign n28 = ~x2 & ~x3 ;
  assign n29 = n28 ^ n27 ;
  assign n44 = n43 ^ n29 ;
  assign n45 = ~x1 & x5 ;
  assign n46 = n45 ^ n43 ;
  assign n47 = n46 ^ n43 ;
  assign n48 = n44 & n47 ;
  assign n49 = n48 ^ n43 ;
  assign n50 = x0 & ~n49 ;
  assign n51 = n50 ^ n27 ;
  assign n52 = n51 ^ n17 ;
  assign n53 = ~n19 & ~n52 ;
  assign n54 = n53 ^ n17 ;
  assign n55 = ~x9 & n54 ;
  assign n56 = ~x10 & ~n55 ;
  assign n57 = x11 ^ x9 ;
  assign n58 = n57 ^ x9 ;
  assign n59 = n58 ^ x13 ;
  assign n60 = x0 & ~x1 ;
  assign n61 = ~n28 & n60 ;
  assign n62 = x14 & ~n61 ;
  assign n63 = n62 ^ x10 ;
  assign n64 = x10 & ~n63 ;
  assign n65 = n64 ^ x9 ;
  assign n66 = n65 ^ x10 ;
  assign n67 = n59 & n66 ;
  assign n68 = n67 ^ n64 ;
  assign n69 = n68 ^ x10 ;
  assign n70 = ~x13 & n69 ;
  assign n71 = n70 ^ x11 ;
  assign n72 = ~n56 & ~n71 ;
  assign y0 = n72 ;
endmodule
