module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 ;
  assign n9 = ~x0 & x2 ;
  assign n10 = ~x7 & ~n9 ;
  assign n11 = ~x5 & n10 ;
  assign n12 = x4 & ~n11 ;
  assign n13 = ~x3 & ~n12 ;
  assign n14 = x1 ^ x0 ;
  assign n15 = x4 ^ x1 ;
  assign n16 = n15 ^ x1 ;
  assign n17 = n14 & ~n16 ;
  assign n18 = n17 ^ x1 ;
  assign n19 = n15 ^ x2 ;
  assign n20 = n19 ^ x7 ;
  assign n21 = n20 ^ n15 ;
  assign n22 = n21 ^ x1 ;
  assign n23 = n15 ^ x5 ;
  assign n27 = n23 ^ n15 ;
  assign n24 = n23 ^ x7 ;
  assign n25 = ~x1 & ~n24 ;
  assign n26 = n25 ^ n17 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = n28 ^ n24 ;
  assign n30 = n29 ^ x1 ;
  assign n31 = n22 & ~n30 ;
  assign n32 = n31 ^ n16 ;
  assign n33 = ~n18 & ~n32 ;
  assign n34 = n33 ^ n17 ;
  assign n35 = n34 ^ n16 ;
  assign n36 = n35 ^ x4 ;
  assign n37 = n36 ^ n15 ;
  assign n38 = n13 & ~n37 ;
  assign n39 = ~x1 & ~x4 ;
  assign n41 = x2 & x7 ;
  assign n40 = ~x2 & ~x7 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = n41 ^ x3 ;
  assign n45 = n44 ^ n41 ;
  assign n46 = n43 & n45 ;
  assign n47 = n46 ^ n41 ;
  assign n48 = x5 & n47 ;
  assign n49 = n48 ^ n41 ;
  assign n50 = n39 & n49 ;
  assign n51 = x0 & n50 ;
  assign n52 = ~n38 & ~n51 ;
  assign y0 = ~n52 ;
endmodule
