// Benchmark "./spla.pla" written by ABC on Thu Apr 23 11:00:03 2020

module \./spla.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15,
    z44  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15;
  output z44;
  wire new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_, new_n24_,
    new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_, new_n31_,
    new_n32_, new_n33_;
  assign new_n18_ = x5 & ~x7;
  assign new_n19_ = x5 & ~x6;
  assign new_n20_ = x10 & x11;
  assign new_n21_ = new_n19_ & ~new_n20_;
  assign new_n22_ = ~x10 & ~x11;
  assign new_n23_ = ~x8 & ~x9;
  assign new_n24_ = ~new_n22_ & new_n23_;
  assign new_n25_ = new_n21_ & new_n24_;
  assign new_n26_ = ~new_n18_ & ~new_n25_;
  assign new_n27_ = new_n19_ & new_n22_;
  assign new_n28_ = x6 & x7;
  assign new_n29_ = ~x5 & new_n28_;
  assign new_n30_ = ~new_n27_ & ~new_n29_;
  assign new_n31_ = x8 & x9;
  assign new_n32_ = ~new_n23_ & ~new_n31_;
  assign new_n33_ = ~new_n30_ & new_n32_;
  assign z44 = ~new_n26_ | new_n33_;
endmodule


