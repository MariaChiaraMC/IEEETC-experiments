module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 ;
  assign n17 = ~x4 & ~x5 ;
  assign n18 = ~x1 & ~x3 ;
  assign n19 = n17 & n18 ;
  assign n20 = ~x6 & n19 ;
  assign n21 = ~x9 & ~x10 ;
  assign n22 = x14 & x15 ;
  assign n23 = n21 & n22 ;
  assign n24 = ~x2 & n23 ;
  assign n25 = n20 & n24 ;
  assign n26 = x6 & x9 ;
  assign n27 = ~x10 & ~x15 ;
  assign n28 = n26 & n27 ;
  assign n29 = n19 & n28 ;
  assign n30 = x5 & ~x6 ;
  assign n31 = ~x1 & n30 ;
  assign n32 = ~x9 & x10 ;
  assign n33 = ~x15 & n32 ;
  assign n34 = n31 & n33 ;
  assign n35 = x6 & x10 ;
  assign n36 = x9 & x15 ;
  assign n37 = x1 & n36 ;
  assign n38 = ~n35 & n37 ;
  assign n39 = ~n34 & ~n38 ;
  assign n40 = x3 & x4 ;
  assign n41 = ~n39 & n40 ;
  assign n42 = ~n29 & ~n41 ;
  assign n43 = x2 & ~x14 ;
  assign n44 = ~n42 & n43 ;
  assign n45 = ~n25 & ~n44 ;
  assign n46 = ~x7 & ~n45 ;
  assign n47 = x2 & x4 ;
  assign n54 = ~x5 & ~x14 ;
  assign n48 = x10 & x14 ;
  assign n49 = n31 & n48 ;
  assign n55 = n54 ^ n49 ;
  assign n56 = n55 ^ n49 ;
  assign n50 = x7 & x10 ;
  assign n51 = x6 & ~n50 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = n52 ^ n49 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n49 ^ x1 ;
  assign n59 = n58 ^ n49 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = n56 & n60 ;
  assign n62 = n61 ^ n56 ;
  assign n63 = ~n57 & n62 ;
  assign n64 = n63 ^ n61 ;
  assign n65 = n64 ^ n49 ;
  assign n66 = n65 ^ n56 ;
  assign n67 = x3 & n66 ;
  assign n68 = n67 ^ n49 ;
  assign n69 = n47 & n68 ;
  assign n70 = n36 & n69 ;
  assign n71 = ~n46 & ~n70 ;
  assign n72 = ~x8 & ~n71 ;
  assign n73 = ~x2 & ~n50 ;
  assign n74 = x8 & n26 ;
  assign n75 = n18 & n74 ;
  assign n76 = x11 & n48 ;
  assign n77 = n76 ^ x14 ;
  assign n78 = n77 ^ n76 ;
  assign n79 = n76 ^ x7 ;
  assign n80 = n79 ^ n76 ;
  assign n81 = ~n78 & n80 ;
  assign n82 = n81 ^ n76 ;
  assign n83 = x15 & n82 ;
  assign n84 = n83 ^ n76 ;
  assign n85 = n75 & n84 ;
  assign n86 = n73 & n85 ;
  assign n87 = n17 & n86 ;
  assign n88 = ~n72 & ~n87 ;
  assign n89 = ~x13 & ~n88 ;
  assign n90 = ~x8 & x9 ;
  assign n91 = n47 & n90 ;
  assign n92 = ~x14 & x15 ;
  assign n93 = x10 & x13 ;
  assign n94 = n92 & n93 ;
  assign n95 = n31 & n94 ;
  assign n96 = n91 & n95 ;
  assign n97 = ~x3 & n96 ;
  assign n98 = ~n89 & ~n97 ;
  assign n99 = ~x0 & ~n98 ;
  assign n100 = ~x12 & n99 ;
  assign y0 = n100 ;
endmodule
