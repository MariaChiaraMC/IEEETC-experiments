module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 ;
  assign n7 = x5 ^ x4 ;
  assign n9 = n7 ^ x3 ;
  assign n10 = n9 ^ x5 ;
  assign n8 = n7 ^ x0 ;
  assign n11 = n10 ^ n8 ;
  assign n12 = n11 ^ n7 ;
  assign n13 = n12 ^ n11 ;
  assign n22 = n11 ^ n10 ;
  assign n20 = n11 ^ n9 ;
  assign n14 = n7 ^ x2 ;
  assign n15 = n14 ^ n9 ;
  assign n16 = n15 ^ n10 ;
  assign n17 = n16 ^ n10 ;
  assign n18 = n17 ^ n7 ;
  assign n19 = n18 ^ n12 ;
  assign n21 = n20 ^ n19 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n13 & ~n23 ;
  assign n25 = n24 ^ n18 ;
  assign n26 = n25 ^ n11 ;
  assign n27 = n16 ^ x1 ;
  assign n28 = n27 ^ n16 ;
  assign n29 = n28 ^ n9 ;
  assign n30 = n29 ^ n11 ;
  assign n31 = n30 ^ n12 ;
  assign n32 = ~n20 & ~n31 ;
  assign n33 = n32 ^ n18 ;
  assign n34 = n33 ^ n29 ;
  assign n35 = n34 ^ n11 ;
  assign n36 = n35 ^ n12 ;
  assign n37 = n36 ^ n22 ;
  assign n38 = n18 ^ n11 ;
  assign n39 = n38 ^ n12 ;
  assign n40 = n39 ^ n22 ;
  assign n41 = n22 ^ n18 ;
  assign n42 = n40 & n41 ;
  assign n43 = n42 ^ n18 ;
  assign n44 = ~n37 & ~n43 ;
  assign n45 = n44 ^ n18 ;
  assign n46 = n45 ^ n12 ;
  assign n47 = ~n26 & ~n46 ;
  assign n48 = n47 ^ n42 ;
  assign n49 = n48 ^ n24 ;
  assign n50 = n49 ^ n44 ;
  assign n51 = n50 ^ n11 ;
  assign n52 = n51 ^ n22 ;
  assign n53 = n52 ^ n7 ;
  assign y0 = ~n53 ;
endmodule
