module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 ;
  assign n9 = ~x0 & x5 ;
  assign n10 = x6 & x7 ;
  assign n11 = n9 & ~n10 ;
  assign n12 = n11 ^ x0 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n11 ^ x2 ;
  assign n15 = n13 & ~n14 ;
  assign n16 = n15 ^ n11 ;
  assign n17 = ~x3 & ~x5 ;
  assign n18 = ~x6 & x7 ;
  assign n19 = n17 & n18 ;
  assign n20 = ~n11 & ~n19 ;
  assign n21 = n20 ^ x4 ;
  assign n22 = ~n16 & n21 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = x4 & n23 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = n25 ^ x3 ;
  assign n27 = x2 & x6 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = ~x4 & n27 ;
  assign n32 = x7 & n31 ;
  assign n33 = ~x0 & ~x5 ;
  assign n34 = n33 ^ n32 ;
  assign n35 = n32 & n34 ;
  assign n36 = n35 ^ n27 ;
  assign n37 = n36 ^ n32 ;
  assign n38 = n30 & n37 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n39 ^ n32 ;
  assign n41 = ~n26 & n40 ;
  assign n42 = n41 ^ n25 ;
  assign n43 = x4 & x5 ;
  assign n44 = ~x2 & ~x6 ;
  assign n45 = n43 & n44 ;
  assign n46 = n45 ^ x0 ;
  assign n47 = n46 ^ n32 ;
  assign n48 = x3 & x7 ;
  assign n49 = n48 ^ x5 ;
  assign n50 = n45 & n49 ;
  assign n51 = n50 ^ x5 ;
  assign n52 = n47 & n51 ;
  assign n53 = n52 ^ n50 ;
  assign n54 = n53 ^ x5 ;
  assign n55 = n54 ^ n45 ;
  assign n56 = ~n32 & n55 ;
  assign n57 = x5 ^ x4 ;
  assign n58 = x0 & n57 ;
  assign n59 = x2 & x3 ;
  assign n60 = n10 & n59 ;
  assign n61 = ~x6 & ~x7 ;
  assign n62 = ~x2 & ~x3 ;
  assign n63 = n61 & n62 ;
  assign n64 = ~n60 & ~n63 ;
  assign n65 = n64 ^ n59 ;
  assign n66 = n59 ^ x5 ;
  assign n67 = n66 ^ n59 ;
  assign n68 = n67 ^ n58 ;
  assign n69 = n65 & ~n68 ;
  assign n70 = n69 ^ n64 ;
  assign n71 = n58 & n70 ;
  assign n72 = ~n56 & ~n71 ;
  assign n73 = x5 ^ x3 ;
  assign n74 = n73 ^ x5 ;
  assign n75 = n33 ^ x5 ;
  assign n76 = n74 & n75 ;
  assign n77 = n76 ^ x5 ;
  assign n78 = n31 & n77 ;
  assign n79 = n72 & ~n78 ;
  assign n80 = n79 ^ x1 ;
  assign n81 = n80 ^ n79 ;
  assign n82 = x0 & ~x2 ;
  assign n83 = n61 & n82 ;
  assign n84 = ~x0 & n31 ;
  assign n85 = n84 ^ x4 ;
  assign n86 = ~n83 & n85 ;
  assign n87 = ~x5 & ~n86 ;
  assign n88 = ~x3 & ~n10 ;
  assign n89 = n88 ^ x0 ;
  assign n90 = n89 ^ n44 ;
  assign n91 = ~x7 & ~n27 ;
  assign n92 = n91 ^ x2 ;
  assign n93 = ~x0 & n92 ;
  assign n94 = n93 ^ x2 ;
  assign n95 = ~n90 & n94 ;
  assign n96 = n95 ^ n93 ;
  assign n97 = n96 ^ x2 ;
  assign n98 = n97 ^ x0 ;
  assign n99 = ~n44 & ~n98 ;
  assign n100 = ~x4 & ~n99 ;
  assign n101 = x6 ^ x0 ;
  assign n102 = n101 ^ x2 ;
  assign n103 = n102 ^ x0 ;
  assign n104 = x2 ^ x0 ;
  assign n105 = n102 & ~n104 ;
  assign n106 = n105 ^ n103 ;
  assign n107 = n48 & n106 ;
  assign n108 = n107 ^ n105 ;
  assign n109 = n103 & n108 ;
  assign n110 = n109 ^ n105 ;
  assign n111 = n43 & n110 ;
  assign n112 = ~n10 & ~n27 ;
  assign n113 = ~x4 & x7 ;
  assign n114 = n33 & ~n113 ;
  assign n115 = ~n112 & n114 ;
  assign n116 = ~n111 & ~n115 ;
  assign n117 = ~n100 & n116 ;
  assign n118 = ~n87 & n117 ;
  assign n119 = n118 ^ n79 ;
  assign n120 = n81 & n119 ;
  assign n121 = n120 ^ n79 ;
  assign n122 = ~n42 & n121 ;
  assign y0 = ~n122 ;
endmodule
