module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 ;
  assign n20 = ~x16 & ~x17 ;
  assign n21 = x14 & ~n20 ;
  assign n22 = x7 & x17 ;
  assign n23 = x8 & ~n22 ;
  assign n24 = n21 & ~n23 ;
  assign n25 = x4 & n23 ;
  assign n26 = ~n20 & ~n25 ;
  assign n27 = x16 & x17 ;
  assign n28 = x6 & n27 ;
  assign n29 = n28 ^ x16 ;
  assign n30 = n29 ^ x6 ;
  assign n31 = n30 ^ n26 ;
  assign n32 = ~x16 & x17 ;
  assign n33 = n32 ^ x7 ;
  assign n34 = ~n29 & n33 ;
  assign n35 = n34 ^ x7 ;
  assign n36 = ~n31 & n35 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = n37 ^ x7 ;
  assign n39 = n38 ^ n29 ;
  assign n40 = ~n26 & ~n39 ;
  assign n41 = ~x3 & ~n40 ;
  assign n42 = ~x11 & ~x12 ;
  assign n43 = x1 & ~n42 ;
  assign n44 = ~x13 & n43 ;
  assign n45 = n20 & ~n44 ;
  assign n46 = ~x14 & ~n45 ;
  assign n47 = ~n41 & n46 ;
  assign n51 = x4 & ~x9 ;
  assign n55 = ~x8 & x16 ;
  assign n56 = ~x7 & ~x17 ;
  assign n57 = ~n22 & ~n56 ;
  assign n58 = n55 & ~n57 ;
  assign n59 = n51 & n58 ;
  assign n48 = ~x7 & x16 ;
  assign n49 = x14 & n48 ;
  assign n50 = x7 & ~x8 ;
  assign n52 = n32 & n51 ;
  assign n53 = n50 & n52 ;
  assign n54 = ~n49 & ~n53 ;
  assign n60 = n59 ^ n54 ;
  assign n61 = n60 ^ n54 ;
  assign n62 = n21 & ~n27 ;
  assign n63 = n62 ^ n54 ;
  assign n64 = n63 ^ n54 ;
  assign n65 = ~n61 & ~n64 ;
  assign n66 = n65 ^ n54 ;
  assign n67 = x6 & n66 ;
  assign n68 = n67 ^ n54 ;
  assign n69 = ~n47 & n68 ;
  assign n70 = ~n24 & n69 ;
  assign n71 = n70 ^ x14 ;
  assign n72 = n71 ^ n70 ;
  assign n74 = ~x2 & ~x10 ;
  assign n75 = x6 & ~x9 ;
  assign n76 = n55 & ~n75 ;
  assign n77 = n74 & ~n76 ;
  assign n73 = x17 ^ x16 ;
  assign n78 = n77 ^ n73 ;
  assign n79 = n77 ^ x17 ;
  assign n80 = n79 ^ x17 ;
  assign n81 = n80 ^ n78 ;
  assign n82 = n48 ^ x6 ;
  assign n83 = ~n48 & ~n82 ;
  assign n84 = n83 ^ x17 ;
  assign n85 = n84 ^ n48 ;
  assign n86 = ~n81 & n85 ;
  assign n87 = n86 ^ n83 ;
  assign n88 = n87 ^ n48 ;
  assign n89 = ~n78 & ~n88 ;
  assign n90 = n89 ^ n77 ;
  assign n91 = n29 ^ x17 ;
  assign n92 = n29 ^ x8 ;
  assign n93 = x8 ^ x7 ;
  assign n94 = n93 ^ n29 ;
  assign n95 = n29 & n94 ;
  assign n96 = n95 ^ n29 ;
  assign n97 = ~n92 & n96 ;
  assign n98 = n97 ^ n95 ;
  assign n99 = n98 ^ n29 ;
  assign n100 = n99 ^ n93 ;
  assign n101 = n91 & n100 ;
  assign n102 = n101 ^ x17 ;
  assign n103 = n90 & ~n102 ;
  assign n104 = n103 ^ n70 ;
  assign n105 = n104 ^ n70 ;
  assign n106 = ~n72 & ~n105 ;
  assign n107 = n106 ^ n70 ;
  assign n108 = x15 & ~n107 ;
  assign n109 = n108 ^ n70 ;
  assign n110 = ~x18 & ~n109 ;
  assign n111 = x14 & ~x15 ;
  assign n112 = ~x14 & x15 ;
  assign n113 = n74 & n112 ;
  assign n114 = ~n111 & ~n113 ;
  assign n115 = ~x6 & ~x16 ;
  assign n116 = ~x8 & n115 ;
  assign n117 = x17 ^ x7 ;
  assign n118 = x18 ^ x17 ;
  assign n119 = n118 ^ x18 ;
  assign n120 = ~x9 & ~n111 ;
  assign n121 = n120 ^ x18 ;
  assign n122 = n119 & ~n121 ;
  assign n123 = n122 ^ x18 ;
  assign n124 = ~n117 & n123 ;
  assign n125 = n116 & n124 ;
  assign n126 = ~n114 & n125 ;
  assign n127 = x6 & ~x8 ;
  assign n128 = x18 & n113 ;
  assign n129 = ~x9 & n128 ;
  assign n130 = ~n127 & ~n129 ;
  assign n131 = ~n111 & ~n128 ;
  assign n132 = x16 ^ x6 ;
  assign n133 = ~n131 & ~n132 ;
  assign n134 = ~n130 & n133 ;
  assign n135 = ~n57 & n134 ;
  assign n136 = ~n126 & ~n135 ;
  assign n137 = ~n110 & n136 ;
  assign y0 = ~n137 ;
endmodule
