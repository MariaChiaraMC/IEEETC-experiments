module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 ;
  assign n9 = x3 & x5 ;
  assign n10 = ~x3 & x6 ;
  assign n11 = x7 ^ x5 ;
  assign n12 = n10 & n11 ;
  assign n13 = ~n9 & ~n12 ;
  assign n14 = x1 & ~n13 ;
  assign n15 = ~x4 & n14 ;
  assign n16 = x4 & x5 ;
  assign n17 = n10 & n16 ;
  assign n18 = x1 & n17 ;
  assign n19 = x2 & ~n18 ;
  assign n20 = ~x4 & ~x5 ;
  assign n21 = x3 ^ x1 ;
  assign n22 = n21 ^ x1 ;
  assign n23 = x7 ^ x1 ;
  assign n24 = ~n22 & n23 ;
  assign n25 = n24 ^ x1 ;
  assign n26 = ~x6 & ~n25 ;
  assign n27 = n20 & n26 ;
  assign n28 = n19 & ~n27 ;
  assign n29 = ~n15 & n28 ;
  assign n30 = ~x2 & ~x6 ;
  assign n32 = ~x1 & n20 ;
  assign n33 = ~n16 & ~n32 ;
  assign n31 = x3 & ~x7 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n34 ^ n33 ;
  assign n36 = n35 ^ x2 ;
  assign n37 = x5 & ~x7 ;
  assign n38 = ~x1 & x4 ;
  assign n39 = ~n37 & n38 ;
  assign n40 = n39 ^ n9 ;
  assign n41 = ~n9 & ~n40 ;
  assign n42 = n41 ^ n33 ;
  assign n43 = n42 ^ n9 ;
  assign n44 = n36 & n43 ;
  assign n45 = n44 ^ n41 ;
  assign n46 = n45 ^ n9 ;
  assign n47 = ~x2 & ~n46 ;
  assign n48 = n47 ^ x2 ;
  assign n49 = ~x0 & n48 ;
  assign n50 = ~n30 & n49 ;
  assign n51 = ~n29 & n50 ;
  assign n52 = x0 & n38 ;
  assign n53 = n9 & n30 ;
  assign n54 = n52 & n53 ;
  assign n55 = x7 & n54 ;
  assign n56 = ~n51 & ~n55 ;
  assign y0 = ~n56 ;
endmodule
