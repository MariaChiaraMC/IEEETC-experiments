module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n10 = x0 & ~x1 ;
  assign n11 = ~x3 & ~n10 ;
  assign n12 = x4 ^ x1 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = x5 ^ x0 ;
  assign n15 = x1 & n14 ;
  assign n16 = n15 ^ x5 ;
  assign n17 = n13 & n16 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n18 ^ x5 ;
  assign n20 = n19 ^ x1 ;
  assign n21 = n11 & n20 ;
  assign n22 = x4 ^ x3 ;
  assign n23 = n22 ^ x4 ;
  assign n24 = x6 ^ x4 ;
  assign n25 = n23 & ~n24 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = n10 & ~n26 ;
  assign n28 = ~n21 & ~n27 ;
  assign n8 = ~x0 & ~x1 ;
  assign n9 = x3 & n8 ;
  assign n29 = n28 ^ n9 ;
  assign n30 = x2 & ~n29 ;
  assign n31 = n30 ^ n28 ;
  assign y0 = ~n31 ;
endmodule
