module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 ;
  output y0 ;
  wire n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 ;
  assign n14 = ~x5 & ~x8 ;
  assign n15 = ~x9 & ~x10 ;
  assign n16 = n14 & n15 ;
  assign n17 = ~x11 & x12 ;
  assign n18 = x7 ^ x6 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = x7 ^ x2 ;
  assign n22 = ~x4 & ~n21 ;
  assign n23 = n22 ^ x2 ;
  assign n24 = ~n20 & n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n25 ^ x2 ;
  assign n27 = n26 ^ x4 ;
  assign n28 = n17 & ~n27 ;
  assign n29 = n16 & n28 ;
  assign n30 = n29 ^ x3 ;
  assign n31 = ~x1 & x2 ;
  assign n32 = ~x4 & ~n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = x3 ^ x0 ;
  assign n35 = n34 ^ x3 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = ~n32 & n36 ;
  assign n38 = n37 ^ n32 ;
  assign n39 = ~n33 & ~n38 ;
  assign n40 = n39 ^ n37 ;
  assign n41 = n40 ^ n32 ;
  assign n42 = n41 ^ n35 ;
  assign n43 = n30 & n42 ;
  assign n44 = n43 ^ n34 ;
  assign y0 = n44 ;
endmodule
