module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 ;
  assign n141 = x7 & ~x10 ;
  assign n18 = x8 & x10 ;
  assign n16 = ~x2 & ~x3 ;
  assign n110 = x0 & ~x1 ;
  assign n111 = ~n16 & n110 ;
  assign n112 = x8 & x11 ;
  assign n113 = ~n111 & n112 ;
  assign n114 = ~n18 & ~n113 ;
  assign n13 = x0 & ~x2 ;
  assign n14 = x10 & n13 ;
  assign n15 = x3 & n14 ;
  assign n17 = n16 ^ x8 ;
  assign n19 = x0 & n18 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = ~x0 & ~x2 ;
  assign n24 = x3 & n23 ;
  assign n25 = x0 & x3 ;
  assign n26 = x2 & ~x10 ;
  assign n27 = x4 & n26 ;
  assign n28 = n27 ^ x5 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = n26 ^ n25 ;
  assign n32 = ~x6 & ~n31 ;
  assign n33 = n32 ^ n27 ;
  assign n34 = n30 & n33 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = ~n25 & n35 ;
  assign n37 = n36 ^ n32 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = ~n24 & ~n38 ;
  assign n40 = n39 ^ n20 ;
  assign n41 = n40 ^ n17 ;
  assign n42 = n22 & n41 ;
  assign n43 = n42 ^ n39 ;
  assign n44 = ~x4 & x10 ;
  assign n45 = ~x0 & ~x10 ;
  assign n46 = ~n44 & ~n45 ;
  assign n47 = n39 & n46 ;
  assign n48 = n47 ^ n17 ;
  assign n49 = n43 & n48 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = n17 & n50 ;
  assign n52 = n51 ^ n42 ;
  assign n53 = n52 ^ x8 ;
  assign n54 = n53 ^ n39 ;
  assign n55 = n54 ^ x1 ;
  assign n56 = n55 ^ n54 ;
  assign n57 = ~x6 & ~x8 ;
  assign n58 = x6 & x10 ;
  assign n59 = ~n57 & ~n58 ;
  assign n60 = n24 & ~n59 ;
  assign n61 = n45 & n57 ;
  assign n62 = n18 & n25 ;
  assign n63 = ~n61 & ~n62 ;
  assign n64 = n63 ^ x3 ;
  assign n65 = n64 ^ x2 ;
  assign n84 = n65 ^ n64 ;
  assign n66 = ~x5 & n27 ;
  assign n67 = x0 & n57 ;
  assign n68 = n66 & n67 ;
  assign n69 = x5 & ~x10 ;
  assign n70 = ~x8 & n69 ;
  assign n71 = ~n44 & ~n70 ;
  assign n72 = n13 & ~n71 ;
  assign n73 = x4 & x5 ;
  assign n74 = n19 & n73 ;
  assign n75 = ~n61 & ~n74 ;
  assign n76 = ~n72 & n75 ;
  assign n77 = ~n68 & n76 ;
  assign n78 = n77 ^ n65 ;
  assign n79 = n78 ^ n64 ;
  assign n80 = n65 ^ n63 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n81 ^ n79 ;
  assign n83 = n79 & n82 ;
  assign n85 = n84 ^ n83 ;
  assign n86 = n85 ^ n79 ;
  assign n87 = x4 ^ x0 ;
  assign n88 = n58 ^ x4 ;
  assign n89 = n88 ^ n58 ;
  assign n90 = x6 & n18 ;
  assign n91 = n90 ^ n58 ;
  assign n92 = n89 & ~n91 ;
  assign n93 = n92 ^ n58 ;
  assign n94 = n87 & n93 ;
  assign n95 = n94 ^ x0 ;
  assign n96 = ~n59 & ~n95 ;
  assign n97 = n96 ^ n64 ;
  assign n98 = n83 ^ n79 ;
  assign n99 = ~n97 & n98 ;
  assign n100 = n99 ^ n64 ;
  assign n101 = n86 & n100 ;
  assign n102 = n101 ^ n64 ;
  assign n103 = n102 ^ x3 ;
  assign n104 = n103 ^ n64 ;
  assign n105 = ~n60 & n104 ;
  assign n106 = n105 ^ n54 ;
  assign n107 = ~n56 & n106 ;
  assign n108 = n107 ^ n54 ;
  assign n109 = ~n15 & n108 ;
  assign n115 = n114 ^ n109 ;
  assign n116 = ~x3 & ~n73 ;
  assign n117 = n110 & ~n116 ;
  assign n118 = n13 ^ x1 ;
  assign n119 = n118 ^ n13 ;
  assign n120 = x6 & n23 ;
  assign n121 = n120 ^ n13 ;
  assign n122 = ~n119 & n121 ;
  assign n123 = n122 ^ n13 ;
  assign n124 = ~x4 & n13 ;
  assign n125 = n124 ^ n117 ;
  assign n126 = n123 & ~n125 ;
  assign n127 = n126 ^ n124 ;
  assign n128 = ~n117 & n127 ;
  assign n129 = n128 ^ n117 ;
  assign n130 = x10 & n129 ;
  assign n131 = n130 ^ n109 ;
  assign n132 = n109 ^ x7 ;
  assign n133 = n109 & ~n132 ;
  assign n134 = n133 ^ n109 ;
  assign n135 = ~n131 & n134 ;
  assign n136 = n135 ^ n133 ;
  assign n137 = n136 ^ n109 ;
  assign n138 = n137 ^ x7 ;
  assign n139 = n115 & ~n138 ;
  assign n140 = n139 ^ n114 ;
  assign n142 = n141 ^ n140 ;
  assign n143 = n142 ^ n140 ;
  assign n144 = n140 ^ x8 ;
  assign n145 = n144 ^ n140 ;
  assign n146 = n143 & n145 ;
  assign n147 = n146 ^ n140 ;
  assign n148 = x9 & ~n147 ;
  assign n149 = n148 ^ n140 ;
  assign y0 = ~n149 ;
endmodule
