module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 ;
  assign n31 = x9 ^ x3 ;
  assign n12 = x7 ^ x2 ;
  assign n14 = x7 ^ x1 ;
  assign n13 = x7 ^ x6 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = n15 ^ n12 ;
  assign n22 = n14 ^ x7 ;
  assign n17 = x7 ^ x5 ;
  assign n18 = n17 ^ x7 ;
  assign n19 = x7 ^ x0 ;
  assign n20 = n19 ^ x7 ;
  assign n21 = n18 & n20 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n16 & n23 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ n14 ;
  assign n27 = n26 ^ n22 ;
  assign n28 = n12 & ~n27 ;
  assign n29 = n28 ^ x2 ;
  assign n30 = n29 ^ x9 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = x9 ^ x8 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n32 & n34 ;
  assign n36 = n35 ^ n31 ;
  assign n37 = x10 ^ x4 ;
  assign n38 = n37 ^ x9 ;
  assign n39 = n38 ^ x10 ;
  assign n40 = ~n36 & n39 ;
  assign n41 = n40 ^ n37 ;
  assign y0 = n41 ;
endmodule
