module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 ;
  assign n8 = ~x1 & ~x2 ;
  assign n9 = x0 & ~n8 ;
  assign n10 = x3 ^ x1 ;
  assign n11 = x5 ^ x1 ;
  assign n12 = x5 ^ x2 ;
  assign n13 = n12 ^ x2 ;
  assign n14 = x6 ^ x2 ;
  assign n15 = ~n13 & ~n14 ;
  assign n16 = n15 ^ x2 ;
  assign n17 = n11 & n16 ;
  assign n18 = n17 ^ x1 ;
  assign n19 = ~n10 & ~n18 ;
  assign n20 = n19 ^ x6 ;
  assign n21 = ~x2 & ~x5 ;
  assign n22 = ~x1 & x3 ;
  assign n23 = ~x2 & x3 ;
  assign n24 = ~n22 & ~n23 ;
  assign n25 = ~n21 & ~n24 ;
  assign n26 = n25 ^ n19 ;
  assign n27 = n19 ^ x4 ;
  assign n28 = ~n19 & n27 ;
  assign n29 = n28 ^ n19 ;
  assign n30 = ~n26 & ~n29 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n31 ^ n19 ;
  assign n33 = n32 ^ x4 ;
  assign n34 = n20 & n33 ;
  assign n35 = n34 ^ x6 ;
  assign n36 = ~n9 & ~n35 ;
  assign n37 = n10 ^ x5 ;
  assign n38 = x5 ^ x4 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = n10 ^ x2 ;
  assign n41 = n40 ^ x2 ;
  assign n42 = n23 ^ x2 ;
  assign n43 = ~n41 & ~n42 ;
  assign n44 = n43 ^ x2 ;
  assign n45 = n44 ^ n37 ;
  assign n46 = ~n39 & ~n45 ;
  assign n47 = n46 ^ n43 ;
  assign n48 = n47 ^ x2 ;
  assign n49 = n48 ^ n38 ;
  assign n50 = ~n37 & n49 ;
  assign n51 = n50 ^ n37 ;
  assign n52 = n51 ^ x4 ;
  assign n53 = n36 & n52 ;
  assign y0 = n53 ;
endmodule
