module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n8 = x2 ^ x1 ;
  assign n9 = x5 ^ x4 ;
  assign n10 = x6 ^ x5 ;
  assign n11 = x6 ^ x3 ;
  assign n12 = x6 & ~n11 ;
  assign n13 = n12 ^ x6 ;
  assign n14 = ~n10 & n13 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n15 ^ x6 ;
  assign n17 = n16 ^ x3 ;
  assign n18 = n9 & ~n17 ;
  assign n19 = n18 ^ x3 ;
  assign n20 = n19 ^ x2 ;
  assign n21 = x1 ^ x0 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = ~n19 & ~n22 ;
  assign n24 = n23 ^ n19 ;
  assign n25 = ~n20 & ~n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n26 ^ n19 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = ~n8 & ~n28 ;
  assign y0 = n29 ;
endmodule
