module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 ;
  assign n8 = x5 & x6 ;
  assign n9 = x2 & ~n8 ;
  assign n10 = x0 & ~x4 ;
  assign n11 = ~x5 & ~x6 ;
  assign n12 = x0 & n11 ;
  assign n13 = ~n10 & ~n12 ;
  assign n14 = ~n9 & n13 ;
  assign n15 = x1 & ~n14 ;
  assign n16 = ~x0 & x2 ;
  assign n17 = x4 & ~n16 ;
  assign n18 = x2 & n11 ;
  assign n19 = ~n16 & ~n18 ;
  assign n20 = ~n17 & ~n19 ;
  assign n21 = ~n15 & ~n20 ;
  assign n22 = ~x3 & ~n21 ;
  assign n23 = ~x2 & x3 ;
  assign n24 = x4 ^ x0 ;
  assign n25 = n8 ^ x4 ;
  assign n26 = ~n24 & n25 ;
  assign n27 = n26 ^ x4 ;
  assign n28 = n23 & n27 ;
  assign n29 = x1 & ~n28 ;
  assign n30 = n17 ^ x3 ;
  assign n31 = n17 ^ x5 ;
  assign n32 = x3 ^ x2 ;
  assign n33 = n32 ^ n17 ;
  assign n34 = n17 & ~n33 ;
  assign n35 = n34 ^ n17 ;
  assign n36 = ~n31 & n35 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = n37 ^ n17 ;
  assign n39 = n38 ^ n32 ;
  assign n40 = n30 & ~n39 ;
  assign n41 = n40 ^ x3 ;
  assign n42 = ~n29 & n41 ;
  assign n43 = x1 & x6 ;
  assign n44 = ~x4 & ~x5 ;
  assign n45 = ~n43 & n44 ;
  assign n46 = n16 & n45 ;
  assign n47 = ~n42 & ~n46 ;
  assign n48 = ~n22 & n47 ;
  assign y0 = n48 ;
endmodule
