module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 ;
  assign n15 = x3 & x4 ;
  assign n16 = ~x0 & n15 ;
  assign n17 = x1 & x6 ;
  assign n20 = n17 ^ x2 ;
  assign n21 = n20 ^ n17 ;
  assign n18 = n17 ^ x9 ;
  assign n19 = n18 ^ n17 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = ~x11 & ~x12 ;
  assign n24 = x7 & n17 ;
  assign n25 = ~x8 & ~x10 ;
  assign n26 = ~x13 & n25 ;
  assign n27 = n24 & n26 ;
  assign n28 = n23 & n27 ;
  assign n29 = n28 ^ n17 ;
  assign n30 = n29 ^ n17 ;
  assign n31 = n30 ^ n21 ;
  assign n32 = n21 & n31 ;
  assign n33 = n32 ^ n21 ;
  assign n34 = n22 & n33 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = n35 ^ n17 ;
  assign n37 = n36 ^ n21 ;
  assign n38 = x5 & ~n37 ;
  assign n39 = n38 ^ n17 ;
  assign n40 = n16 & ~n39 ;
  assign y0 = n40 ;
endmodule
