module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 ;
  assign n18 = x16 ^ x14 ;
  assign n19 = n18 ^ x16 ;
  assign n20 = n19 ^ x12 ;
  assign n21 = ~x9 & ~x10 ;
  assign n22 = ~x7 & ~x8 ;
  assign n23 = ~x4 & ~x5 ;
  assign n24 = n22 & ~n23 ;
  assign n25 = n21 & n24 ;
  assign n26 = ~x2 & ~x11 ;
  assign n27 = ~n25 & n26 ;
  assign n28 = x13 & ~n27 ;
  assign n29 = ~x15 & n28 ;
  assign n30 = x7 ^ x1 ;
  assign n31 = n30 ^ x1 ;
  assign n32 = n31 ^ x11 ;
  assign n33 = ~x2 & ~x8 ;
  assign n34 = n33 ^ x11 ;
  assign n35 = ~n21 & ~n34 ;
  assign n36 = n35 ^ x1 ;
  assign n37 = ~n32 & n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = ~x11 & n38 ;
  assign n40 = n39 ^ n35 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n41 ^ x11 ;
  assign n43 = n29 & ~n42 ;
  assign n44 = n43 ^ x16 ;
  assign n60 = n44 ^ x16 ;
  assign n45 = x13 ^ x11 ;
  assign n46 = x13 ^ x6 ;
  assign n47 = x13 ^ x3 ;
  assign n48 = ~x13 & ~n47 ;
  assign n49 = n48 ^ x13 ;
  assign n50 = n46 & ~n49 ;
  assign n51 = n50 ^ n48 ;
  assign n52 = n51 ^ x13 ;
  assign n53 = n52 ^ x3 ;
  assign n54 = n45 & ~n53 ;
  assign n55 = n54 ^ x16 ;
  assign n56 = n55 ^ n44 ;
  assign n57 = n44 ^ x0 ;
  assign n58 = n57 ^ n44 ;
  assign n59 = n56 & n58 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = n20 & n61 ;
  assign n63 = n62 ^ n59 ;
  assign n64 = n63 ^ x16 ;
  assign n65 = n64 ^ n60 ;
  assign n66 = ~x12 & ~n65 ;
  assign n67 = n66 ^ x16 ;
  assign y0 = ~n67 ;
endmodule
