module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n10 = ~x5 & ~x7 ;
  assign n11 = ~x1 & ~n10 ;
  assign n12 = ~x2 & x4 ;
  assign n13 = ~x8 & ~n12 ;
  assign n14 = ~n11 & n13 ;
  assign n15 = ~x0 & ~x6 ;
  assign n16 = ~x3 & n15 ;
  assign n17 = x2 ^ x1 ;
  assign n18 = n17 ^ x2 ;
  assign n19 = x7 ^ x2 ;
  assign n20 = n18 & ~n19 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = x2 & ~x4 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = n21 & n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n16 & n25 ;
  assign n27 = n26 ^ n16 ;
  assign n28 = n14 & n27 ;
  assign y0 = n28 ;
endmodule
