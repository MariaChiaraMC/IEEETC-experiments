module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 ;
  assign n16 = x12 ^ x11 ;
  assign n17 = ~x1 & ~x8 ;
  assign n18 = ~x0 & ~x13 ;
  assign n19 = x9 & n18 ;
  assign n20 = x11 & n19 ;
  assign n21 = ~n17 & n20 ;
  assign n22 = x10 & ~n21 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = n23 ^ x12 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = ~x2 & ~x3 ;
  assign n27 = x4 & n26 ;
  assign n28 = ~x10 & ~n27 ;
  assign n29 = x2 & x3 ;
  assign n30 = x13 ^ x5 ;
  assign n31 = ~x0 & ~n30 ;
  assign n32 = n31 ^ x5 ;
  assign n33 = ~n29 & n32 ;
  assign n34 = ~x9 & ~n33 ;
  assign n35 = n28 & n34 ;
  assign n36 = n35 ^ x0 ;
  assign n38 = ~x3 & ~x7 ;
  assign n39 = x6 & ~n38 ;
  assign n37 = x3 ^ x2 ;
  assign n40 = n39 ^ n37 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n37 ^ x3 ;
  assign n43 = n41 & n42 ;
  assign n44 = n43 ^ n37 ;
  assign n45 = ~x5 & ~n37 ;
  assign n46 = n45 ^ x4 ;
  assign n47 = ~n44 & n46 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = x4 & n48 ;
  assign n50 = n49 ^ n37 ;
  assign n51 = n50 ^ x4 ;
  assign n52 = ~x13 & n51 ;
  assign n53 = n52 ^ n35 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = ~x9 & ~x14 ;
  assign n56 = ~x12 & ~n55 ;
  assign n57 = ~x13 & ~n56 ;
  assign n58 = x10 & ~n57 ;
  assign n59 = n58 ^ n52 ;
  assign n60 = ~n54 & ~n59 ;
  assign n61 = n60 ^ n52 ;
  assign n62 = ~n36 & n61 ;
  assign n63 = n62 ^ x0 ;
  assign n64 = x1 & ~n63 ;
  assign n65 = n64 ^ n23 ;
  assign n66 = n65 ^ n16 ;
  assign n67 = n25 & n66 ;
  assign n68 = n67 ^ n64 ;
  assign n69 = ~x13 & ~n64 ;
  assign n70 = n69 ^ n16 ;
  assign n71 = ~n68 & n70 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = n16 & n72 ;
  assign n74 = n73 ^ n67 ;
  assign n75 = n74 ^ x11 ;
  assign n76 = n75 ^ n64 ;
  assign y0 = n76 ;
endmodule
