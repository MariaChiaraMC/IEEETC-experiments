module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 ;
  assign n7 = ~x0 & x1 ;
  assign n8 = x3 ^ x2 ;
  assign n9 = n8 ^ x2 ;
  assign n10 = n9 ^ n7 ;
  assign n11 = x5 ^ x2 ;
  assign n12 = x4 ^ x2 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n11 & n13 ;
  assign n15 = n14 ^ x2 ;
  assign n16 = n15 ^ n11 ;
  assign n17 = n10 & n16 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = n18 ^ n11 ;
  assign n20 = n7 & n19 ;
  assign y0 = n20 ;
endmodule
