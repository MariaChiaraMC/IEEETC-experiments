module top( x0 , x1 , x2 , x3 , x4 , y0 );
  input x0 , x1 , x2 , x3 , x4 ;
  output y0 ;
  wire n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 ;
  assign n6 = x4 ^ x3 ;
  assign n14 = n6 ^ x4 ;
  assign n7 = n6 ^ x1 ;
  assign n8 = n7 ^ n6 ;
  assign n9 = n8 ^ x4 ;
  assign n10 = n6 ^ x0 ;
  assign n11 = n10 ^ n7 ;
  assign n12 = n11 ^ n9 ;
  assign n13 = n9 & ~n12 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = n15 ^ n9 ;
  assign n17 = x3 ^ x2 ;
  assign n18 = n17 ^ x4 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = n19 ^ x4 ;
  assign n21 = n13 ^ n9 ;
  assign n22 = n20 & n21 ;
  assign n23 = n22 ^ x4 ;
  assign n24 = ~n16 & ~n23 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = n25 ^ n18 ;
  assign n27 = n26 ^ x4 ;
  assign y0 = n27 ;
endmodule
