// Benchmark "./pla/b11.pla_res_5NonExact" written by ABC on Fri Nov 20 10:19:57 2020

module \./pla/b11.pla_res_5NonExact  ( 
    x0, x1,
    z0  );
  input  x0, x1;
  output z0;
  assign z0 = ~x0 & ~x1;
endmodule


