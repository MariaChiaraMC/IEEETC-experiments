module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n8 = x0 & x1 ;
  assign n9 = ~x0 & ~x1 ;
  assign n10 = ~x4 & x5 ;
  assign n11 = ~x2 & ~n10 ;
  assign n12 = n9 & ~n11 ;
  assign n13 = ~n8 & ~n12 ;
  assign n14 = x3 & ~n13 ;
  assign n15 = x1 ^ x0 ;
  assign n16 = x3 ^ x1 ;
  assign n17 = n16 ^ x3 ;
  assign n18 = x5 ^ x3 ;
  assign n19 = n17 & ~n18 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = ~n15 & ~n20 ;
  assign n22 = x4 & n21 ;
  assign n23 = x0 & x6 ;
  assign n24 = x3 & ~n23 ;
  assign n25 = ~n9 & ~n24 ;
  assign n26 = ~x2 & n25 ;
  assign n27 = ~n22 & ~n26 ;
  assign n28 = ~n14 & n27 ;
  assign y0 = ~n28 ;
endmodule
