module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n16 = x9 & ~x14 ;
  assign n17 = n16 ^ x10 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = ~x0 & x6 ;
  assign n20 = ~x3 & x7 ;
  assign n21 = x4 & n20 ;
  assign n22 = n19 & ~n21 ;
  assign n23 = ~x2 & ~x9 ;
  assign n24 = ~x1 & n23 ;
  assign n25 = n22 & n24 ;
  assign n26 = n25 ^ n16 ;
  assign n27 = ~n18 & ~n26 ;
  assign n28 = n27 ^ n16 ;
  assign n29 = ~x13 & ~n28 ;
  assign n30 = n29 ^ x10 ;
  assign y0 = n30 ;
endmodule
