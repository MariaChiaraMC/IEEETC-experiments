module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n8 = ~x0 & x3 ;
  assign n9 = x2 & x5 ;
  assign n10 = ~n8 & ~n9 ;
  assign n7 = x2 & x4 ;
  assign n11 = n10 ^ n7 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = x0 & ~x5 ;
  assign n14 = n13 ^ n10 ;
  assign n15 = n14 ^ n10 ;
  assign n16 = ~n12 & ~n15 ;
  assign n17 = n16 ^ n10 ;
  assign n18 = ~x1 & ~n17 ;
  assign n19 = n18 ^ n10 ;
  assign n20 = ~x1 & ~n7 ;
  assign n21 = ~x2 & ~x4 ;
  assign n22 = x0 & ~n21 ;
  assign n23 = ~n20 & n22 ;
  assign n24 = ~x1 & x3 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = ~x3 & n7 ;
  assign n28 = ~n21 & ~n27 ;
  assign n29 = n28 ^ n24 ;
  assign n30 = ~n26 & ~n29 ;
  assign n31 = n30 ^ n24 ;
  assign n32 = ~x4 & n24 ;
  assign n33 = n32 ^ n23 ;
  assign n34 = n31 & ~n33 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = ~n23 & n35 ;
  assign n37 = n36 ^ n23 ;
  assign n38 = n19 & ~n37 ;
  assign y0 = ~n38 ;
endmodule
