module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 ;
  assign n9 = x2 & x7 ;
  assign n10 = ~x0 & n9 ;
  assign n11 = x4 & ~x7 ;
  assign n12 = ~n10 & ~n11 ;
  assign n13 = x1 & ~n12 ;
  assign n14 = ~x0 & ~x1 ;
  assign n15 = n14 ^ x3 ;
  assign n20 = n15 ^ x5 ;
  assign n21 = n20 ^ n14 ;
  assign n16 = x7 ^ x2 ;
  assign n17 = n16 ^ x7 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n18 ^ n14 ;
  assign n22 = n21 ^ n19 ;
  assign n25 = n15 ^ n14 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = n21 & ~n26 ;
  assign n23 = n15 & n16 ;
  assign n30 = n27 ^ n23 ;
  assign n24 = n23 ^ n22 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = n24 & n28 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n22 & n31 ;
  assign n33 = n32 ^ n27 ;
  assign n34 = n33 ^ n29 ;
  assign n35 = n34 ^ x3 ;
  assign n36 = ~n13 & ~n35 ;
  assign y0 = ~n36 ;
endmodule
