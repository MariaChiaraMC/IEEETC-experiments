module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 ;
  output y0 ;
  wire n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 ;
  assign n28 = x1 & x2 ;
  assign n19 = x13 & x14 ;
  assign n20 = x15 ^ x5 ;
  assign n21 = n20 ^ x15 ;
  assign n22 = ~x3 & ~x12 ;
  assign n23 = n22 ^ x15 ;
  assign n24 = n21 & n23 ;
  assign n25 = n24 ^ x15 ;
  assign n26 = x16 & ~n25 ;
  assign n27 = n19 & ~n26 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = x12 & x14 ;
  assign n34 = x3 & ~x13 ;
  assign n35 = n33 & ~n34 ;
  assign n36 = x5 & x15 ;
  assign n37 = ~n35 & n36 ;
  assign n38 = n37 ^ n30 ;
  assign n39 = n38 ^ n29 ;
  assign n40 = n32 & n39 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = x3 & x12 ;
  assign n43 = ~n22 & ~n42 ;
  assign n44 = ~n37 & n43 ;
  assign n45 = n44 ^ n29 ;
  assign n46 = ~n41 & ~n45 ;
  assign n47 = n46 ^ n44 ;
  assign n48 = ~n29 & n47 ;
  assign n49 = n48 ^ n40 ;
  assign n50 = n49 ^ n28 ;
  assign n51 = n50 ^ n37 ;
  assign n52 = x4 & ~n51 ;
  assign n63 = ~x1 & ~x2 ;
  assign n53 = x2 & x12 ;
  assign n54 = x2 ^ x1 ;
  assign n55 = n54 ^ x2 ;
  assign n56 = x10 & x12 ;
  assign n57 = n56 ^ x2 ;
  assign n58 = n55 & n57 ;
  assign n59 = n58 ^ x2 ;
  assign n60 = x9 & n59 ;
  assign n61 = ~n53 & n60 ;
  assign n62 = ~x5 & ~n61 ;
  assign n64 = n63 ^ n62 ;
  assign n65 = n64 ^ x0 ;
  assign n73 = n65 ^ n64 ;
  assign n66 = ~x8 & n42 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = n67 ^ n64 ;
  assign n69 = n65 ^ n62 ;
  assign n70 = n69 ^ n66 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = n68 & ~n71 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = n74 ^ n68 ;
  assign n76 = n64 ^ n22 ;
  assign n77 = n72 ^ n68 ;
  assign n78 = n76 & n77 ;
  assign n79 = n78 ^ n64 ;
  assign n80 = ~n75 & ~n79 ;
  assign n81 = n80 ^ n64 ;
  assign n82 = n81 ^ n63 ;
  assign n83 = n82 ^ n64 ;
  assign n84 = n52 & n83 ;
  assign n85 = ~x16 & x17 ;
  assign n86 = n19 & n85 ;
  assign n87 = ~n43 & n86 ;
  assign n88 = x6 ^ x3 ;
  assign n89 = n88 ^ x6 ;
  assign n90 = x7 ^ x6 ;
  assign n91 = n89 & n90 ;
  assign n92 = n91 ^ x6 ;
  assign n93 = x15 & n92 ;
  assign n94 = ~n87 & ~n93 ;
  assign n95 = ~x0 & x5 ;
  assign n96 = ~n94 & n95 ;
  assign n97 = n28 & n96 ;
  assign n98 = ~n84 & ~n97 ;
  assign n99 = x11 & ~n98 ;
  assign y0 = n99 ;
endmodule
