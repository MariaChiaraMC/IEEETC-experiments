module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 ;
  output y0 ;
  wire n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 ;
  assign n34 = ~x6 & ~x29 ;
  assign n35 = ~x8 & n34 ;
  assign n36 = ~x7 & n35 ;
  assign n37 = ~x9 & n36 ;
  assign n38 = x12 ^ x0 ;
  assign n39 = ~x2 & ~x3 ;
  assign n40 = ~x1 & n39 ;
  assign n41 = ~x10 & x11 ;
  assign n42 = x15 & x17 ;
  assign n43 = x16 & n42 ;
  assign n44 = ~x13 & n43 ;
  assign n45 = ~x16 & ~x17 ;
  assign n46 = x13 & ~x15 ;
  assign n47 = n45 & n46 ;
  assign n48 = ~n44 & ~n47 ;
  assign n49 = x4 ^ x0 ;
  assign n50 = x5 & ~n49 ;
  assign n51 = n50 ^ x0 ;
  assign n52 = x14 & n51 ;
  assign n53 = ~n48 & n52 ;
  assign n54 = ~x16 & x17 ;
  assign n55 = ~x4 & ~x14 ;
  assign n56 = x0 & ~x5 ;
  assign n57 = n55 & n56 ;
  assign n58 = n54 & n57 ;
  assign n59 = n46 & n58 ;
  assign n60 = ~n53 & ~n59 ;
  assign n61 = n41 & ~n60 ;
  assign n62 = x10 & ~x11 ;
  assign n63 = ~x13 & x15 ;
  assign n64 = n45 & n63 ;
  assign n65 = n57 & n64 ;
  assign n66 = n62 & n65 ;
  assign n67 = ~n61 & ~n66 ;
  assign n68 = n40 & ~n67 ;
  assign n69 = n68 ^ n38 ;
  assign n70 = n69 ^ x12 ;
  assign n71 = n70 ^ n69 ;
  assign n72 = ~x4 & n39 ;
  assign n73 = ~x5 & n72 ;
  assign n74 = ~x1 & x32 ;
  assign n75 = n73 & n74 ;
  assign n76 = ~x14 & x15 ;
  assign n77 = n41 & n76 ;
  assign n78 = n62 ^ x12 ;
  assign n79 = ~x14 & ~x15 ;
  assign n80 = x16 & n79 ;
  assign n81 = x11 & n80 ;
  assign n82 = n81 ^ n62 ;
  assign n83 = n82 ^ n81 ;
  assign n84 = n83 ^ n78 ;
  assign n85 = n42 ^ x16 ;
  assign n86 = n85 ^ x14 ;
  assign n87 = ~x14 & ~n86 ;
  assign n88 = n87 ^ n81 ;
  assign n89 = n88 ^ x14 ;
  assign n90 = n84 & n89 ;
  assign n91 = n90 ^ n87 ;
  assign n92 = n91 ^ x14 ;
  assign n93 = n78 & ~n92 ;
  assign n94 = n93 ^ x12 ;
  assign n95 = ~n77 & ~n94 ;
  assign n96 = x13 & ~n95 ;
  assign n97 = x16 & ~x17 ;
  assign n98 = ~x13 & x14 ;
  assign n99 = ~x10 & n98 ;
  assign n100 = ~n97 & n99 ;
  assign n101 = ~x12 & ~n100 ;
  assign n102 = x11 & n45 ;
  assign n103 = n98 & n102 ;
  assign n104 = ~x15 & n103 ;
  assign n105 = ~n41 & ~n104 ;
  assign n106 = ~n101 & ~n105 ;
  assign n107 = ~n96 & ~n106 ;
  assign n108 = n75 & ~n107 ;
  assign n109 = n108 ^ n69 ;
  assign n110 = n109 ^ n38 ;
  assign n111 = ~n71 & ~n110 ;
  assign n112 = n111 ^ n108 ;
  assign n113 = ~x18 & x19 ;
  assign n114 = n76 & n113 ;
  assign n115 = ~n98 & ~n114 ;
  assign n116 = x16 & x32 ;
  assign n117 = ~x5 & ~x17 ;
  assign n118 = ~x4 & n117 ;
  assign n119 = n116 & n118 ;
  assign n120 = ~n115 & n119 ;
  assign n121 = ~x4 & ~x5 ;
  assign n122 = x30 & x31 ;
  assign n123 = n122 ^ x16 ;
  assign n124 = ~x17 & n123 ;
  assign n125 = n124 ^ x16 ;
  assign n126 = x32 & ~n125 ;
  assign n127 = n121 & n126 ;
  assign n128 = x14 & ~n127 ;
  assign n129 = x18 & ~x19 ;
  assign n130 = x20 & x21 ;
  assign n131 = n113 & ~n130 ;
  assign n132 = ~x22 & n131 ;
  assign n133 = ~n129 & ~n132 ;
  assign n134 = x24 & n97 ;
  assign n135 = ~n133 & n134 ;
  assign n136 = n135 ^ x4 ;
  assign n137 = n136 ^ n135 ;
  assign n138 = n137 ^ n63 ;
  assign n139 = n129 ^ x5 ;
  assign n140 = n129 ^ n116 ;
  assign n141 = n140 ^ n116 ;
  assign n142 = x24 & n113 ;
  assign n143 = n142 ^ x22 ;
  assign n144 = n142 ^ n131 ;
  assign n145 = n144 ^ n131 ;
  assign n146 = x23 & n130 ;
  assign n147 = n146 ^ n131 ;
  assign n148 = n145 & n147 ;
  assign n149 = n148 ^ n131 ;
  assign n150 = ~n143 & ~n149 ;
  assign n151 = n150 ^ x22 ;
  assign n152 = x16 & n151 ;
  assign n153 = n152 ^ n116 ;
  assign n154 = ~n141 & n153 ;
  assign n155 = n154 ^ n116 ;
  assign n156 = n139 & n155 ;
  assign n157 = n156 ^ x5 ;
  assign n158 = ~x17 & n157 ;
  assign n159 = n158 ^ x14 ;
  assign n160 = ~n158 & n159 ;
  assign n161 = n160 ^ n135 ;
  assign n162 = n161 ^ n158 ;
  assign n163 = ~n138 & n162 ;
  assign n164 = n163 ^ n160 ;
  assign n165 = n164 ^ n158 ;
  assign n166 = n63 & ~n165 ;
  assign n167 = n166 ^ n63 ;
  assign n168 = ~n128 & n167 ;
  assign n169 = ~n120 & ~n168 ;
  assign n170 = n40 & ~n169 ;
  assign n171 = n62 & n170 ;
  assign n172 = x5 & n72 ;
  assign n173 = n64 & n172 ;
  assign n174 = ~x1 & n173 ;
  assign n175 = n44 ^ x1 ;
  assign n176 = n72 ^ n44 ;
  assign n177 = n176 ^ n72 ;
  assign n178 = n72 ^ n47 ;
  assign n179 = ~n177 & n178 ;
  assign n180 = n179 ^ n72 ;
  assign n181 = n175 & ~n180 ;
  assign n182 = n181 ^ x1 ;
  assign n183 = ~n174 & ~n182 ;
  assign n184 = x14 & ~n183 ;
  assign n185 = n73 ^ x1 ;
  assign n186 = x32 ^ x1 ;
  assign n187 = x1 & ~x14 ;
  assign n188 = ~n172 & ~n187 ;
  assign n189 = x17 & ~n188 ;
  assign n190 = n189 ^ x1 ;
  assign n191 = ~x1 & n190 ;
  assign n192 = n191 ^ x1 ;
  assign n193 = ~n186 & ~n192 ;
  assign n194 = n193 ^ n191 ;
  assign n195 = n194 ^ x1 ;
  assign n196 = n195 ^ n189 ;
  assign n197 = n185 & n196 ;
  assign n198 = n46 & ~n197 ;
  assign n199 = ~x16 & n198 ;
  assign n200 = ~n184 & ~n199 ;
  assign n201 = n200 ^ x10 ;
  assign n202 = n201 ^ n200 ;
  assign n203 = n202 ^ x11 ;
  assign n204 = x27 & x28 ;
  assign n205 = n204 ^ x26 ;
  assign n206 = x25 & ~n205 ;
  assign n207 = n206 ^ x26 ;
  assign n208 = n207 ^ n75 ;
  assign n209 = n75 & ~n208 ;
  assign n210 = n209 ^ n200 ;
  assign n211 = n210 ^ n75 ;
  assign n212 = n203 & ~n211 ;
  assign n213 = n212 ^ n209 ;
  assign n214 = n213 ^ n75 ;
  assign n215 = x11 & n214 ;
  assign n216 = ~n171 & ~n215 ;
  assign n217 = ~n108 & n216 ;
  assign n218 = n217 ^ n38 ;
  assign n219 = ~n112 & ~n218 ;
  assign n220 = n219 ^ n217 ;
  assign n221 = ~n38 & n220 ;
  assign n222 = n221 ^ n111 ;
  assign n223 = n222 ^ x0 ;
  assign n224 = n223 ^ n108 ;
  assign n225 = n37 & n224 ;
  assign y0 = n225 ;
endmodule
