module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 ;
  assign n9 = x2 & x7 ;
  assign n10 = x4 & n9 ;
  assign n11 = x0 & x1 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = ~x3 & ~x6 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = n13 ^ x6 ;
  assign n17 = n15 & n16 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = n18 ^ n10 ;
  assign n20 = n12 & n19 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n21 ^ n13 ;
  assign n23 = n22 ^ n11 ;
  assign n24 = n10 & n23 ;
  assign n25 = n24 ^ n10 ;
  assign y0 = n25 ;
endmodule
