module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 ;
  output y0 ;
  wire n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 ;
  assign n19 = x13 & ~x17 ;
  assign n20 = x12 & n19 ;
  assign n21 = x15 ^ x13 ;
  assign n22 = ~x8 & ~x10 ;
  assign n23 = ~x7 & ~x9 ;
  assign n24 = ~x4 & ~x5 ;
  assign n25 = n23 & ~n24 ;
  assign n26 = n22 & n25 ;
  assign n27 = ~x2 & ~x11 ;
  assign n28 = ~n26 & n27 ;
  assign n29 = x14 & ~n28 ;
  assign n30 = ~x16 & n29 ;
  assign n31 = x7 ^ x1 ;
  assign n32 = n31 ^ x1 ;
  assign n33 = n32 ^ x11 ;
  assign n34 = ~x2 & ~x9 ;
  assign n35 = n34 ^ x11 ;
  assign n36 = ~n22 & ~n35 ;
  assign n37 = n36 ^ x1 ;
  assign n38 = ~n33 & n37 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = ~x11 & n39 ;
  assign n41 = n40 ^ n36 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = n42 ^ x11 ;
  assign n44 = n30 & ~n43 ;
  assign n45 = n44 ^ x0 ;
  assign n46 = n45 ^ n44 ;
  assign n47 = x14 ^ x11 ;
  assign n48 = x14 ^ x6 ;
  assign n49 = x14 ^ x3 ;
  assign n50 = ~x14 & ~n49 ;
  assign n51 = n50 ^ x14 ;
  assign n52 = n48 & ~n51 ;
  assign n53 = n52 ^ n50 ;
  assign n54 = n53 ^ x14 ;
  assign n55 = n54 ^ x3 ;
  assign n56 = n47 & ~n55 ;
  assign n57 = n56 ^ n44 ;
  assign n58 = n46 & n57 ;
  assign n59 = n58 ^ n44 ;
  assign n60 = n59 ^ x15 ;
  assign n61 = n21 & ~n60 ;
  assign n62 = n61 ^ n58 ;
  assign n63 = n62 ^ n44 ;
  assign n64 = n63 ^ x13 ;
  assign n65 = ~x15 & ~n64 ;
  assign n66 = n65 ^ x15 ;
  assign n67 = ~n20 & n66 ;
  assign y0 = ~n67 ;
endmodule
