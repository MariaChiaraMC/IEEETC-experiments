module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ;
  assign n7 = ~x2 & ~x3 ;
  assign n8 = ~x5 & ~n7 ;
  assign n9 = ~x0 & ~n8 ;
  assign n11 = x4 ^ x0 ;
  assign n14 = n11 ^ x4 ;
  assign n15 = n14 ^ n11 ;
  assign n10 = x4 ^ x2 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = n12 ^ n10 ;
  assign n16 = n15 ^ n13 ;
  assign n20 = n10 ^ x5 ;
  assign n18 = n14 ^ x1 ;
  assign n17 = n10 ^ x3 ;
  assign n19 = n18 ^ n17 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = ~n12 & ~n21 ;
  assign n23 = n22 ^ n17 ;
  assign n24 = n23 ^ n19 ;
  assign n25 = n24 ^ n12 ;
  assign n26 = n25 ^ n20 ;
  assign n27 = n16 & ~n26 ;
  assign n28 = n27 ^ n12 ;
  assign n29 = n28 ^ n13 ;
  assign n30 = n25 ^ n13 ;
  assign n31 = ~n13 & ~n30 ;
  assign n32 = n31 ^ n12 ;
  assign n33 = n29 & ~n32 ;
  assign n34 = n33 ^ n17 ;
  assign n35 = n34 ^ n12 ;
  assign n36 = n35 ^ n13 ;
  assign n37 = n36 ^ x4 ;
  assign n38 = n37 ^ n17 ;
  assign n39 = ~n9 & ~n38 ;
  assign y0 = n39 ;
endmodule
