module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 ;
  assign n13 = ~x1 & x3 ;
  assign n14 = x5 & n13 ;
  assign n15 = x0 & ~n14 ;
  assign n16 = ~x4 & ~n15 ;
  assign n17 = ~x2 & ~n16 ;
  assign n18 = x7 & x10 ;
  assign n19 = x8 & x11 ;
  assign n20 = x6 & n19 ;
  assign n21 = n18 & n20 ;
  assign n22 = x9 & n21 ;
  assign n23 = x3 ^ x0 ;
  assign n31 = n23 ^ x0 ;
  assign n32 = x4 ^ x0 ;
  assign n33 = n32 ^ x2 ;
  assign n34 = n33 ^ x0 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = ~n31 & ~n35 ;
  assign n24 = n23 ^ x2 ;
  assign n25 = n24 ^ x0 ;
  assign n26 = n25 ^ x1 ;
  assign n27 = n25 & ~n26 ;
  assign n41 = n36 ^ n27 ;
  assign n28 = n27 ^ n23 ;
  assign n29 = n28 ^ n25 ;
  assign n30 = n29 ^ n22 ;
  assign n37 = n36 ^ n25 ;
  assign n38 = n37 ^ n31 ;
  assign n39 = n38 ^ n22 ;
  assign n40 = ~n30 & n39 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = ~n22 & n42 ;
  assign n44 = n43 ^ n36 ;
  assign n45 = n44 ^ n27 ;
  assign n46 = n45 ^ n40 ;
  assign n47 = ~n17 & n46 ;
  assign y0 = n47 ;
endmodule
