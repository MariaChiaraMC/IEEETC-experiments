module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 ;
  assign n16 = x6 & x7 ;
  assign n17 = ~x8 & n16 ;
  assign n18 = ~x3 & ~n17 ;
  assign n19 = ~x0 & ~x1 ;
  assign n20 = x13 & n19 ;
  assign n21 = ~x2 & ~x10 ;
  assign n22 = x9 & ~n21 ;
  assign n23 = n20 & ~n22 ;
  assign n24 = x12 & ~n19 ;
  assign n25 = ~x2 & n24 ;
  assign n26 = ~x3 & ~x4 ;
  assign n27 = n19 ^ x11 ;
  assign n28 = n27 ^ x11 ;
  assign n29 = x14 ^ x11 ;
  assign n30 = n28 & n29 ;
  assign n31 = n30 ^ x11 ;
  assign n32 = x2 & n31 ;
  assign n33 = ~n26 & n32 ;
  assign n34 = ~n25 & ~n33 ;
  assign n35 = ~n23 & n34 ;
  assign n36 = ~n18 & ~n35 ;
  assign n37 = ~n20 & ~n24 ;
  assign n38 = x7 ^ x6 ;
  assign n39 = n38 ^ x8 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = n38 ^ x7 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = ~n40 & n42 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = x5 & ~n44 ;
  assign n46 = n45 ^ n38 ;
  assign n47 = ~n37 & ~n46 ;
  assign n48 = ~x4 & n47 ;
  assign n49 = ~n36 & ~n48 ;
  assign y0 = ~n49 ;
endmodule
