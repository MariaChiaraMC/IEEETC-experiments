module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 ;
  assign n11 = ~x3 & x5 ;
  assign n12 = x0 & x7 ;
  assign n13 = n11 & n12 ;
  assign n14 = ~x4 & ~x8 ;
  assign n15 = n13 & n14 ;
  assign n16 = ~x0 & x3 ;
  assign n17 = ~x5 & x8 ;
  assign n18 = ~x7 & n17 ;
  assign n19 = x4 & n18 ;
  assign n20 = n16 & n19 ;
  assign n21 = ~n15 & ~n20 ;
  assign n22 = ~x2 & ~x9 ;
  assign n23 = ~n21 & n22 ;
  assign n24 = x1 & n23 ;
  assign n204 = x2 & ~x4 ;
  assign n129 = x8 ^ x7 ;
  assign n205 = n129 ^ x9 ;
  assign n206 = x9 ^ x5 ;
  assign n214 = n206 ^ x9 ;
  assign n215 = n214 ^ x9 ;
  assign n216 = ~n214 & ~n215 ;
  assign n208 = n206 ^ x1 ;
  assign n207 = n206 ^ x8 ;
  assign n209 = n208 ^ n207 ;
  assign n210 = n207 ^ n206 ;
  assign n211 = n210 ^ x9 ;
  assign n212 = ~n209 & n211 ;
  assign n219 = n216 ^ n212 ;
  assign n213 = n212 ^ n205 ;
  assign n217 = n216 ^ n214 ;
  assign n218 = n213 & ~n217 ;
  assign n220 = n219 ^ n218 ;
  assign n221 = n205 & n220 ;
  assign n222 = n221 ^ n212 ;
  assign n223 = n222 ^ n216 ;
  assign n224 = n223 ^ n218 ;
  assign n225 = n204 & n224 ;
  assign n92 = ~x4 & x9 ;
  assign n226 = x1 & ~x2 ;
  assign n227 = n92 & n226 ;
  assign n228 = n227 ^ x5 ;
  assign n229 = n228 ^ n18 ;
  assign n230 = n229 ^ n227 ;
  assign n231 = n230 ^ n229 ;
  assign n62 = x7 & ~x9 ;
  assign n232 = ~x8 & n62 ;
  assign n233 = n232 ^ x2 ;
  assign n234 = n233 ^ n232 ;
  assign n235 = n232 ^ x1 ;
  assign n236 = n234 & ~n235 ;
  assign n237 = n236 ^ n232 ;
  assign n66 = ~x7 & x9 ;
  assign n238 = ~n66 & ~n232 ;
  assign n239 = n238 ^ n14 ;
  assign n240 = ~n237 & ~n239 ;
  assign n241 = n240 ^ n238 ;
  assign n242 = ~n14 & n241 ;
  assign n243 = n242 ^ n14 ;
  assign n244 = n243 ^ n229 ;
  assign n245 = n244 ^ n228 ;
  assign n246 = n231 & n245 ;
  assign n247 = n246 ^ n243 ;
  assign n248 = x7 & ~x8 ;
  assign n249 = n243 & ~n248 ;
  assign n250 = n249 ^ n228 ;
  assign n251 = n247 & ~n250 ;
  assign n252 = n251 ^ n249 ;
  assign n253 = ~n228 & n252 ;
  assign n254 = n253 ^ n246 ;
  assign n255 = n254 ^ x5 ;
  assign n256 = n255 ^ n243 ;
  assign n257 = ~n225 & ~n256 ;
  assign n258 = x3 & ~n257 ;
  assign n46 = ~x1 & x4 ;
  assign n259 = ~x2 & n46 ;
  assign n43 = ~x8 & ~x9 ;
  assign n44 = ~x7 & n43 ;
  assign n260 = ~x5 & n44 ;
  assign n261 = n259 & n260 ;
  assign n166 = ~x3 & ~x5 ;
  assign n153 = x4 & ~x8 ;
  assign n262 = ~x1 & ~x2 ;
  assign n263 = ~n153 & n262 ;
  assign n25 = ~x4 & x8 ;
  assign n264 = ~x9 & n25 ;
  assign n265 = ~n263 & ~n264 ;
  assign n266 = ~x7 & ~n265 ;
  assign n267 = ~x1 & ~x4 ;
  assign n268 = n43 & n267 ;
  assign n269 = ~x2 & n268 ;
  assign n270 = n204 & n248 ;
  assign n169 = x4 & ~x7 ;
  assign n271 = n22 & ~n169 ;
  assign n272 = ~n14 & n271 ;
  assign n273 = ~n270 & ~n272 ;
  assign n274 = x1 & ~n273 ;
  assign n275 = ~n269 & ~n274 ;
  assign n276 = ~n266 & n275 ;
  assign n277 = n166 & ~n276 ;
  assign n278 = ~n261 & ~n277 ;
  assign n279 = ~n258 & n278 ;
  assign n280 = x0 & ~n279 ;
  assign n50 = ~x8 & x9 ;
  assign n167 = x8 & ~x9 ;
  assign n281 = ~n50 & ~n167 ;
  assign n91 = ~x5 & x7 ;
  assign n282 = ~x3 & n259 ;
  assign n74 = x1 & ~x3 ;
  assign n283 = n50 & n74 ;
  assign n284 = n204 & n283 ;
  assign n285 = ~n282 & ~n284 ;
  assign n286 = n91 & ~n285 ;
  assign n287 = ~n281 & n286 ;
  assign n65 = x1 & x3 ;
  assign n117 = x5 & ~x7 ;
  assign n288 = n14 & n117 ;
  assign n289 = ~n19 & ~n288 ;
  assign n290 = n22 & ~n289 ;
  assign n291 = n65 & n290 ;
  assign n121 = x0 & ~x3 ;
  assign n292 = ~x7 & n121 ;
  assign n93 = x4 & ~x9 ;
  assign n94 = ~n92 & ~n93 ;
  assign n293 = x4 & ~x5 ;
  assign n294 = x1 & x8 ;
  assign n295 = ~n293 & n294 ;
  assign n296 = n94 & n295 ;
  assign n297 = ~n268 & ~n296 ;
  assign n298 = n297 ^ n46 ;
  assign n299 = n298 ^ n297 ;
  assign n142 = x8 & x9 ;
  assign n300 = n297 ^ n142 ;
  assign n301 = n300 ^ n297 ;
  assign n302 = n299 & n301 ;
  assign n303 = n302 ^ n297 ;
  assign n304 = ~x2 & ~n303 ;
  assign n305 = n304 ^ n297 ;
  assign n306 = n292 & ~n305 ;
  assign n307 = ~n291 & ~n306 ;
  assign n308 = ~n287 & n307 ;
  assign n309 = ~n280 & n308 ;
  assign n310 = n93 & n166 ;
  assign n115 = x3 & x5 ;
  assign n52 = x9 & n25 ;
  assign n311 = ~x9 & n153 ;
  assign n312 = ~n52 & ~n311 ;
  assign n313 = n115 & ~n312 ;
  assign n314 = x1 & ~n313 ;
  assign n315 = ~n310 & n314 ;
  assign n147 = x5 & n50 ;
  assign n148 = ~x3 & n147 ;
  assign n316 = x4 & n148 ;
  assign n317 = ~x5 & ~x9 ;
  assign n103 = ~x3 & ~x4 ;
  assign n318 = x3 & x4 ;
  assign n319 = ~n103 & ~n318 ;
  assign n320 = n319 ^ x8 ;
  assign n321 = n320 ^ n319 ;
  assign n322 = n319 ^ x3 ;
  assign n323 = ~n321 & ~n322 ;
  assign n324 = n323 ^ n319 ;
  assign n325 = n317 & ~n324 ;
  assign n326 = ~x1 & ~n325 ;
  assign n327 = ~n316 & n326 ;
  assign n328 = x2 & ~n327 ;
  assign n329 = ~n315 & n328 ;
  assign n330 = n283 & n293 ;
  assign n331 = n17 & n92 ;
  assign n332 = n331 ^ x5 ;
  assign n333 = n332 ^ n331 ;
  assign n334 = n331 ^ n311 ;
  assign n335 = n334 ^ n331 ;
  assign n336 = n333 & n335 ;
  assign n337 = n336 ^ n331 ;
  assign n338 = ~x3 & n337 ;
  assign n339 = n338 ^ n331 ;
  assign n340 = n226 & n339 ;
  assign n341 = ~n330 & ~n340 ;
  assign n342 = ~n329 & n341 ;
  assign n343 = n342 ^ x7 ;
  assign n344 = n343 ^ n342 ;
  assign n345 = n344 ^ x0 ;
  assign n350 = n50 & n267 ;
  assign n352 = n350 ^ x5 ;
  assign n360 = n352 ^ n350 ;
  assign n351 = n350 ^ x9 ;
  assign n353 = n352 ^ n351 ;
  assign n354 = n353 ^ n352 ;
  assign n355 = n354 ^ n350 ;
  assign n356 = n353 ^ n294 ;
  assign n357 = n356 ^ n353 ;
  assign n358 = n357 ^ n355 ;
  assign n359 = ~n355 & ~n358 ;
  assign n361 = n360 ^ n359 ;
  assign n362 = n361 ^ n355 ;
  assign n363 = n350 ^ x4 ;
  assign n364 = n359 ^ n355 ;
  assign n365 = ~n363 & ~n364 ;
  assign n366 = n365 ^ n350 ;
  assign n367 = n362 & ~n366 ;
  assign n368 = n367 ^ n350 ;
  assign n369 = n368 ^ x5 ;
  assign n370 = n369 ^ n350 ;
  assign n371 = x3 & ~n370 ;
  assign n346 = n74 & n331 ;
  assign n108 = x4 & n74 ;
  assign n347 = ~n17 & n108 ;
  assign n348 = ~n281 & n347 ;
  assign n349 = ~n346 & ~n348 ;
  assign n372 = n371 ^ n349 ;
  assign n373 = n372 ^ n371 ;
  assign n374 = n115 & n167 ;
  assign n375 = ~n148 & ~n374 ;
  assign n376 = n267 & ~n375 ;
  assign n377 = n376 ^ n371 ;
  assign n378 = n377 ^ n371 ;
  assign n379 = n373 & ~n378 ;
  assign n380 = n379 ^ n371 ;
  assign n381 = x2 & ~n380 ;
  assign n382 = n381 ^ n371 ;
  assign n383 = n43 & n293 ;
  assign n384 = n65 & n383 ;
  assign n385 = n148 & n259 ;
  assign n386 = ~n384 & ~n385 ;
  assign n387 = n386 ^ n382 ;
  assign n388 = ~n382 & ~n387 ;
  assign n389 = n388 ^ n342 ;
  assign n390 = n389 ^ n382 ;
  assign n391 = n345 & ~n390 ;
  assign n392 = n391 ^ n388 ;
  assign n393 = n392 ^ n382 ;
  assign n394 = ~x0 & ~n393 ;
  assign n395 = n394 ^ x0 ;
  assign n396 = n309 & n395 ;
  assign n26 = x5 & n25 ;
  assign n27 = x7 ^ x3 ;
  assign n28 = n27 ^ x9 ;
  assign n29 = x9 ^ x0 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = x9 ^ x1 ;
  assign n32 = x7 ^ x1 ;
  assign n33 = ~n31 & ~n32 ;
  assign n34 = n33 ^ x1 ;
  assign n35 = n34 ^ n28 ;
  assign n36 = n30 & n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ x1 ;
  assign n39 = n38 ^ n29 ;
  assign n40 = ~n28 & n39 ;
  assign n41 = n40 ^ n28 ;
  assign n42 = n26 & ~n41 ;
  assign n45 = x7 & x8 ;
  assign n47 = ~n45 & n46 ;
  assign n48 = ~n44 & n47 ;
  assign n49 = n16 & ~n48 ;
  assign n51 = ~x7 & n50 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = n52 ^ x4 ;
  assign n56 = n55 ^ n52 ;
  assign n57 = ~n54 & ~n56 ;
  assign n58 = n57 ^ n52 ;
  assign n59 = ~x1 & ~n58 ;
  assign n60 = n59 ^ n52 ;
  assign n61 = n49 & n60 ;
  assign n63 = ~x3 & ~x8 ;
  assign n64 = n62 & n63 ;
  assign n67 = ~x9 & n45 ;
  assign n68 = ~n66 & ~n67 ;
  assign n69 = n65 & ~n68 ;
  assign n70 = ~n64 & ~n69 ;
  assign n71 = n70 ^ x4 ;
  assign n72 = n71 ^ n70 ;
  assign n73 = n72 ^ x0 ;
  assign n75 = ~n51 & ~n67 ;
  assign n76 = n74 & ~n75 ;
  assign n77 = ~n45 & ~n63 ;
  assign n78 = x9 & n77 ;
  assign n79 = ~x1 & n78 ;
  assign n80 = n79 ^ n76 ;
  assign n81 = ~n76 & n80 ;
  assign n82 = n81 ^ n70 ;
  assign n83 = n82 ^ n76 ;
  assign n84 = n73 & ~n83 ;
  assign n85 = n84 ^ n81 ;
  assign n86 = n85 ^ n76 ;
  assign n87 = x0 & ~n86 ;
  assign n88 = n87 ^ x0 ;
  assign n89 = ~n61 & ~n88 ;
  assign n90 = x5 & ~n89 ;
  assign n95 = n91 & ~n94 ;
  assign n96 = x0 & n95 ;
  assign n97 = x1 & ~n96 ;
  assign n98 = ~x5 & n66 ;
  assign n99 = ~n62 & ~n98 ;
  assign n100 = x4 & n16 ;
  assign n101 = ~n99 & n100 ;
  assign n102 = ~x0 & ~x9 ;
  assign n104 = ~x1 & ~n103 ;
  assign n105 = n91 & ~n104 ;
  assign n106 = ~n102 & n105 ;
  assign n107 = ~n101 & ~n106 ;
  assign n109 = ~n107 & ~n108 ;
  assign n110 = x8 & n109 ;
  assign n111 = ~n97 & n110 ;
  assign n112 = ~n90 & ~n111 ;
  assign n113 = n112 ^ x2 ;
  assign n114 = n113 ^ n112 ;
  assign n149 = ~x7 & n148 ;
  assign n150 = ~x4 & n64 ;
  assign n151 = ~n149 & ~n150 ;
  assign n152 = ~x0 & ~n151 ;
  assign n154 = n66 & n153 ;
  assign n155 = x5 & n67 ;
  assign n156 = ~n154 & ~n155 ;
  assign n157 = n16 & ~n156 ;
  assign n158 = ~n152 & ~n157 ;
  assign n122 = ~n91 & ~n117 ;
  assign n159 = x4 & x5 ;
  assign n160 = n142 & ~n159 ;
  assign n161 = ~n122 & n160 ;
  assign n162 = ~x3 & n161 ;
  assign n163 = n158 & ~n162 ;
  assign n116 = ~n66 & ~n115 ;
  assign n118 = ~x0 & ~x4 ;
  assign n119 = ~n117 & n118 ;
  assign n120 = ~n116 & n119 ;
  assign n123 = n93 & ~n122 ;
  assign n124 = n121 & n123 ;
  assign n125 = ~n120 & ~n124 ;
  assign n126 = ~x8 & ~n125 ;
  assign n127 = x9 ^ x4 ;
  assign n128 = n127 ^ n16 ;
  assign n130 = x8 ^ x4 ;
  assign n131 = n130 ^ x8 ;
  assign n132 = n129 & n131 ;
  assign n133 = n132 ^ x8 ;
  assign n134 = n133 ^ n127 ;
  assign n135 = ~n128 & ~n134 ;
  assign n136 = n135 ^ n132 ;
  assign n137 = n136 ^ x8 ;
  assign n138 = n137 ^ n16 ;
  assign n139 = ~n127 & n138 ;
  assign n140 = n139 ^ n127 ;
  assign n141 = ~x5 & ~n140 ;
  assign n143 = ~n14 & ~n142 ;
  assign n144 = n13 & ~n143 ;
  assign n145 = ~n141 & ~n144 ;
  assign n146 = ~n126 & n145 ;
  assign n164 = n163 ^ n146 ;
  assign n165 = n164 ^ n146 ;
  assign n168 = ~n166 & ~n167 ;
  assign n170 = ~n117 & ~n169 ;
  assign n171 = ~n168 & ~n170 ;
  assign n172 = x7 ^ x4 ;
  assign n173 = n172 ^ n50 ;
  assign n174 = x7 ^ x5 ;
  assign n175 = x5 ^ x3 ;
  assign n176 = n174 & ~n175 ;
  assign n177 = n176 ^ x5 ;
  assign n178 = n177 ^ n172 ;
  assign n179 = ~n173 & n178 ;
  assign n180 = n179 ^ n176 ;
  assign n181 = n180 ^ x5 ;
  assign n182 = n181 ^ n50 ;
  assign n183 = ~n172 & ~n182 ;
  assign n184 = n183 ^ n172 ;
  assign n185 = ~n171 & n184 ;
  assign n186 = x0 & ~n185 ;
  assign n187 = n186 ^ n146 ;
  assign n188 = n187 ^ n146 ;
  assign n189 = n165 & ~n188 ;
  assign n190 = n189 ^ n146 ;
  assign n191 = x1 & n190 ;
  assign n192 = n191 ^ n146 ;
  assign n193 = x0 & ~x9 ;
  assign n194 = ~n91 & ~n193 ;
  assign n195 = x4 & ~n62 ;
  assign n196 = ~n194 & n195 ;
  assign n197 = x8 & n196 ;
  assign n198 = ~n175 & n197 ;
  assign n199 = n192 & ~n198 ;
  assign n200 = n199 ^ n112 ;
  assign n201 = n114 & n200 ;
  assign n202 = n201 ^ n112 ;
  assign n203 = ~n42 & n202 ;
  assign n397 = n396 ^ n203 ;
  assign n398 = x6 & n397 ;
  assign n399 = n398 ^ n203 ;
  assign n400 = ~n24 & n399 ;
  assign y0 = ~n400 ;
endmodule
