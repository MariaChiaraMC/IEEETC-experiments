module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 ;
  assign n22 = x0 & ~x1 ;
  assign n23 = x5 & n22 ;
  assign n24 = ~x0 & x1 ;
  assign n25 = ~x2 & n24 ;
  assign n26 = ~n23 & ~n25 ;
  assign n27 = x5 ^ x3 ;
  assign n28 = ~x4 & ~n27 ;
  assign n29 = ~n26 & n28 ;
  assign n30 = ~x19 & ~x20 ;
  assign n31 = x2 & n22 ;
  assign n32 = ~x6 & ~x7 ;
  assign n33 = ~x12 & ~x13 ;
  assign n34 = n32 & n33 ;
  assign n35 = ~x5 & n34 ;
  assign n36 = n31 & n35 ;
  assign n37 = x10 ^ x8 ;
  assign n38 = x9 & x11 ;
  assign n39 = n38 ^ x11 ;
  assign n40 = x11 ^ x10 ;
  assign n41 = n40 ^ x11 ;
  assign n42 = ~n39 & ~n41 ;
  assign n43 = n42 ^ x11 ;
  assign n44 = n37 & ~n43 ;
  assign n45 = n36 & n44 ;
  assign n46 = x9 & x10 ;
  assign n47 = ~x12 & n46 ;
  assign n48 = x8 & n47 ;
  assign n49 = x12 & ~x13 ;
  assign n50 = x7 & ~x16 ;
  assign n51 = n49 & ~n50 ;
  assign n52 = ~x6 & n51 ;
  assign n53 = ~n48 & ~n52 ;
  assign n54 = x8 & n32 ;
  assign n55 = ~x16 & n54 ;
  assign n56 = ~x8 & x10 ;
  assign n57 = ~x11 & n56 ;
  assign n58 = x15 & n32 ;
  assign n59 = n57 & n58 ;
  assign n60 = ~n55 & ~n59 ;
  assign n62 = ~x9 & x10 ;
  assign n61 = x15 ^ x13 ;
  assign n63 = n62 ^ n61 ;
  assign n64 = n63 ^ n61 ;
  assign n65 = n63 ^ x15 ;
  assign n66 = n65 ^ n63 ;
  assign n67 = n66 ^ n61 ;
  assign n68 = n67 ^ n61 ;
  assign n69 = ~n64 & ~n68 ;
  assign n70 = n69 ^ n67 ;
  assign n71 = n67 ^ x12 ;
  assign n72 = n71 ^ n70 ;
  assign n73 = n46 ^ x11 ;
  assign n74 = ~n67 & ~n73 ;
  assign n75 = n74 ^ n46 ;
  assign n76 = n75 ^ n73 ;
  assign n77 = ~n72 & ~n76 ;
  assign n78 = n77 ^ n67 ;
  assign n79 = ~n70 & ~n78 ;
  assign n80 = n79 ^ n69 ;
  assign n81 = n80 ^ n67 ;
  assign n82 = n81 ^ x13 ;
  assign n83 = n60 & n82 ;
  assign n84 = x7 & x11 ;
  assign n85 = x9 & ~x12 ;
  assign n86 = n84 & n85 ;
  assign n87 = ~x13 & ~n86 ;
  assign n88 = x6 & ~n87 ;
  assign n89 = ~x17 & ~n88 ;
  assign n90 = x11 & n54 ;
  assign n91 = x11 & ~x16 ;
  assign n92 = ~x8 & ~n91 ;
  assign n93 = n92 ^ x13 ;
  assign n94 = n93 ^ n90 ;
  assign n95 = ~x10 & n32 ;
  assign n96 = n95 ^ n38 ;
  assign n97 = n92 & ~n96 ;
  assign n98 = n97 ^ n95 ;
  assign n99 = n94 & ~n98 ;
  assign n100 = n99 ^ n97 ;
  assign n101 = n100 ^ n95 ;
  assign n102 = n101 ^ n92 ;
  assign n103 = ~n90 & ~n102 ;
  assign n104 = n89 & n103 ;
  assign n105 = n83 & n104 ;
  assign n106 = n53 & n105 ;
  assign n107 = x2 & ~n106 ;
  assign n108 = ~x8 & x9 ;
  assign n109 = ~x12 & n108 ;
  assign n110 = ~x1 & n109 ;
  assign n111 = ~n47 & ~n110 ;
  assign n112 = x11 & ~n111 ;
  assign n113 = ~x12 & x13 ;
  assign n114 = n84 & n113 ;
  assign n115 = x13 ^ x1 ;
  assign n116 = n115 ^ n114 ;
  assign n117 = ~x10 & ~x11 ;
  assign n118 = n108 & n117 ;
  assign n119 = n118 ^ x0 ;
  assign n120 = ~x1 & n119 ;
  assign n121 = n120 ^ x0 ;
  assign n122 = ~n116 & n121 ;
  assign n123 = n122 ^ n120 ;
  assign n124 = n123 ^ x0 ;
  assign n125 = n124 ^ x1 ;
  assign n126 = ~n114 & ~n125 ;
  assign n127 = ~n112 & n126 ;
  assign n128 = ~n107 & n127 ;
  assign n129 = x5 & ~n128 ;
  assign n130 = ~n22 & ~n129 ;
  assign n131 = n130 ^ x4 ;
  assign n132 = n131 ^ n130 ;
  assign n133 = ~x11 & n108 ;
  assign n134 = ~n44 & ~n133 ;
  assign n135 = x1 & n35 ;
  assign n136 = ~n134 & n135 ;
  assign n137 = x2 & x5 ;
  assign n138 = ~x1 & ~x2 ;
  assign n139 = ~n137 & ~n138 ;
  assign n140 = ~x0 & n139 ;
  assign n141 = ~n136 & n140 ;
  assign n142 = x5 ^ x2 ;
  assign n143 = n142 ^ x5 ;
  assign n144 = n143 ^ x0 ;
  assign n145 = ~x11 & ~x13 ;
  assign n146 = x1 & n145 ;
  assign n147 = n146 ^ n48 ;
  assign n148 = n48 & n147 ;
  assign n149 = n148 ^ x5 ;
  assign n150 = n149 ^ n48 ;
  assign n151 = n144 & n150 ;
  assign n152 = n151 ^ n148 ;
  assign n153 = n152 ^ n48 ;
  assign n154 = x0 & n153 ;
  assign n155 = n154 ^ x0 ;
  assign n156 = ~n141 & ~n155 ;
  assign n157 = n156 ^ n130 ;
  assign n158 = ~n132 & ~n157 ;
  assign n159 = n158 ^ n130 ;
  assign n160 = ~n45 & n159 ;
  assign n161 = ~x3 & ~n160 ;
  assign n162 = x1 & n137 ;
  assign n163 = x3 & ~x4 ;
  assign n165 = x2 & ~n56 ;
  assign n164 = x0 & ~n117 ;
  assign n166 = n165 ^ n164 ;
  assign n167 = ~x9 & n166 ;
  assign n168 = n167 ^ n165 ;
  assign n169 = n163 & n168 ;
  assign n170 = ~x9 & ~x10 ;
  assign n171 = ~n145 & ~n170 ;
  assign n172 = n46 ^ n32 ;
  assign n173 = n172 ^ n46 ;
  assign n174 = n46 ^ x13 ;
  assign n175 = n174 ^ n46 ;
  assign n176 = ~n173 & ~n175 ;
  assign n177 = n176 ^ n46 ;
  assign n178 = ~x8 & ~n177 ;
  assign n179 = n178 ^ n46 ;
  assign n180 = ~n171 & n179 ;
  assign n181 = n169 & n180 ;
  assign n182 = n181 ^ n138 ;
  assign n183 = n182 ^ x3 ;
  assign n184 = n182 ^ n181 ;
  assign n185 = n184 ^ n183 ;
  assign n186 = ~n183 & ~n185 ;
  assign n187 = n186 ^ n182 ;
  assign n188 = n187 ^ n183 ;
  assign n189 = x13 ^ x12 ;
  assign n190 = n181 ^ x13 ;
  assign n191 = n189 & n190 ;
  assign n192 = n191 ^ n182 ;
  assign n193 = ~n188 & n192 ;
  assign n194 = n193 ^ n182 ;
  assign n195 = n194 ^ n181 ;
  assign n196 = n195 ^ x5 ;
  assign n197 = n196 ^ n195 ;
  assign n198 = n197 ^ n162 ;
  assign n199 = x3 & n24 ;
  assign n200 = ~n22 & ~n199 ;
  assign n201 = n200 ^ x4 ;
  assign n202 = x4 & ~n201 ;
  assign n203 = n202 ^ n195 ;
  assign n204 = n203 ^ x4 ;
  assign n205 = n198 & n204 ;
  assign n206 = n205 ^ n202 ;
  assign n207 = n206 ^ x4 ;
  assign n208 = ~n162 & n207 ;
  assign n209 = n208 ^ n162 ;
  assign n210 = ~n161 & ~n209 ;
  assign n211 = n210 ^ x18 ;
  assign n212 = n30 & n211 ;
  assign n213 = n212 ^ x18 ;
  assign n214 = ~n29 & n213 ;
  assign n215 = x14 & ~n214 ;
  assign y0 = n215 ;
endmodule
