module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n7 = x5 ^ x2 ;
  assign n17 = n7 ^ x0 ;
  assign n8 = n7 ^ x1 ;
  assign n9 = n8 ^ n7 ;
  assign n18 = n9 ^ x3 ;
  assign n19 = n17 & n18 ;
  assign n10 = x5 ^ x4 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = n10 ^ x5 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n11 & ~n13 ;
  assign n25 = n19 ^ n14 ;
  assign n15 = n14 ^ n9 ;
  assign n16 = n15 ^ n11 ;
  assign n20 = n10 ^ n7 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = n21 ^ n17 ;
  assign n23 = n22 ^ x3 ;
  assign n24 = n16 & ~n23 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n26 ^ n20 ;
  assign n28 = n27 ^ n17 ;
  assign n29 = n28 ^ x3 ;
  assign n30 = x3 & ~n29 ;
  assign n31 = n30 ^ x3 ;
  assign n32 = n31 ^ x5 ;
  assign n33 = n32 ^ x3 ;
  assign y0 = n33 ;
endmodule
