module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 ;
  assign n9 = x5 & x7 ;
  assign n10 = ~x4 & ~n9 ;
  assign n11 = ~x2 & x3 ;
  assign n12 = x6 & ~x7 ;
  assign n13 = ~n9 & ~n12 ;
  assign n14 = n11 & ~n13 ;
  assign n15 = ~n10 & n14 ;
  assign n16 = ~x1 & x7 ;
  assign n17 = ~x2 & x4 ;
  assign n18 = ~x1 & n17 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = ~n16 & ~n19 ;
  assign n21 = x4 & x6 ;
  assign n22 = ~x5 & ~x7 ;
  assign n23 = ~n9 & ~n22 ;
  assign n24 = n21 & ~n23 ;
  assign n25 = ~n20 & ~n24 ;
  assign n26 = x7 ^ x5 ;
  assign n27 = x6 ^ x1 ;
  assign n28 = n27 ^ x1 ;
  assign n29 = x4 ^ x1 ;
  assign n30 = ~n28 & n29 ;
  assign n31 = n30 ^ x1 ;
  assign n32 = n31 ^ x7 ;
  assign n33 = ~n26 & ~n32 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ x1 ;
  assign n36 = n35 ^ x5 ;
  assign n37 = ~x7 & n36 ;
  assign n38 = n37 ^ x7 ;
  assign n39 = n25 & n38 ;
  assign n40 = x5 ^ x4 ;
  assign n41 = n40 ^ x4 ;
  assign n42 = x7 ^ x4 ;
  assign n43 = ~n41 & n42 ;
  assign n44 = n43 ^ x4 ;
  assign n45 = x2 & n44 ;
  assign n46 = n39 & ~n45 ;
  assign n47 = n46 ^ x3 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = n48 ^ n15 ;
  assign n50 = x2 & ~n16 ;
  assign n51 = x6 & x7 ;
  assign n52 = ~n22 & ~n51 ;
  assign n53 = ~n50 & n52 ;
  assign n54 = n53 ^ x4 ;
  assign n55 = ~n53 & n54 ;
  assign n56 = n55 ^ n46 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = ~n49 & n57 ;
  assign n59 = n58 ^ n55 ;
  assign n60 = n59 ^ n53 ;
  assign n61 = ~n15 & ~n60 ;
  assign n62 = n61 ^ n15 ;
  assign n63 = ~x0 & n62 ;
  assign n64 = ~n17 & ~n21 ;
  assign n65 = ~x5 & n64 ;
  assign n66 = ~n11 & ~n65 ;
  assign n67 = ~x0 & ~n66 ;
  assign n68 = x3 & x7 ;
  assign n69 = ~x2 & ~x5 ;
  assign n70 = ~n68 & ~n69 ;
  assign n74 = x6 ^ x4 ;
  assign n75 = n74 ^ x7 ;
  assign n71 = x7 ^ x3 ;
  assign n73 = n71 ^ x6 ;
  assign n76 = n75 ^ n73 ;
  assign n72 = n71 ^ x7 ;
  assign n77 = n76 ^ n72 ;
  assign n78 = n77 ^ n76 ;
  assign n81 = x5 & x6 ;
  assign n82 = x2 & n81 ;
  assign n83 = x0 & n82 ;
  assign n84 = n83 ^ n76 ;
  assign n85 = ~n76 & n84 ;
  assign n79 = n71 & ~n75 ;
  assign n88 = n85 ^ n79 ;
  assign n80 = n79 ^ n78 ;
  assign n86 = n85 ^ n76 ;
  assign n87 = ~n80 & ~n86 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = ~n78 & n89 ;
  assign n91 = n90 ^ n85 ;
  assign n92 = n91 ^ n87 ;
  assign n93 = ~n70 & n92 ;
  assign n94 = ~n67 & ~n93 ;
  assign n95 = ~x1 & ~n94 ;
  assign n96 = x1 & ~x2 ;
  assign n97 = ~x3 & n96 ;
  assign n98 = n22 ^ x4 ;
  assign n99 = n98 ^ n22 ;
  assign n100 = n99 ^ n97 ;
  assign n101 = n9 ^ x6 ;
  assign n102 = ~n9 & ~n101 ;
  assign n103 = n102 ^ n22 ;
  assign n104 = n103 ^ n9 ;
  assign n105 = ~n100 & n104 ;
  assign n106 = n105 ^ n102 ;
  assign n107 = n106 ^ n9 ;
  assign n108 = n97 & ~n107 ;
  assign n109 = n108 ^ n97 ;
  assign n110 = ~n95 & ~n109 ;
  assign n111 = ~n63 & n110 ;
  assign y0 = ~n111 ;
endmodule
