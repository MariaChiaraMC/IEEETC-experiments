// Benchmark "./p3.pla" written by ABC on Thu Apr 23 11:00:00 2020

module \./p3.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z12  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z12;
  assign z12 = 1'b1;
endmodule


