module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 ;
  assign n21 = ~x7 & x17 ;
  assign n23 = x7 & ~x17 ;
  assign n42 = ~n21 & ~n23 ;
  assign n43 = x9 ^ x8 ;
  assign n44 = x18 ^ x9 ;
  assign n45 = n43 & n44 ;
  assign n46 = n45 ^ x8 ;
  assign n47 = n42 & ~n46 ;
  assign n22 = x8 & ~x18 ;
  assign n48 = x6 & ~n21 ;
  assign n49 = n22 & ~n48 ;
  assign n50 = ~n47 & ~n49 ;
  assign n35 = n22 & n23 ;
  assign n51 = ~x6 & ~n35 ;
  assign n52 = x16 & ~n51 ;
  assign n53 = ~x10 & x15 ;
  assign n54 = ~x2 & n53 ;
  assign n55 = n52 & n54 ;
  assign n56 = ~n50 & n55 ;
  assign n57 = x7 & n53 ;
  assign n58 = x15 & ~x18 ;
  assign n59 = x17 & ~n58 ;
  assign n60 = ~n57 & n59 ;
  assign n61 = ~x8 & n21 ;
  assign n62 = ~x6 & ~n61 ;
  assign n63 = x17 ^ x7 ;
  assign n64 = n63 ^ x2 ;
  assign n65 = x8 & x9 ;
  assign n66 = n65 ^ n46 ;
  assign n67 = ~x7 & ~n66 ;
  assign n68 = n67 ^ n46 ;
  assign n69 = n64 & ~n68 ;
  assign n70 = n69 ^ n67 ;
  assign n71 = n70 ^ n46 ;
  assign n72 = n71 ^ x7 ;
  assign n73 = ~x2 & n72 ;
  assign n74 = n62 & n73 ;
  assign n75 = ~x10 & ~n74 ;
  assign n76 = x12 & x13 ;
  assign n77 = x1 & ~x18 ;
  assign n78 = x10 & ~x11 ;
  assign n79 = n77 & n78 ;
  assign n80 = ~n76 & n79 ;
  assign n81 = n80 ^ x15 ;
  assign n82 = n81 ^ n80 ;
  assign n83 = n82 ^ x16 ;
  assign n84 = x18 ^ x17 ;
  assign n85 = ~x18 & n84 ;
  assign n86 = n85 ^ n80 ;
  assign n87 = n86 ^ x18 ;
  assign n88 = ~n83 & n87 ;
  assign n89 = n88 ^ n85 ;
  assign n90 = n89 ^ x18 ;
  assign n91 = ~x16 & ~n90 ;
  assign n92 = n91 ^ x16 ;
  assign n93 = ~n75 & ~n92 ;
  assign n94 = ~n60 & n93 ;
  assign n95 = ~n56 & ~n94 ;
  assign n20 = x16 ^ x6 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = ~x8 & x18 ;
  assign n27 = n26 ^ n22 ;
  assign n28 = n27 ^ n22 ;
  assign n29 = ~n25 & n28 ;
  assign n30 = n29 ^ n22 ;
  assign n31 = ~n21 & n30 ;
  assign n32 = n31 ^ n22 ;
  assign n33 = n32 ^ x16 ;
  assign n34 = n33 ^ n32 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ n32 ;
  assign n38 = n34 & n37 ;
  assign n39 = n38 ^ n32 ;
  assign n40 = n20 & n39 ;
  assign n41 = n40 ^ n32 ;
  assign n96 = n95 ^ n41 ;
  assign n97 = n96 ^ n95 ;
  assign n98 = n95 ^ x15 ;
  assign n99 = n98 ^ n95 ;
  assign n100 = n97 & ~n99 ;
  assign n101 = n100 ^ n95 ;
  assign n102 = x14 & ~n101 ;
  assign n103 = n102 ^ n95 ;
  assign y0 = ~n103 ;
endmodule
