// Benchmark "./p82.pla" written by ABC on Thu Apr 23 11:00:00 2020

module \./p82.pla  ( 
    x0, x1, x2, x3, x4,
    z9  );
  input  x0, x1, x2, x3, x4;
  output z9;
  assign z9 = ~x0 | ~x1;
endmodule


