module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 ;
  assign n9 = x3 & ~x6 ;
  assign n10 = x0 & ~n9 ;
  assign n11 = ~x5 & ~n10 ;
  assign n12 = ~x4 & ~n11 ;
  assign n13 = ~x1 & ~n12 ;
  assign n14 = x3 ^ x2 ;
  assign n15 = n14 ^ x0 ;
  assign n16 = ~x4 & ~x7 ;
  assign n17 = x6 & n16 ;
  assign n18 = n17 ^ x4 ;
  assign n19 = ~x2 & n18 ;
  assign n20 = n19 ^ x4 ;
  assign n21 = n15 & n20 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ x4 ;
  assign n24 = n23 ^ x2 ;
  assign n25 = ~x0 & ~n24 ;
  assign n26 = n25 ^ x2 ;
  assign n27 = n13 & ~n26 ;
  assign y0 = ~n27 ;
endmodule
