module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 ;
  assign n9 = x0 & ~x2 ;
  assign n10 = x6 ^ x1 ;
  assign n11 = ~x5 & n10 ;
  assign n12 = n11 ^ x1 ;
  assign n13 = ~x2 & ~n12 ;
  assign n14 = ~n9 & ~n13 ;
  assign n15 = ~x2 & x4 ;
  assign n16 = ~x0 & ~n15 ;
  assign n17 = x4 & x6 ;
  assign n18 = x5 & x7 ;
  assign n19 = n17 & n18 ;
  assign n20 = n16 & ~n19 ;
  assign n21 = ~x3 & ~n20 ;
  assign n22 = n14 & n21 ;
  assign n23 = ~x6 & ~x7 ;
  assign n24 = x5 & ~n23 ;
  assign n25 = n15 ^ x0 ;
  assign n26 = n25 ^ n15 ;
  assign n27 = ~x3 & ~x4 ;
  assign n28 = n27 ^ n15 ;
  assign n29 = n26 & n28 ;
  assign n30 = n29 ^ n15 ;
  assign n31 = ~n24 & n30 ;
  assign n32 = ~x5 & ~x6 ;
  assign n33 = ~x5 & ~x7 ;
  assign n34 = ~n32 & ~n33 ;
  assign n35 = ~n23 & n27 ;
  assign n36 = ~n34 & n35 ;
  assign n37 = ~x4 & x6 ;
  assign n38 = ~x3 & ~n37 ;
  assign n39 = n17 ^ x7 ;
  assign n40 = n39 ^ x7 ;
  assign n41 = ~x0 & x7 ;
  assign n42 = n41 ^ x7 ;
  assign n43 = ~n40 & ~n42 ;
  assign n44 = n43 ^ x7 ;
  assign n45 = x5 & ~n44 ;
  assign n46 = ~n38 & n45 ;
  assign n47 = ~n36 & ~n46 ;
  assign n48 = n47 ^ n27 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = ~x3 & n34 ;
  assign n51 = x5 & x6 ;
  assign n52 = ~x4 & ~n51 ;
  assign n53 = ~x4 & ~x7 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = ~n50 & n54 ;
  assign n56 = n55 ^ n47 ;
  assign n57 = n56 ^ n47 ;
  assign n58 = ~n49 & ~n57 ;
  assign n59 = n58 ^ n47 ;
  assign n60 = x2 & ~n59 ;
  assign n61 = n60 ^ n47 ;
  assign n62 = ~n31 & n61 ;
  assign n63 = ~x1 & ~n62 ;
  assign n64 = ~n17 & ~n52 ;
  assign n65 = ~x1 & ~n64 ;
  assign n66 = x4 & ~n33 ;
  assign n67 = ~x0 & ~n66 ;
  assign n68 = ~n65 & n67 ;
  assign n69 = ~x0 & x1 ;
  assign n70 = n32 & n53 ;
  assign n71 = ~n69 & ~n70 ;
  assign n72 = n71 ^ x2 ;
  assign n73 = n72 ^ n71 ;
  assign n74 = n73 ^ n68 ;
  assign n75 = x4 ^ x1 ;
  assign n76 = n18 ^ x4 ;
  assign n77 = n76 ^ n18 ;
  assign n78 = n34 ^ n18 ;
  assign n79 = ~n77 & ~n78 ;
  assign n80 = n79 ^ n18 ;
  assign n81 = n75 & n80 ;
  assign n82 = n81 ^ x1 ;
  assign n83 = n82 ^ x0 ;
  assign n84 = x0 & n83 ;
  assign n85 = n84 ^ n71 ;
  assign n86 = n85 ^ x0 ;
  assign n87 = n74 & ~n86 ;
  assign n88 = n87 ^ n84 ;
  assign n89 = n88 ^ x0 ;
  assign n90 = ~n68 & n89 ;
  assign n91 = n90 ^ n68 ;
  assign n92 = x3 & n91 ;
  assign n93 = n15 & n41 ;
  assign n94 = n32 & n93 ;
  assign n95 = ~n92 & ~n94 ;
  assign n96 = ~n63 & n95 ;
  assign n97 = ~n22 & n96 ;
  assign y0 = ~n97 ;
endmodule
