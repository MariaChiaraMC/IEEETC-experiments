module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n15 = x11 ^ x9 ;
  assign n16 = x11 ^ x10 ;
  assign n18 = n16 ^ x13 ;
  assign n17 = n16 ^ x12 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = n16 ^ x11 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = ~n18 & n22 ;
  assign n24 = n23 ^ n18 ;
  assign n25 = n19 & ~n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n26 ^ n16 ;
  assign n28 = n27 ^ n18 ;
  assign n29 = ~n15 & ~n28 ;
  assign n30 = n29 ^ x10 ;
  assign y0 = ~n30 ;
endmodule
