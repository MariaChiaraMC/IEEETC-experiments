module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 ;
  assign n15 = x3 & x11 ;
  assign n16 = x12 & n15 ;
  assign n17 = x10 & x13 ;
  assign n18 = n16 & n17 ;
  assign n19 = x9 & n18 ;
  assign n20 = ~x4 & ~x8 ;
  assign n21 = ~x6 & x7 ;
  assign n22 = ~x2 & n21 ;
  assign n23 = n20 & n22 ;
  assign n24 = x0 & ~n23 ;
  assign n25 = n24 ^ n19 ;
  assign n26 = ~x2 & x4 ;
  assign n27 = n26 ^ x1 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = x2 & ~n21 ;
  assign n30 = ~x0 & ~n29 ;
  assign n31 = ~x5 & ~n30 ;
  assign n32 = n31 ^ n26 ;
  assign n33 = ~n28 & n32 ;
  assign n34 = n33 ^ n26 ;
  assign n35 = n34 ^ n19 ;
  assign n36 = ~n25 & n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ n26 ;
  assign n39 = n38 ^ n24 ;
  assign n40 = n19 & ~n39 ;
  assign n41 = n40 ^ n19 ;
  assign y0 = n41 ;
endmodule
