module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 ;
  assign n121 = ~x11 & x14 ;
  assign n18 = ~x2 & ~x3 ;
  assign n19 = x7 & ~n18 ;
  assign n20 = ~x1 & n19 ;
  assign n21 = x6 ^ x0 ;
  assign n22 = ~x3 & ~x4 ;
  assign n23 = x2 & ~n22 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n24 ^ x6 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = ~x2 & ~x7 ;
  assign n28 = n27 ^ n24 ;
  assign n29 = n28 ^ n21 ;
  assign n30 = ~n26 & ~n29 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = x1 & ~n27 ;
  assign n33 = n32 ^ n21 ;
  assign n34 = ~n31 & ~n33 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = ~n21 & n35 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = n37 ^ x0 ;
  assign n39 = n38 ^ n27 ;
  assign n40 = ~n20 & ~n39 ;
  assign n41 = x5 & ~n40 ;
  assign n42 = x5 ^ x4 ;
  assign n43 = n42 ^ x6 ;
  assign n44 = n43 ^ x4 ;
  assign n45 = n44 ^ x4 ;
  assign n46 = x4 & ~n45 ;
  assign n47 = n46 ^ x4 ;
  assign n48 = n47 ^ n44 ;
  assign n49 = n48 ^ x3 ;
  assign n50 = n45 ^ x3 ;
  assign n51 = n27 ^ x6 ;
  assign n52 = n51 ^ x4 ;
  assign n53 = ~n50 & n52 ;
  assign n54 = n53 ^ x6 ;
  assign n55 = n54 ^ n44 ;
  assign n56 = x6 ^ x2 ;
  assign n57 = ~x2 & ~n56 ;
  assign n58 = n57 ^ x2 ;
  assign n59 = n58 ^ x4 ;
  assign n60 = n59 ^ n44 ;
  assign n61 = n60 ^ x3 ;
  assign n62 = ~n55 & n61 ;
  assign n63 = n62 ^ x4 ;
  assign n64 = ~n49 & n63 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = n65 ^ x4 ;
  assign n67 = x1 & n66 ;
  assign n68 = x3 & x5 ;
  assign n69 = x3 & ~x4 ;
  assign n70 = x0 & ~n69 ;
  assign n71 = x2 & n70 ;
  assign n72 = ~n68 & n71 ;
  assign n73 = ~n67 & ~n72 ;
  assign n74 = ~x0 & x1 ;
  assign n75 = n74 ^ x3 ;
  assign n76 = ~x5 & ~x7 ;
  assign n77 = ~x4 & n76 ;
  assign n78 = x2 & ~n77 ;
  assign n79 = n78 ^ n74 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = n80 ^ n75 ;
  assign n82 = ~x2 & ~x4 ;
  assign n83 = n82 ^ x5 ;
  assign n84 = n82 & n83 ;
  assign n85 = n84 ^ n78 ;
  assign n86 = n85 ^ n82 ;
  assign n87 = ~n81 & n86 ;
  assign n88 = n87 ^ n84 ;
  assign n89 = n88 ^ n82 ;
  assign n90 = n75 & n89 ;
  assign n91 = n90 ^ n74 ;
  assign n92 = x9 ^ x3 ;
  assign n93 = x0 & ~x1 ;
  assign n94 = n93 ^ x9 ;
  assign n95 = n94 ^ n93 ;
  assign n96 = ~x0 & n82 ;
  assign n97 = n96 ^ n93 ;
  assign n98 = n95 & n97 ;
  assign n99 = n98 ^ n93 ;
  assign n100 = n92 & ~n99 ;
  assign n101 = n100 ^ x3 ;
  assign n102 = ~n91 & ~n101 ;
  assign n103 = ~x13 & n102 ;
  assign n104 = n73 & n103 ;
  assign n105 = ~n41 & n104 ;
  assign n106 = n105 ^ x9 ;
  assign n107 = n105 ^ x13 ;
  assign n108 = n107 ^ x13 ;
  assign n109 = n108 ^ n106 ;
  assign n110 = n96 ^ x5 ;
  assign n111 = n96 & n110 ;
  assign n112 = n111 ^ x13 ;
  assign n113 = n112 ^ n96 ;
  assign n114 = n109 & n113 ;
  assign n115 = n114 ^ n111 ;
  assign n116 = n115 ^ n96 ;
  assign n117 = n106 & n116 ;
  assign n118 = n117 ^ n105 ;
  assign n119 = ~x10 & n118 ;
  assign n16 = x10 & ~x13 ;
  assign n17 = x9 & n16 ;
  assign n120 = n119 ^ n17 ;
  assign n122 = n121 ^ n120 ;
  assign n130 = n122 ^ n120 ;
  assign n123 = ~x11 & ~n16 ;
  assign n124 = n123 ^ n122 ;
  assign n125 = n124 ^ n120 ;
  assign n126 = n122 ^ n17 ;
  assign n127 = n126 ^ n123 ;
  assign n128 = n127 ^ n125 ;
  assign n129 = n125 & n128 ;
  assign n131 = n130 ^ n129 ;
  assign n132 = n131 ^ n125 ;
  assign n133 = ~n18 & n93 ;
  assign n134 = n133 ^ n120 ;
  assign n135 = n129 ^ n125 ;
  assign n136 = ~n134 & n135 ;
  assign n137 = n136 ^ n120 ;
  assign n138 = ~n132 & ~n137 ;
  assign n139 = n138 ^ n120 ;
  assign n140 = n139 ^ n119 ;
  assign n141 = n140 ^ n120 ;
  assign y0 = ~n141 ;
endmodule
