// Benchmark "./m3.pla" written by ABC on Thu Apr 23 10:59:55 2020

module \./m3.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z1  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z1;
  assign z1 = 1'b1;
endmodule


