module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 ;
  output y0 ;
  wire n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 ;
  assign n19 = ~x0 & ~x14 ;
  assign n20 = x16 ^ x6 ;
  assign n28 = n20 ^ x13 ;
  assign n21 = n20 ^ x16 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n20 ^ x15 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = ~n22 & n24 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = n26 ^ x13 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = x15 ^ x5 ;
  assign n31 = n30 ^ n20 ;
  assign n32 = n31 ^ x13 ;
  assign n33 = n32 ^ n28 ;
  assign n34 = ~x13 & ~n33 ;
  assign n35 = n34 ^ n28 ;
  assign n36 = ~x7 & ~x8 ;
  assign n37 = x3 & n36 ;
  assign n38 = n28 & ~n37 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = n39 ^ n31 ;
  assign n41 = n40 ^ n28 ;
  assign n42 = n35 & ~n41 ;
  assign n43 = n42 ^ x13 ;
  assign n44 = n43 ^ n31 ;
  assign n45 = n29 & ~n44 ;
  assign n46 = n45 ^ x13 ;
  assign n47 = n46 ^ n28 ;
  assign n48 = n47 ^ n20 ;
  assign n49 = ~x17 & n48 ;
  assign n54 = ~x5 & x15 ;
  assign n50 = x5 & ~x15 ;
  assign n51 = x7 & ~n50 ;
  assign n52 = x16 & ~n51 ;
  assign n53 = ~x17 & ~n52 ;
  assign n55 = n54 ^ n53 ;
  assign n56 = n53 ^ x7 ;
  assign n57 = n56 ^ n55 ;
  assign n58 = x6 & x16 ;
  assign n59 = ~x6 & ~x16 ;
  assign n60 = ~n58 & ~n59 ;
  assign n61 = ~n50 & ~n60 ;
  assign n62 = n61 ^ x16 ;
  assign n63 = x7 & ~n62 ;
  assign n64 = n63 ^ n61 ;
  assign n65 = n57 & ~n64 ;
  assign n66 = n65 ^ n63 ;
  assign n67 = n66 ^ n61 ;
  assign n68 = n67 ^ x7 ;
  assign n69 = ~n55 & ~n68 ;
  assign n70 = n69 ^ n54 ;
  assign n71 = n70 ^ x13 ;
  assign n72 = n71 ^ n70 ;
  assign n100 = x3 & ~n36 ;
  assign n101 = ~n60 & n100 ;
  assign n73 = x3 & x8 ;
  assign n74 = n73 ^ n51 ;
  assign n75 = n54 ^ x6 ;
  assign n76 = n75 ^ x6 ;
  assign n77 = n20 & ~n76 ;
  assign n78 = n77 ^ x6 ;
  assign n79 = n78 ^ n73 ;
  assign n80 = n74 & n79 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n81 ^ x6 ;
  assign n83 = n82 ^ n51 ;
  assign n84 = n73 & n83 ;
  assign n85 = n84 ^ n73 ;
  assign n86 = ~n58 & n85 ;
  assign n87 = ~x4 & ~x16 ;
  assign n88 = ~x9 & ~x15 ;
  assign n89 = x1 & x2 ;
  assign n90 = n88 & n89 ;
  assign n91 = n87 & n90 ;
  assign n92 = x11 ^ x10 ;
  assign n93 = n92 ^ n90 ;
  assign n94 = x11 & ~x12 ;
  assign n95 = n94 ^ n91 ;
  assign n96 = ~n93 & n95 ;
  assign n97 = n96 ^ n94 ;
  assign n98 = n91 & n97 ;
  assign n99 = ~n86 & ~n98 ;
  assign n102 = n101 ^ n99 ;
  assign n103 = n102 ^ n99 ;
  assign n104 = x7 & x8 ;
  assign n105 = ~n30 & ~n104 ;
  assign n106 = n105 ^ n99 ;
  assign n107 = n106 ^ n99 ;
  assign n108 = n103 & n107 ;
  assign n109 = n108 ^ n99 ;
  assign n110 = x17 & ~n109 ;
  assign n111 = n110 ^ n99 ;
  assign n112 = n111 ^ n70 ;
  assign n113 = ~n72 & ~n112 ;
  assign n114 = n113 ^ n70 ;
  assign n115 = ~n49 & ~n114 ;
  assign n116 = n19 & ~n115 ;
  assign y0 = n116 ;
endmodule
