module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 ;
  assign n9 = ~x6 & ~x7 ;
  assign n10 = x4 & ~n9 ;
  assign n11 = x5 & n10 ;
  assign n12 = ~x2 & ~x3 ;
  assign n13 = ~x4 & ~x6 ;
  assign n14 = ~n12 & ~n13 ;
  assign n15 = ~x4 & ~x5 ;
  assign n16 = x2 & x3 ;
  assign n17 = ~n15 & ~n16 ;
  assign n18 = n14 & n17 ;
  assign n19 = ~n11 & n18 ;
  assign n20 = x3 ^ x2 ;
  assign n29 = n20 ^ x4 ;
  assign n30 = n29 ^ n20 ;
  assign n31 = n30 ^ x5 ;
  assign n21 = x5 ^ x3 ;
  assign n22 = n21 ^ x5 ;
  assign n32 = n22 ^ n20 ;
  assign n33 = n31 & n32 ;
  assign n23 = x6 ^ x5 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = n26 ^ n20 ;
  assign n28 = ~n20 & n27 ;
  assign n34 = n33 ^ n28 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n35 ^ n20 ;
  assign n37 = n36 ^ n31 ;
  assign n38 = n29 ^ x7 ;
  assign n39 = n38 ^ n20 ;
  assign n40 = n39 ^ n20 ;
  assign n41 = ~n22 & ~n40 ;
  assign n42 = n41 ^ n33 ;
  assign n43 = n42 ^ n30 ;
  assign n44 = n43 ^ n31 ;
  assign n45 = n31 & ~n44 ;
  assign n46 = n45 ^ n20 ;
  assign n47 = n46 ^ n31 ;
  assign n48 = n37 & ~n47 ;
  assign n49 = n48 ^ n28 ;
  assign n50 = ~n19 & ~n49 ;
  assign n51 = ~x1 & ~n50 ;
  assign n52 = x6 & n15 ;
  assign n53 = ~x1 & ~n52 ;
  assign n54 = n12 & ~n53 ;
  assign n55 = ~n11 & n54 ;
  assign n56 = ~x0 & ~n55 ;
  assign n57 = ~n51 & n56 ;
  assign y0 = n57 ;
endmodule
