module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 ;
  assign n12 = x5 & x6 ;
  assign n13 = x7 & n12 ;
  assign n16 = ~x9 & ~x10 ;
  assign n17 = ~x4 & n16 ;
  assign n18 = n17 ^ x10 ;
  assign n19 = n13 & ~n18 ;
  assign n20 = x10 ^ x7 ;
  assign n21 = n20 ^ x9 ;
  assign n22 = x4 & n12 ;
  assign n23 = n22 ^ x6 ;
  assign n24 = ~x7 & ~n23 ;
  assign n25 = n24 ^ x6 ;
  assign n26 = n21 & ~n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n27 ^ x6 ;
  assign n29 = n28 ^ x7 ;
  assign n30 = ~x9 & n29 ;
  assign n31 = ~n19 & ~n30 ;
  assign n14 = ~x10 & ~n13 ;
  assign n15 = x9 & ~n14 ;
  assign n32 = n31 ^ n15 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = x3 & x4 ;
  assign n35 = n12 & n34 ;
  assign n36 = x5 & n34 ;
  assign n37 = ~x6 & ~n36 ;
  assign n38 = x7 & ~n37 ;
  assign n39 = ~n35 & n38 ;
  assign n40 = x1 & x2 ;
  assign n43 = x0 & n40 ;
  assign n44 = ~n34 & n43 ;
  assign n41 = x3 & n40 ;
  assign n42 = n41 ^ x4 ;
  assign n45 = n44 ^ n42 ;
  assign n46 = n45 ^ n42 ;
  assign n47 = x3 ^ x2 ;
  assign n48 = x4 & n47 ;
  assign n49 = n48 ^ x2 ;
  assign n50 = ~n43 & n49 ;
  assign n51 = n50 ^ n42 ;
  assign n52 = n51 ^ n42 ;
  assign n53 = ~n46 & ~n52 ;
  assign n54 = n53 ^ n42 ;
  assign n55 = ~x5 & ~n54 ;
  assign n56 = n55 ^ n42 ;
  assign n57 = n56 ^ x6 ;
  assign n58 = n57 ^ n56 ;
  assign n59 = x2 & n34 ;
  assign n60 = n59 ^ x5 ;
  assign n61 = n60 ^ n56 ;
  assign n62 = n58 & n61 ;
  assign n63 = n62 ^ n56 ;
  assign n64 = ~x7 & n63 ;
  assign n65 = ~n39 & ~n64 ;
  assign n66 = n16 & ~n65 ;
  assign n67 = n66 ^ n31 ;
  assign n68 = n67 ^ n31 ;
  assign n69 = ~n33 & ~n68 ;
  assign n70 = n69 ^ n31 ;
  assign n71 = ~x8 & ~n70 ;
  assign n72 = n71 ^ n31 ;
  assign y0 = n72 ;
endmodule
