// Benchmark "./pla/pdc.pla_dbb_orig_14NonExact" written by ABC on Fri Nov 20 10:27:51 2020

module \./pla/pdc.pla_dbb_orig_14NonExact  ( 
    x0, x1,
    z0  );
  input  x0, x1;
  output z0;
  assign z0 = x0 & ~x1;
endmodule


