module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 ;
  assign n25 = x14 & ~x20 ;
  assign n26 = ~x19 & n25 ;
  assign n27 = ~x0 & x5 ;
  assign n28 = x1 & x2 ;
  assign n29 = n27 & n28 ;
  assign n30 = x5 ^ x1 ;
  assign n31 = ~x2 & x3 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = x21 ^ x5 ;
  assign n34 = n33 ^ x21 ;
  assign n35 = x21 ^ x0 ;
  assign n36 = ~n34 & ~n35 ;
  assign n37 = n36 ^ x21 ;
  assign n38 = n37 ^ n30 ;
  assign n39 = n32 & n38 ;
  assign n40 = n39 ^ n36 ;
  assign n41 = n40 ^ x21 ;
  assign n42 = n41 ^ n31 ;
  assign n43 = n30 & n42 ;
  assign n44 = n43 ^ n30 ;
  assign n45 = ~n29 & ~n44 ;
  assign n46 = x3 ^ x1 ;
  assign n47 = n46 ^ x1 ;
  assign n48 = n30 & n47 ;
  assign n49 = n48 ^ x1 ;
  assign n50 = x1 & x23 ;
  assign n51 = n50 ^ x0 ;
  assign n52 = n49 & n51 ;
  assign n53 = n52 ^ n50 ;
  assign n54 = x0 & n53 ;
  assign n55 = n54 ^ x0 ;
  assign n56 = n55 ^ x3 ;
  assign n57 = n56 ^ n45 ;
  assign n58 = ~x6 & ~x7 ;
  assign n59 = x12 & ~x13 ;
  assign n60 = ~x10 & ~x16 ;
  assign n61 = ~x8 & ~n60 ;
  assign n62 = x15 & ~n61 ;
  assign n63 = x11 & n62 ;
  assign n64 = ~n59 & ~n63 ;
  assign n65 = n58 & ~n64 ;
  assign n66 = ~x9 & x10 ;
  assign n67 = ~x6 & ~n66 ;
  assign n68 = x13 & ~n67 ;
  assign n69 = x9 & x10 ;
  assign n70 = ~x13 & ~n69 ;
  assign n71 = ~n59 & ~n70 ;
  assign n72 = ~x11 & n58 ;
  assign n73 = x10 & n72 ;
  assign n74 = ~x8 & n73 ;
  assign n75 = ~n71 & ~n74 ;
  assign n76 = x15 & ~n75 ;
  assign n77 = x8 & n58 ;
  assign n78 = ~x13 & ~n77 ;
  assign n79 = ~x10 & ~x11 ;
  assign n80 = ~n78 & n79 ;
  assign n81 = ~x17 & ~n80 ;
  assign n82 = ~n76 & n81 ;
  assign n83 = ~n68 & n82 ;
  assign n84 = x11 & ~x12 ;
  assign n85 = ~x8 & n84 ;
  assign n86 = x11 ^ x10 ;
  assign n87 = x6 & x7 ;
  assign n88 = n87 ^ x11 ;
  assign n89 = n88 ^ x11 ;
  assign n90 = n89 ^ n86 ;
  assign n91 = x18 ^ x8 ;
  assign n92 = ~x11 & n91 ;
  assign n93 = n92 ^ x18 ;
  assign n94 = n90 & n93 ;
  assign n95 = n94 ^ n92 ;
  assign n96 = n95 ^ x18 ;
  assign n97 = n96 ^ x11 ;
  assign n98 = n86 & ~n97 ;
  assign n99 = n98 ^ x10 ;
  assign n100 = n99 ^ x13 ;
  assign n101 = ~x12 & n100 ;
  assign n102 = n101 ^ x13 ;
  assign n103 = ~n85 & ~n102 ;
  assign n104 = x9 & ~n103 ;
  assign n105 = x10 & x11 ;
  assign n106 = x7 & n105 ;
  assign n107 = ~x13 & ~n106 ;
  assign n108 = x8 & ~n107 ;
  assign n109 = ~n59 & n108 ;
  assign n110 = x8 & x10 ;
  assign n111 = n84 & n110 ;
  assign n112 = ~x6 & n111 ;
  assign n113 = ~x1 & ~n112 ;
  assign n114 = ~n109 & n113 ;
  assign n115 = ~n104 & n114 ;
  assign n116 = n83 & n115 ;
  assign n117 = ~n65 & n116 ;
  assign n118 = x2 & ~n117 ;
  assign n119 = ~x0 & x1 ;
  assign n120 = x15 & n119 ;
  assign n121 = ~x13 & ~n84 ;
  assign n122 = x0 & ~n70 ;
  assign n123 = ~n121 & n122 ;
  assign n124 = ~n120 & ~n123 ;
  assign n125 = ~n118 & n124 ;
  assign n126 = x5 & ~n125 ;
  assign n127 = n126 ^ x2 ;
  assign n128 = x3 & ~n127 ;
  assign n129 = n128 ^ n126 ;
  assign n130 = ~n57 & ~n129 ;
  assign n131 = n130 ^ n128 ;
  assign n132 = n131 ^ n126 ;
  assign n133 = n132 ^ x3 ;
  assign n134 = n45 & ~n133 ;
  assign n135 = x4 & ~n134 ;
  assign n139 = ~x4 & x5 ;
  assign n136 = x3 & ~n27 ;
  assign n137 = ~x1 & ~x2 ;
  assign n138 = ~n136 & n137 ;
  assign n140 = n139 ^ n138 ;
  assign n141 = ~x4 & ~x15 ;
  assign n142 = x23 & n141 ;
  assign n143 = x22 & n142 ;
  assign n144 = ~x3 & ~n143 ;
  assign n145 = ~x0 & ~n144 ;
  assign n146 = n145 ^ n138 ;
  assign n147 = n146 ^ n145 ;
  assign n148 = n147 ^ n140 ;
  assign n149 = n28 ^ x3 ;
  assign n150 = n28 & n149 ;
  assign n151 = n150 ^ n145 ;
  assign n152 = n151 ^ n28 ;
  assign n153 = ~n148 & ~n152 ;
  assign n154 = n153 ^ n150 ;
  assign n155 = n154 ^ n28 ;
  assign n156 = n140 & n155 ;
  assign n157 = n156 ^ n138 ;
  assign n158 = ~n135 & ~n157 ;
  assign n159 = n26 & ~n158 ;
  assign y0 = n159 ;
endmodule
