module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 ;
  assign n11 = x3 & x4 ;
  assign n12 = x2 & ~x5 ;
  assign n13 = ~x1 & x6 ;
  assign n14 = ~x7 & n13 ;
  assign n15 = n12 & n14 ;
  assign n16 = n11 & n15 ;
  assign n19 = x5 ^ x2 ;
  assign n38 = ~x3 & x7 ;
  assign n39 = ~x4 & n38 ;
  assign n40 = n39 ^ x5 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = n39 ^ x7 ;
  assign n43 = n42 ^ n39 ;
  assign n44 = n41 & ~n43 ;
  assign n45 = n44 ^ n39 ;
  assign n46 = ~n11 & ~n39 ;
  assign n47 = n46 ^ n19 ;
  assign n48 = ~n45 & n47 ;
  assign n49 = n48 ^ n46 ;
  assign n50 = n19 & n49 ;
  assign n51 = n50 ^ n39 ;
  assign n52 = n51 ^ n19 ;
  assign n53 = x1 & n52 ;
  assign n17 = ~x4 & ~x7 ;
  assign n18 = ~n11 & ~n17 ;
  assign n20 = x5 ^ x1 ;
  assign n21 = n19 & ~n20 ;
  assign n22 = n18 & n21 ;
  assign n23 = n22 ^ x3 ;
  assign n24 = n22 ^ x7 ;
  assign n25 = n24 ^ x7 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = x7 ^ x4 ;
  assign n28 = x1 & ~n27 ;
  assign n29 = n28 ^ n12 ;
  assign n30 = n12 & n29 ;
  assign n31 = n30 ^ x7 ;
  assign n32 = n31 ^ n12 ;
  assign n33 = ~n26 & n32 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ n12 ;
  assign n36 = n23 & n35 ;
  assign n37 = n36 ^ n22 ;
  assign n54 = n53 ^ n37 ;
  assign n55 = n54 ^ n37 ;
  assign n56 = ~x1 & x7 ;
  assign n57 = ~x2 & x5 ;
  assign n58 = n56 & n57 ;
  assign n59 = n58 ^ n37 ;
  assign n60 = n59 ^ n37 ;
  assign n61 = ~n55 & ~n60 ;
  assign n62 = n61 ^ n37 ;
  assign n63 = x6 & ~n62 ;
  assign n64 = n63 ^ n37 ;
  assign n65 = n64 ^ x0 ;
  assign n66 = n65 ^ n64 ;
  assign n70 = ~x3 & ~x4 ;
  assign n71 = x2 & ~n70 ;
  assign n68 = ~x6 & x7 ;
  assign n67 = x6 & ~x7 ;
  assign n69 = n68 ^ n67 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = n72 ^ n69 ;
  assign n74 = n73 ^ x1 ;
  assign n75 = n67 ^ n11 ;
  assign n76 = n11 & n75 ;
  assign n77 = n76 ^ n69 ;
  assign n78 = n77 ^ n11 ;
  assign n79 = ~n74 & n78 ;
  assign n80 = n79 ^ n76 ;
  assign n81 = n80 ^ n11 ;
  assign n82 = ~x1 & n81 ;
  assign n83 = n82 ^ n67 ;
  assign n84 = ~x5 & n83 ;
  assign n85 = n84 ^ n64 ;
  assign n86 = n66 & n85 ;
  assign n87 = n86 ^ n64 ;
  assign n88 = ~n16 & ~n87 ;
  assign n89 = ~x8 & n88 ;
  assign n90 = x2 & x5 ;
  assign n91 = n39 & n90 ;
  assign n92 = n13 & n91 ;
  assign n93 = n92 ^ x0 ;
  assign n94 = n93 ^ n92 ;
  assign n95 = x7 ^ x1 ;
  assign n96 = x6 ^ x3 ;
  assign n97 = n95 & ~n96 ;
  assign n98 = n97 ^ x3 ;
  assign n99 = n98 ^ n97 ;
  assign n100 = x6 ^ x1 ;
  assign n101 = x7 ^ x6 ;
  assign n102 = n100 & n101 ;
  assign n103 = n102 ^ n97 ;
  assign n104 = n103 ^ n97 ;
  assign n105 = ~n99 & n104 ;
  assign n106 = n105 ^ n97 ;
  assign n107 = x4 & n106 ;
  assign n108 = n107 ^ n97 ;
  assign n109 = n90 & n108 ;
  assign n110 = ~x5 & n28 ;
  assign n111 = ~x2 & n110 ;
  assign n112 = ~n96 & n111 ;
  assign n113 = ~n109 & ~n112 ;
  assign n114 = n113 ^ n92 ;
  assign n115 = ~n94 & ~n114 ;
  assign n116 = n115 ^ n92 ;
  assign n117 = x8 & ~n116 ;
  assign n118 = ~x9 & ~n117 ;
  assign n119 = ~n89 & n118 ;
  assign y0 = n119 ;
endmodule
