module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 ;
  assign n9 = x2 & ~x4 ;
  assign n10 = x3 & ~n9 ;
  assign n12 = x2 & ~x3 ;
  assign n13 = ~x0 & ~x1 ;
  assign n14 = ~n12 & n13 ;
  assign n15 = x5 & n14 ;
  assign n11 = x0 & x1 ;
  assign n16 = n15 ^ n11 ;
  assign n17 = n16 ^ n11 ;
  assign n18 = x6 & x7 ;
  assign n19 = n18 ^ n11 ;
  assign n20 = n19 ^ n11 ;
  assign n21 = n17 & n20 ;
  assign n22 = n21 ^ n11 ;
  assign n23 = ~x4 & n22 ;
  assign n24 = n23 ^ n11 ;
  assign n25 = ~n10 & n24 ;
  assign y0 = ~n25 ;
endmodule
