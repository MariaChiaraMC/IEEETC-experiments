module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 ;
  assign n9 = x2 & x7 ;
  assign n10 = ~x6 & ~n9 ;
  assign n11 = ~x5 & ~n10 ;
  assign n13 = x4 ^ x2 ;
  assign n12 = x6 ^ x4 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n14 ^ n12 ;
  assign n20 = n15 ^ x4 ;
  assign n18 = x7 ^ x4 ;
  assign n16 = x4 ^ x1 ;
  assign n17 = n16 ^ n15 ;
  assign n19 = n18 ^ n17 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = n15 ^ n12 ;
  assign n23 = n22 ^ n17 ;
  assign n24 = n21 & n23 ;
  assign n25 = n24 ^ n15 ;
  assign n29 = n20 ^ n15 ;
  assign n30 = n17 ^ n15 ;
  assign n31 = n30 ^ n20 ;
  assign n32 = ~n29 & ~n31 ;
  assign n26 = x5 ^ x4 ;
  assign n27 = n22 ^ n20 ;
  assign n28 = n26 & ~n27 ;
  assign n33 = n32 ^ n28 ;
  assign n34 = n33 ^ n20 ;
  assign n35 = n34 ^ n22 ;
  assign n36 = n22 & ~n35 ;
  assign n37 = n36 ^ n28 ;
  assign n38 = n37 ^ n15 ;
  assign n39 = n38 ^ n22 ;
  assign n40 = n25 & n39 ;
  assign n41 = n40 ^ n32 ;
  assign n42 = n41 ^ n15 ;
  assign n43 = n42 ^ n20 ;
  assign n44 = n43 ^ x4 ;
  assign n45 = ~n11 & ~n44 ;
  assign y0 = ~n45 ;
endmodule
