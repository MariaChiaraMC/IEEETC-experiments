module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 ;
  assign n8 = ~x0 & x2 ;
  assign n9 = x4 & n8 ;
  assign n10 = x6 ^ x0 ;
  assign n11 = n10 ^ x6 ;
  assign n12 = n11 ^ x1 ;
  assign n13 = n12 ^ x1 ;
  assign n14 = n13 ^ n10 ;
  assign n15 = n10 ^ x5 ;
  assign n16 = n15 ^ x1 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = ~n14 & ~n18 ;
  assign n20 = n19 ^ n15 ;
  assign n21 = x3 & x4 ;
  assign n22 = n21 ^ x1 ;
  assign n23 = n22 ^ n13 ;
  assign n24 = n22 ^ n15 ;
  assign n25 = n23 & n24 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = n26 ^ n14 ;
  assign n28 = n21 ^ n14 ;
  assign n29 = x2 & n28 ;
  assign n30 = n29 ^ x2 ;
  assign n31 = n30 ^ n15 ;
  assign n32 = n31 ^ n13 ;
  assign n33 = n32 ^ n14 ;
  assign n34 = n27 & ~n33 ;
  assign n35 = n34 ^ n13 ;
  assign n36 = n35 ^ n14 ;
  assign n37 = ~n20 & n36 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = n38 ^ n13 ;
  assign n40 = n39 ^ n14 ;
  assign n41 = n40 ^ x0 ;
  assign n42 = ~n9 & ~n41 ;
  assign y0 = n42 ;
endmodule
