module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 ;
  assign n12 = x7 & ~x8 ;
  assign n13 = x3 & ~x5 ;
  assign n14 = ~n12 & ~n13 ;
  assign n15 = n14 ^ x3 ;
  assign n16 = n15 ^ x4 ;
  assign n24 = n16 ^ n15 ;
  assign n17 = ~x5 & x8 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n16 ^ n14 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n19 & n22 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ n19 ;
  assign n27 = n15 ^ x6 ;
  assign n28 = n23 ^ n19 ;
  assign n29 = n27 & n28 ;
  assign n30 = n29 ^ n15 ;
  assign n31 = ~n26 & n30 ;
  assign n32 = n31 ^ n15 ;
  assign n33 = n32 ^ x3 ;
  assign n34 = n33 ^ n15 ;
  assign n10 = x8 ^ x2 ;
  assign n11 = n10 ^ x8 ;
  assign n35 = n34 ^ n11 ;
  assign n36 = n35 ^ n34 ;
  assign n38 = x7 ^ x6 ;
  assign n39 = n38 ^ x5 ;
  assign n37 = n10 ^ x5 ;
  assign n40 = n39 ^ n37 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = n41 ^ n34 ;
  assign n43 = n42 ^ n36 ;
  assign n44 = n36 & n43 ;
  assign n45 = n44 ^ n41 ;
  assign n46 = n45 ^ n36 ;
  assign n47 = n10 ^ x6 ;
  assign n48 = n47 ^ n39 ;
  assign n49 = n48 ^ n40 ;
  assign n50 = n49 ^ n10 ;
  assign n51 = n50 ^ n10 ;
  assign n52 = n51 ^ n34 ;
  assign n53 = n50 ^ n40 ;
  assign n57 = n53 ^ n41 ;
  assign n58 = n57 ^ n34 ;
  assign n59 = ~n10 & n58 ;
  assign n54 = n53 ^ n34 ;
  assign n55 = n40 ^ n36 ;
  assign n56 = n54 & n55 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = n60 ^ n40 ;
  assign n62 = n61 ^ n50 ;
  assign n63 = n62 ^ n34 ;
  assign n64 = ~n52 & n63 ;
  assign n65 = n64 ^ n56 ;
  assign n66 = n65 ^ n40 ;
  assign n67 = n66 ^ n50 ;
  assign n68 = n67 ^ n10 ;
  assign n69 = n68 ^ n34 ;
  assign n70 = n46 & ~n69 ;
  assign n71 = n70 ^ x2 ;
  assign n72 = x3 & ~x6 ;
  assign n73 = x5 ^ x4 ;
  assign n74 = n72 & n73 ;
  assign n75 = ~n71 & ~n74 ;
  assign n76 = ~x0 & ~n75 ;
  assign n77 = ~x0 & x3 ;
  assign n78 = n12 & n77 ;
  assign n79 = ~x7 & x8 ;
  assign n80 = x3 ^ x0 ;
  assign n81 = x6 ^ x3 ;
  assign n82 = ~n80 & ~n81 ;
  assign n83 = n79 & ~n82 ;
  assign n84 = ~x5 & n12 ;
  assign n85 = ~x5 & x6 ;
  assign n86 = x5 & ~x6 ;
  assign n87 = ~n85 & ~n86 ;
  assign n88 = ~x0 & ~n87 ;
  assign n89 = ~n84 & ~n88 ;
  assign n90 = n89 ^ x4 ;
  assign n91 = n90 ^ n89 ;
  assign n92 = ~x6 & x7 ;
  assign n93 = x8 & n92 ;
  assign n94 = n93 ^ n89 ;
  assign n95 = ~n91 & ~n94 ;
  assign n96 = n95 ^ n89 ;
  assign n97 = ~n83 & n96 ;
  assign n98 = ~n78 & n97 ;
  assign n99 = ~x2 & ~n98 ;
  assign n100 = x0 & ~x8 ;
  assign n101 = ~x3 & x6 ;
  assign n102 = ~n86 & ~n101 ;
  assign n103 = n100 & ~n102 ;
  assign n104 = ~x3 & x8 ;
  assign n105 = x0 & ~x5 ;
  assign n106 = ~x6 & n105 ;
  assign n107 = ~n104 & ~n106 ;
  assign n108 = n73 & ~n107 ;
  assign n109 = ~n103 & ~n108 ;
  assign n110 = ~x7 & ~n109 ;
  assign n111 = x1 & ~n110 ;
  assign n112 = ~n99 & n111 ;
  assign n113 = n105 ^ x4 ;
  assign n114 = ~x8 & n92 ;
  assign n115 = n114 ^ n113 ;
  assign n116 = n115 ^ n105 ;
  assign n117 = n116 ^ n115 ;
  assign n118 = n92 & n104 ;
  assign n119 = x2 & ~n118 ;
  assign n120 = ~x0 & x7 ;
  assign n121 = x3 & ~x8 ;
  assign n122 = ~n120 & ~n121 ;
  assign n123 = x6 & ~n122 ;
  assign n124 = x0 & n13 ;
  assign n125 = ~n118 & ~n124 ;
  assign n126 = ~n123 & n125 ;
  assign n127 = ~n119 & ~n126 ;
  assign n128 = n127 ^ n115 ;
  assign n129 = n128 ^ n113 ;
  assign n130 = n117 & ~n129 ;
  assign n131 = n130 ^ n127 ;
  assign n132 = x2 & ~x3 ;
  assign n133 = ~n127 & ~n132 ;
  assign n134 = n133 ^ n113 ;
  assign n135 = ~n131 & n134 ;
  assign n136 = n135 ^ n133 ;
  assign n137 = n113 & n136 ;
  assign n138 = n137 ^ n130 ;
  assign n139 = n138 ^ x4 ;
  assign n140 = n139 ^ n127 ;
  assign n141 = n112 & ~n140 ;
  assign n142 = ~n76 & n141 ;
  assign n144 = ~x7 & ~x8 ;
  assign n145 = n132 & ~n144 ;
  assign n143 = x7 ^ x5 ;
  assign n146 = n145 ^ n143 ;
  assign n147 = n145 ^ x7 ;
  assign n148 = n147 ^ x7 ;
  assign n149 = ~x2 & x8 ;
  assign n150 = n149 ^ x7 ;
  assign n151 = ~n148 & n150 ;
  assign n152 = n151 ^ x7 ;
  assign n153 = n146 & n152 ;
  assign n154 = n153 ^ n145 ;
  assign n156 = ~x4 & x5 ;
  assign n157 = x3 & ~x7 ;
  assign n158 = ~x0 & x2 ;
  assign n159 = n157 & n158 ;
  assign n160 = ~n156 & ~n159 ;
  assign n161 = n160 ^ n77 ;
  assign n155 = n77 ^ x2 ;
  assign n162 = n161 ^ n155 ;
  assign n163 = n162 ^ x7 ;
  assign n164 = n163 ^ n161 ;
  assign n165 = n164 ^ n77 ;
  assign n166 = x5 & ~x8 ;
  assign n167 = ~n105 & ~n166 ;
  assign n168 = n167 ^ n163 ;
  assign n169 = ~x7 & ~n168 ;
  assign n170 = n161 ^ n77 ;
  assign n171 = ~n164 & ~n170 ;
  assign n172 = n171 ^ n165 ;
  assign n173 = n169 & n172 ;
  assign n174 = n173 ^ n171 ;
  assign n175 = n165 & n174 ;
  assign n176 = n175 ^ n171 ;
  assign n177 = n176 ^ n160 ;
  assign n178 = ~n154 & n177 ;
  assign n179 = x6 & ~n178 ;
  assign n180 = x5 & x8 ;
  assign n181 = ~n144 & ~n180 ;
  assign n182 = x2 & n181 ;
  assign n183 = ~x4 & n182 ;
  assign n184 = ~x4 & n93 ;
  assign n185 = n79 & n156 ;
  assign n186 = ~n184 & ~n185 ;
  assign n187 = ~n183 & n186 ;
  assign n188 = x3 & ~n187 ;
  assign n189 = ~x1 & ~n188 ;
  assign n190 = ~n179 & n189 ;
  assign n191 = x3 & x7 ;
  assign n192 = n100 & n191 ;
  assign n193 = x0 & ~x3 ;
  assign n194 = ~n92 & ~n193 ;
  assign n195 = n180 & ~n194 ;
  assign n196 = ~n192 & ~n195 ;
  assign n197 = n196 ^ n118 ;
  assign n198 = n197 ^ n196 ;
  assign n199 = ~n12 & ~n86 ;
  assign n200 = x5 & x7 ;
  assign n201 = x0 & ~n200 ;
  assign n202 = ~n199 & n201 ;
  assign n203 = x7 & n156 ;
  assign n204 = ~x3 & n203 ;
  assign n205 = ~n202 & ~n204 ;
  assign n206 = n205 ^ n196 ;
  assign n207 = n206 ^ n196 ;
  assign n208 = ~n198 & n207 ;
  assign n209 = n208 ^ n196 ;
  assign n210 = x2 & n209 ;
  assign n211 = n210 ^ n196 ;
  assign n212 = n190 & n211 ;
  assign n213 = ~n142 & ~n212 ;
  assign n214 = x6 & n144 ;
  assign n215 = n124 & n214 ;
  assign n216 = ~x2 & x7 ;
  assign n217 = n86 & n121 ;
  assign n218 = n216 & n217 ;
  assign n219 = ~n215 & ~n218 ;
  assign n220 = ~n213 & n219 ;
  assign n221 = ~x1 & x5 ;
  assign n222 = ~n77 & ~n79 ;
  assign n223 = n221 & ~n222 ;
  assign n224 = n104 & n120 ;
  assign n225 = n166 & n193 ;
  assign n226 = ~n224 & ~n225 ;
  assign n227 = ~x5 & n191 ;
  assign n228 = ~n17 & ~n227 ;
  assign n229 = ~n72 & ~n101 ;
  assign n230 = ~n157 & n229 ;
  assign n231 = ~n228 & ~n230 ;
  assign n232 = n226 & ~n231 ;
  assign n233 = ~n223 & n232 ;
  assign n234 = ~x2 & ~n233 ;
  assign n235 = x0 & ~x6 ;
  assign n236 = ~n158 & ~n235 ;
  assign n237 = n79 & ~n236 ;
  assign n238 = n92 & n166 ;
  assign n239 = ~n84 & ~n106 ;
  assign n240 = x2 & ~n239 ;
  assign n241 = ~n238 & ~n240 ;
  assign n242 = ~n237 & n241 ;
  assign n243 = ~x3 & ~n242 ;
  assign n244 = ~n234 & ~n243 ;
  assign n245 = n77 & n85 ;
  assign n246 = ~n72 & ~n166 ;
  assign n247 = n158 & ~n246 ;
  assign n248 = ~n14 & n235 ;
  assign n249 = ~n247 & ~n248 ;
  assign n250 = ~n245 & n249 ;
  assign n251 = ~x1 & ~n250 ;
  assign n252 = n221 ^ x8 ;
  assign n253 = n252 ^ x0 ;
  assign n261 = n253 ^ n252 ;
  assign n254 = ~n158 & ~n216 ;
  assign n255 = n254 ^ n253 ;
  assign n256 = n255 ^ n252 ;
  assign n257 = n253 ^ n221 ;
  assign n258 = n257 ^ n254 ;
  assign n259 = n258 ^ n256 ;
  assign n260 = ~n256 & n259 ;
  assign n262 = n261 ^ n260 ;
  assign n263 = n262 ^ n256 ;
  assign n264 = n252 ^ x1 ;
  assign n265 = n260 ^ n256 ;
  assign n266 = ~n264 & ~n265 ;
  assign n267 = n266 ^ n252 ;
  assign n268 = n263 & ~n267 ;
  assign n269 = n268 ^ n252 ;
  assign n270 = n269 ^ x8 ;
  assign n271 = n270 ^ n252 ;
  assign n272 = n101 & ~n271 ;
  assign n273 = ~n251 & ~n272 ;
  assign n274 = x4 & n273 ;
  assign n275 = n244 & n274 ;
  assign n276 = n12 & n13 ;
  assign n277 = ~x5 & ~x7 ;
  assign n278 = n100 & ~n277 ;
  assign n279 = n278 ^ n149 ;
  assign n280 = n279 ^ n193 ;
  assign n281 = n279 ^ n278 ;
  assign n282 = n281 ^ n280 ;
  assign n283 = ~n280 & ~n282 ;
  assign n284 = n283 ^ n279 ;
  assign n285 = n284 ^ n280 ;
  assign n286 = n278 ^ x7 ;
  assign n287 = x3 & ~n286 ;
  assign n288 = n287 ^ n279 ;
  assign n289 = ~n285 & n288 ;
  assign n290 = n289 ^ n279 ;
  assign n291 = n290 ^ n278 ;
  assign n292 = ~n276 & ~n291 ;
  assign n293 = x6 & ~n292 ;
  assign n294 = ~n157 & ~n166 ;
  assign n295 = ~n144 & n235 ;
  assign n296 = ~n294 & n295 ;
  assign n297 = ~n72 & ~n79 ;
  assign n298 = n105 & ~n297 ;
  assign n299 = x2 & n298 ;
  assign n300 = ~n296 & ~n299 ;
  assign n301 = ~n104 & ~n157 ;
  assign n302 = x5 & ~n301 ;
  assign n303 = n158 & n302 ;
  assign n304 = ~x4 & ~n303 ;
  assign n305 = n300 & n304 ;
  assign n306 = ~n293 & n305 ;
  assign n307 = ~n275 & ~n306 ;
  assign n308 = n157 & n166 ;
  assign n309 = ~n118 & ~n308 ;
  assign n310 = x0 & ~n309 ;
  assign n311 = ~x2 & n310 ;
  assign n312 = ~n307 & ~n311 ;
  assign n313 = n220 & n312 ;
  assign y0 = ~n313 ;
endmodule
