module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n18 = x13 & x15 ;
  assign n19 = x11 & ~n18 ;
  assign n20 = x16 & ~n19 ;
  assign n21 = ~x13 & ~x15 ;
  assign n22 = n21 ^ x14 ;
  assign n23 = x1 & x3 ;
  assign n24 = x2 & ~x6 ;
  assign n25 = ~x4 & ~n24 ;
  assign n26 = n23 & n25 ;
  assign n27 = n26 ^ n21 ;
  assign n28 = x14 ^ x11 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = ~n26 & n29 ;
  assign n31 = n30 ^ n26 ;
  assign n32 = ~n27 & ~n31 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ n26 ;
  assign n35 = n34 ^ n28 ;
  assign n36 = n22 & n35 ;
  assign n37 = n36 ^ x11 ;
  assign n38 = ~n20 & n37 ;
  assign y0 = n38 ;
endmodule
