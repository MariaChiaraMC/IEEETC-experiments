// Benchmark "./exp.pla" written by ABC on Thu Apr 23 10:59:51 2020

module \./exp.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z13  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z13;
  assign z13 = x4 | x5;
endmodule


