module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 ;
  assign n9 = x1 & x3 ;
  assign n10 = ~x4 & ~n9 ;
  assign n11 = ~x2 & ~n10 ;
  assign n12 = ~x1 & ~x3 ;
  assign n13 = ~x3 & ~x5 ;
  assign n14 = ~n12 & ~n13 ;
  assign n15 = x6 & n14 ;
  assign n16 = x7 & n15 ;
  assign n17 = ~x1 & ~x5 ;
  assign n18 = x3 & ~n17 ;
  assign n19 = x2 & ~n18 ;
  assign n20 = x4 & ~n12 ;
  assign n21 = n19 & ~n20 ;
  assign n22 = ~n16 & n21 ;
  assign n23 = n22 ^ n11 ;
  assign n25 = ~x3 & ~x7 ;
  assign n26 = ~n17 & ~n25 ;
  assign n27 = ~x6 & ~n26 ;
  assign n28 = n14 & ~n27 ;
  assign n24 = n22 ^ x0 ;
  assign n29 = n28 ^ n24 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = x3 ^ x1 ;
  assign n32 = x5 ^ x3 ;
  assign n33 = n31 & n32 ;
  assign n34 = n33 ^ x3 ;
  assign n35 = n25 ^ n15 ;
  assign n36 = ~n34 & ~n35 ;
  assign n37 = n36 ^ n25 ;
  assign n38 = ~n15 & n37 ;
  assign n39 = n38 ^ n15 ;
  assign n40 = n39 ^ n15 ;
  assign n41 = n40 ^ n28 ;
  assign n42 = ~n30 & ~n41 ;
  assign n43 = n42 ^ n28 ;
  assign n44 = n43 ^ n11 ;
  assign n45 = ~n23 & n44 ;
  assign n46 = n45 ^ n42 ;
  assign n47 = n46 ^ n28 ;
  assign n48 = n47 ^ n22 ;
  assign n49 = n11 & ~n48 ;
  assign n50 = n49 ^ n11 ;
  assign n51 = n50 ^ n24 ;
  assign y0 = n51 ;
endmodule
