module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 ;
  assign n20 = ~x4 & ~x10 ;
  assign n21 = x2 & x3 ;
  assign n22 = ~n20 & n21 ;
  assign n23 = ~x7 & ~x8 ;
  assign n24 = ~n22 & n23 ;
  assign n25 = x9 & n24 ;
  assign n26 = ~x2 & x3 ;
  assign n27 = x7 & ~n26 ;
  assign n13 = x8 & x9 ;
  assign n28 = n13 ^ x4 ;
  assign n29 = n28 ^ n13 ;
  assign n30 = x3 & ~x8 ;
  assign n31 = n30 ^ n13 ;
  assign n32 = n29 & n31 ;
  assign n33 = n32 ^ n13 ;
  assign n34 = n27 & n33 ;
  assign n35 = ~n25 & ~n34 ;
  assign n36 = ~x11 & ~n35 ;
  assign n14 = x4 & ~x10 ;
  assign n15 = x7 & n14 ;
  assign n16 = n13 & n15 ;
  assign n37 = ~x2 & n16 ;
  assign n38 = ~n36 & ~n37 ;
  assign n17 = x2 & ~x3 ;
  assign n18 = ~x11 & n17 ;
  assign n19 = n16 & n18 ;
  assign n39 = n38 ^ n19 ;
  assign n40 = ~x5 & ~n39 ;
  assign n41 = n40 ^ n38 ;
  assign y0 = ~n41 ;
endmodule
