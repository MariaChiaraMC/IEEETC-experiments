module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 ;
  assign n11 = ~x6 & x9 ;
  assign n12 = ~x2 & n11 ;
  assign n13 = x5 & x7 ;
  assign n14 = x1 & x4 ;
  assign n15 = x0 & n14 ;
  assign n16 = n13 & n15 ;
  assign n17 = n16 ^ x7 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = ~x4 & ~x5 ;
  assign n20 = ~x0 & ~x1 ;
  assign n21 = n19 & n20 ;
  assign n22 = n21 ^ n16 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = ~n18 & n23 ;
  assign n25 = n24 ^ n16 ;
  assign n26 = x8 & n25 ;
  assign n27 = n26 ^ n16 ;
  assign n28 = n12 & n27 ;
  assign n29 = ~x5 & x9 ;
  assign n30 = x0 & ~x1 ;
  assign n31 = x6 & ~x7 ;
  assign n32 = ~x8 & n31 ;
  assign n33 = n30 & n32 ;
  assign n34 = x1 & x7 ;
  assign n35 = ~x6 & x8 ;
  assign n36 = n34 & n35 ;
  assign n37 = ~n33 & ~n36 ;
  assign n38 = n29 & ~n37 ;
  assign n39 = ~x0 & ~x5 ;
  assign n40 = x7 & ~x9 ;
  assign n41 = ~x1 & x6 ;
  assign n42 = n40 & n41 ;
  assign n43 = ~x6 & ~x7 ;
  assign n44 = x1 & ~x8 ;
  assign n45 = n43 & n44 ;
  assign n46 = ~n42 & ~n45 ;
  assign n47 = n39 & ~n46 ;
  assign n48 = x1 & x5 ;
  assign n49 = x0 & x5 ;
  assign n50 = ~x6 & ~x9 ;
  assign n51 = n49 & n50 ;
  assign n52 = ~n48 & ~n51 ;
  assign n53 = x1 & ~x9 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = ~x7 & x8 ;
  assign n56 = n55 ^ x0 ;
  assign n57 = n56 ^ n55 ;
  assign n58 = x6 & ~x8 ;
  assign n59 = n58 ^ n55 ;
  assign n60 = ~n57 & n59 ;
  assign n61 = n60 ^ n55 ;
  assign n62 = n61 ^ n52 ;
  assign n63 = n54 & ~n62 ;
  assign n64 = n63 ^ n60 ;
  assign n65 = n64 ^ n55 ;
  assign n66 = n65 ^ n53 ;
  assign n67 = ~n52 & ~n66 ;
  assign n68 = n67 ^ n52 ;
  assign n69 = ~n47 & n68 ;
  assign n70 = ~n38 & n69 ;
  assign n71 = x4 & ~n70 ;
  assign n72 = x7 & x9 ;
  assign n73 = ~x4 & x5 ;
  assign n74 = n41 & n73 ;
  assign n75 = n74 ^ x8 ;
  assign n87 = n75 ^ n74 ;
  assign n76 = n75 ^ x6 ;
  assign n77 = n76 ^ n74 ;
  assign n78 = ~x0 & x1 ;
  assign n79 = n73 & n78 ;
  assign n80 = x0 & x1 ;
  assign n81 = ~x5 & n80 ;
  assign n82 = ~n79 & ~n81 ;
  assign n83 = n82 ^ x6 ;
  assign n84 = n83 ^ x6 ;
  assign n85 = n84 ^ n77 ;
  assign n86 = n77 & ~n85 ;
  assign n88 = n87 ^ n86 ;
  assign n89 = n88 ^ n77 ;
  assign n90 = n74 ^ n19 ;
  assign n91 = n86 ^ n77 ;
  assign n92 = ~n90 & n91 ;
  assign n93 = n92 ^ n74 ;
  assign n94 = n89 & ~n93 ;
  assign n95 = n94 ^ n74 ;
  assign n96 = n95 ^ x8 ;
  assign n97 = n96 ^ n74 ;
  assign n98 = n72 & n97 ;
  assign n99 = x5 & ~x8 ;
  assign n100 = n20 & n40 ;
  assign n101 = n99 & n100 ;
  assign n102 = x6 & n101 ;
  assign n103 = ~n98 & ~n102 ;
  assign n104 = x6 & x9 ;
  assign n105 = ~x0 & ~n104 ;
  assign n106 = ~x4 & ~n105 ;
  assign n107 = ~n50 & ~n106 ;
  assign n108 = ~x5 & ~x7 ;
  assign n109 = x0 & ~n11 ;
  assign n110 = n44 & ~n109 ;
  assign n111 = n108 & n110 ;
  assign n112 = ~n107 & n111 ;
  assign n113 = ~x2 & ~n112 ;
  assign n114 = n103 & n113 ;
  assign n115 = ~n71 & n114 ;
  assign n118 = ~x1 & x4 ;
  assign n119 = ~n20 & ~n118 ;
  assign n120 = n32 & ~n119 ;
  assign n121 = ~x4 & ~x7 ;
  assign n122 = x4 & x7 ;
  assign n123 = ~n121 & ~n122 ;
  assign n124 = x7 & ~x8 ;
  assign n125 = ~x6 & ~n124 ;
  assign n126 = ~n123 & n125 ;
  assign n127 = n78 & n126 ;
  assign n128 = ~n120 & ~n127 ;
  assign n116 = ~x0 & n43 ;
  assign n117 = ~n44 & n116 ;
  assign n129 = n128 ^ n117 ;
  assign n130 = n129 ^ x5 ;
  assign n138 = n130 ^ n129 ;
  assign n131 = x1 & ~x4 ;
  assign n132 = n131 ^ n130 ;
  assign n133 = n132 ^ n129 ;
  assign n134 = n131 ^ n117 ;
  assign n135 = n134 ^ n131 ;
  assign n136 = n135 ^ n133 ;
  assign n137 = ~n133 & ~n136 ;
  assign n139 = n138 ^ n137 ;
  assign n140 = n139 ^ n133 ;
  assign n141 = n129 ^ x8 ;
  assign n142 = n137 ^ n133 ;
  assign n143 = ~n141 & ~n142 ;
  assign n144 = n143 ^ n129 ;
  assign n145 = ~n140 & ~n144 ;
  assign n146 = n145 ^ n129 ;
  assign n147 = n146 ^ n117 ;
  assign n148 = n147 ^ n129 ;
  assign n149 = ~x9 & n148 ;
  assign n171 = n108 & n118 ;
  assign n172 = n11 & n171 ;
  assign n175 = n42 ^ x9 ;
  assign n176 = n175 ^ n42 ;
  assign n173 = n43 ^ n42 ;
  assign n174 = n173 ^ n42 ;
  assign n177 = n176 ^ n174 ;
  assign n178 = n131 ^ n42 ;
  assign n179 = n178 ^ n42 ;
  assign n180 = n179 ^ n176 ;
  assign n181 = n176 & n180 ;
  assign n182 = n181 ^ n176 ;
  assign n183 = ~n177 & n182 ;
  assign n184 = n183 ^ n181 ;
  assign n185 = n184 ^ n42 ;
  assign n186 = n185 ^ n176 ;
  assign n187 = x5 & n186 ;
  assign n188 = n187 ^ n42 ;
  assign n189 = ~n172 & ~n188 ;
  assign n150 = x6 & x7 ;
  assign n151 = n150 ^ x5 ;
  assign n152 = n151 ^ x4 ;
  assign n161 = n152 ^ n150 ;
  assign n153 = n150 ^ x9 ;
  assign n154 = n153 ^ n152 ;
  assign n155 = n154 ^ n152 ;
  assign n156 = n155 ^ n150 ;
  assign n157 = n154 ^ x4 ;
  assign n158 = n157 ^ n154 ;
  assign n159 = n158 ^ n156 ;
  assign n160 = n156 & n159 ;
  assign n162 = n161 ^ n160 ;
  assign n163 = n162 ^ n156 ;
  assign n164 = n150 ^ n43 ;
  assign n165 = n160 ^ n156 ;
  assign n166 = n164 & n165 ;
  assign n167 = n166 ^ n150 ;
  assign n168 = n163 & n167 ;
  assign n169 = n168 ^ n150 ;
  assign n170 = n169 ^ n150 ;
  assign n190 = n189 ^ n170 ;
  assign n191 = n190 ^ n189 ;
  assign n192 = n189 ^ x1 ;
  assign n193 = n192 ^ n189 ;
  assign n194 = n191 & n193 ;
  assign n195 = n194 ^ n189 ;
  assign n196 = ~x8 & ~n195 ;
  assign n197 = n196 ^ n189 ;
  assign n198 = n197 ^ x0 ;
  assign n199 = n198 ^ n197 ;
  assign n200 = n199 ^ x2 ;
  assign n201 = ~x4 & ~x6 ;
  assign n202 = n29 & n34 ;
  assign n203 = n202 ^ n201 ;
  assign n204 = n201 & n203 ;
  assign n205 = n204 ^ n197 ;
  assign n206 = n205 ^ n201 ;
  assign n207 = ~n200 & ~n206 ;
  assign n208 = n207 ^ n204 ;
  assign n209 = n208 ^ n201 ;
  assign n210 = x2 & n209 ;
  assign n211 = n210 ^ x2 ;
  assign n212 = ~n149 & n211 ;
  assign n213 = ~n115 & ~n212 ;
  assign n214 = n213 ^ x3 ;
  assign n215 = n214 ^ n213 ;
  assign n216 = n215 ^ n28 ;
  assign n217 = n15 & n104 ;
  assign n218 = ~x2 & n217 ;
  assign n219 = x6 ^ x2 ;
  assign n220 = n219 ^ x9 ;
  assign n221 = x1 ^ x0 ;
  assign n222 = n221 ^ x2 ;
  assign n223 = n222 ^ n220 ;
  assign n224 = x9 ^ x6 ;
  assign n225 = x6 ^ x1 ;
  assign n226 = n225 ^ x6 ;
  assign n227 = ~n224 & n226 ;
  assign n228 = n227 ^ x6 ;
  assign n229 = n228 ^ n220 ;
  assign n230 = ~n223 & n229 ;
  assign n231 = n230 ^ n227 ;
  assign n232 = n231 ^ x6 ;
  assign n233 = n232 ^ n222 ;
  assign n234 = n220 & ~n233 ;
  assign n235 = n234 ^ n220 ;
  assign n236 = n121 & n235 ;
  assign n237 = ~x5 & ~x8 ;
  assign n238 = ~n236 & n237 ;
  assign n239 = ~n218 & n238 ;
  assign n240 = x2 & x4 ;
  assign n241 = n72 & n240 ;
  assign n242 = n41 & n241 ;
  assign n243 = n99 & ~n242 ;
  assign n244 = ~n31 & ~n122 ;
  assign n245 = ~x2 & ~n201 ;
  assign n246 = x0 & n245 ;
  assign n247 = n244 & n246 ;
  assign n248 = x2 & ~x4 ;
  assign n249 = n116 & n248 ;
  assign n250 = ~n247 & ~n249 ;
  assign n251 = ~x1 & ~x9 ;
  assign n252 = ~n250 & n251 ;
  assign n253 = n243 & ~n252 ;
  assign n254 = x6 ^ x4 ;
  assign n255 = ~x7 & n254 ;
  assign n256 = ~x2 & n255 ;
  assign n257 = n256 ^ x0 ;
  assign n258 = n257 ^ n256 ;
  assign n259 = n258 ^ n53 ;
  assign n260 = n31 & n240 ;
  assign n261 = ~x2 & n201 ;
  assign n262 = n261 ^ n260 ;
  assign n263 = ~n260 & n262 ;
  assign n264 = n263 ^ n256 ;
  assign n265 = n264 ^ n260 ;
  assign n266 = n259 & n265 ;
  assign n267 = n266 ^ n263 ;
  assign n268 = n267 ^ n260 ;
  assign n269 = n53 & ~n268 ;
  assign n270 = n269 ^ n53 ;
  assign n271 = n253 & ~n270 ;
  assign n272 = ~n239 & ~n271 ;
  assign n273 = ~x2 & n118 ;
  assign n274 = ~n80 & ~n273 ;
  assign n275 = x5 & ~x6 ;
  assign n276 = ~n274 & n275 ;
  assign n277 = n276 ^ n248 ;
  assign n278 = n277 ^ n276 ;
  assign n279 = n39 ^ x6 ;
  assign n280 = n279 ^ n39 ;
  assign n281 = n49 ^ n39 ;
  assign n282 = n281 ^ n39 ;
  assign n283 = n280 & n282 ;
  assign n284 = n283 ^ n39 ;
  assign n285 = ~n225 & n284 ;
  assign n286 = n285 ^ n39 ;
  assign n287 = n286 ^ n276 ;
  assign n288 = n278 & n287 ;
  assign n289 = n288 ^ n276 ;
  assign n290 = n40 & n289 ;
  assign n291 = x8 & ~n290 ;
  assign n292 = ~x2 & n43 ;
  assign n293 = n21 & n292 ;
  assign n294 = n291 & ~n293 ;
  assign n343 = x0 & x2 ;
  assign n295 = ~n49 & ~n108 ;
  assign n296 = n108 & n240 ;
  assign n297 = n296 ^ n261 ;
  assign n298 = n297 ^ n261 ;
  assign n299 = n261 ^ x0 ;
  assign n300 = n299 ^ n261 ;
  assign n301 = n298 & n300 ;
  assign n302 = n301 ^ n261 ;
  assign n303 = x1 & n302 ;
  assign n304 = n303 ^ n261 ;
  assign n305 = ~n295 & n304 ;
  assign n306 = n31 & n73 ;
  assign n307 = n20 & n306 ;
  assign n308 = x1 & x6 ;
  assign n309 = n308 ^ n123 ;
  assign n310 = x5 ^ x0 ;
  assign n311 = n310 ^ x5 ;
  assign n312 = n108 ^ x5 ;
  assign n313 = ~n311 & n312 ;
  assign n314 = n313 ^ x5 ;
  assign n315 = n314 ^ n308 ;
  assign n316 = ~n309 & n315 ;
  assign n317 = n316 ^ n313 ;
  assign n318 = n317 ^ x5 ;
  assign n319 = n318 ^ n123 ;
  assign n320 = n308 & ~n319 ;
  assign n321 = n320 ^ n308 ;
  assign n322 = ~n307 & ~n321 ;
  assign n323 = n322 ^ x2 ;
  assign n324 = n323 ^ n322 ;
  assign n325 = n19 & n31 ;
  assign n326 = x7 ^ x5 ;
  assign n327 = n326 ^ x7 ;
  assign n328 = n150 ^ x7 ;
  assign n329 = ~n327 & ~n328 ;
  assign n330 = n329 ^ x7 ;
  assign n331 = x4 & ~n330 ;
  assign n332 = ~n325 & ~n331 ;
  assign n333 = n20 & ~n332 ;
  assign n334 = ~x0 & n13 ;
  assign n335 = n308 & n334 ;
  assign n336 = ~n333 & ~n335 ;
  assign n337 = n336 ^ n322 ;
  assign n338 = n324 & n337 ;
  assign n339 = n338 ^ n322 ;
  assign n340 = ~n305 & n339 ;
  assign n344 = n343 ^ n340 ;
  assign n345 = n344 ^ n340 ;
  assign n341 = n340 ^ n325 ;
  assign n342 = n341 ^ n340 ;
  assign n346 = n345 ^ n342 ;
  assign n347 = n340 ^ x1 ;
  assign n348 = n347 ^ n340 ;
  assign n349 = n348 ^ n345 ;
  assign n350 = n345 & n349 ;
  assign n351 = n350 ^ n345 ;
  assign n352 = n346 & n351 ;
  assign n353 = n352 ^ n350 ;
  assign n354 = n353 ^ n340 ;
  assign n355 = n354 ^ n345 ;
  assign n356 = ~x9 & ~n355 ;
  assign n357 = n356 ^ n340 ;
  assign n358 = n294 & n357 ;
  assign n359 = n358 ^ n272 ;
  assign n360 = n272 & ~n359 ;
  assign n361 = n360 ^ n213 ;
  assign n362 = n361 ^ n272 ;
  assign n363 = n216 & n362 ;
  assign n364 = n363 ^ n360 ;
  assign n365 = n364 ^ n272 ;
  assign n366 = ~n28 & n365 ;
  assign n367 = n366 ^ n28 ;
  assign y0 = n367 ;
endmodule
