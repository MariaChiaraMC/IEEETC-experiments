module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 ;
  assign n20 = x9 & ~x14 ;
  assign n21 = ~x8 & x18 ;
  assign n22 = x7 & x17 ;
  assign n23 = ~x7 & ~x17 ;
  assign n24 = ~n22 & ~n23 ;
  assign n25 = n21 & ~n24 ;
  assign n26 = x8 & ~x18 ;
  assign n27 = x17 & n26 ;
  assign n28 = ~x7 & n27 ;
  assign n29 = ~n25 & ~n28 ;
  assign n30 = n20 & ~n29 ;
  assign n31 = ~n21 & ~n26 ;
  assign n32 = ~n24 & n31 ;
  assign n33 = ~x9 & n32 ;
  assign n34 = ~n30 & ~n33 ;
  assign n49 = x4 & ~n34 ;
  assign n39 = ~x17 & ~x18 ;
  assign n50 = ~n30 & n39 ;
  assign n51 = ~x6 & ~n50 ;
  assign n52 = n49 & n51 ;
  assign n68 = x6 & ~n39 ;
  assign n53 = x1 & x3 ;
  assign n54 = ~x5 & n53 ;
  assign n55 = x12 ^ x11 ;
  assign n56 = x13 ^ x11 ;
  assign n57 = n39 ^ x11 ;
  assign n58 = x11 & n57 ;
  assign n59 = n58 ^ x11 ;
  assign n60 = ~n56 & n59 ;
  assign n61 = n60 ^ n58 ;
  assign n62 = n61 ^ x11 ;
  assign n63 = n62 ^ n39 ;
  assign n64 = ~n55 & n63 ;
  assign n65 = n64 ^ n39 ;
  assign n66 = n54 & n65 ;
  assign n67 = ~x10 & n66 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = ~x14 & n69 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = ~n52 & ~n71 ;
  assign n35 = n34 ^ x6 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = n36 ^ x4 ;
  assign n38 = x7 & x8 ;
  assign n40 = n38 & n39 ;
  assign n41 = n40 ^ x4 ;
  assign n42 = n20 & ~n41 ;
  assign n43 = n42 ^ n34 ;
  assign n44 = ~n37 & ~n43 ;
  assign n45 = n44 ^ n42 ;
  assign n46 = ~x4 & n45 ;
  assign n47 = n46 ^ n42 ;
  assign n48 = n47 ^ n44 ;
  assign n73 = n72 ^ n48 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = ~x6 & n38 ;
  assign n76 = x14 & ~n68 ;
  assign n77 = ~n75 & n76 ;
  assign n78 = n77 ^ n72 ;
  assign n79 = n78 ^ n72 ;
  assign n80 = ~n74 & ~n79 ;
  assign n81 = n80 ^ n72 ;
  assign n82 = x16 & n81 ;
  assign n83 = n82 ^ n72 ;
  assign n84 = x18 ^ x8 ;
  assign n85 = x17 ^ x7 ;
  assign n86 = n85 ^ x18 ;
  assign n87 = n84 & n86 ;
  assign n88 = n87 ^ x14 ;
  assign n89 = n39 & n88 ;
  assign n90 = n89 ^ n87 ;
  assign n91 = x14 & n90 ;
  assign n92 = n91 ^ x14 ;
  assign n93 = n83 & ~n92 ;
  assign y0 = ~n93 ;
endmodule
