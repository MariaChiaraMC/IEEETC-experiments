module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 ;
  output y0 ;
  wire n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 ;
  assign n24 = x2 ^ x1 ;
  assign n25 = x1 ^ x0 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = x3 ^ x2 ;
  assign n28 = x5 ^ x2 ;
  assign n29 = n27 & ~n28 ;
  assign n30 = n29 ^ x2 ;
  assign n31 = n30 ^ n24 ;
  assign n32 = n26 & ~n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ x2 ;
  assign n35 = n34 ^ n25 ;
  assign n36 = n24 & ~n35 ;
  assign n37 = n36 ^ n24 ;
  assign n38 = ~x4 & n37 ;
  assign n39 = x19 ^ x18 ;
  assign n40 = n39 ^ x18 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = x2 & x4 ;
  assign n43 = x0 & ~x1 ;
  assign n44 = ~x9 & ~x10 ;
  assign n45 = x8 & x11 ;
  assign n46 = ~x6 & n45 ;
  assign n47 = ~n44 & n46 ;
  assign n48 = ~x6 & ~x7 ;
  assign n49 = x8 & ~x10 ;
  assign n50 = n48 & n49 ;
  assign n51 = ~x11 & n50 ;
  assign n52 = ~n47 & ~n51 ;
  assign n53 = ~x10 & ~x13 ;
  assign n54 = x10 & ~x11 ;
  assign n55 = ~x8 & n54 ;
  assign n56 = x9 & ~n55 ;
  assign n57 = ~n53 & n56 ;
  assign n58 = n52 & ~n57 ;
  assign n59 = ~x15 & ~n58 ;
  assign n60 = ~x8 & n48 ;
  assign n61 = x11 & ~x16 ;
  assign n62 = x10 & ~x13 ;
  assign n63 = ~n61 & ~n62 ;
  assign n64 = n60 & ~n63 ;
  assign n65 = x10 & x11 ;
  assign n66 = ~x15 & ~n65 ;
  assign n67 = n64 & n66 ;
  assign n68 = x7 & ~n44 ;
  assign n69 = ~x13 & n68 ;
  assign n70 = n45 & n69 ;
  assign n71 = ~n67 & ~n70 ;
  assign n72 = n71 ^ x9 ;
  assign n73 = n72 ^ n71 ;
  assign n76 = ~x8 & ~x11 ;
  assign n74 = n48 & n53 ;
  assign n75 = n74 ^ n68 ;
  assign n77 = n76 ^ n75 ;
  assign n85 = n77 ^ n75 ;
  assign n78 = n46 & n53 ;
  assign n79 = n78 ^ n77 ;
  assign n80 = n79 ^ n75 ;
  assign n81 = n77 ^ n74 ;
  assign n82 = n81 ^ n78 ;
  assign n83 = n82 ^ n80 ;
  assign n84 = ~n80 & ~n83 ;
  assign n86 = n85 ^ n84 ;
  assign n87 = n86 ^ n80 ;
  assign n88 = x6 & ~n49 ;
  assign n89 = n88 ^ n75 ;
  assign n90 = n84 ^ n80 ;
  assign n91 = ~n89 & ~n90 ;
  assign n92 = n91 ^ n75 ;
  assign n93 = ~n87 & n92 ;
  assign n94 = n93 ^ n75 ;
  assign n95 = n94 ^ n68 ;
  assign n96 = n95 ^ n75 ;
  assign n97 = n96 ^ n71 ;
  assign n98 = n73 & ~n97 ;
  assign n99 = n98 ^ n71 ;
  assign n100 = ~n59 & n99 ;
  assign n101 = ~x12 & ~n100 ;
  assign n102 = x13 & ~x15 ;
  assign n103 = n44 ^ x16 ;
  assign n104 = ~x11 & ~n103 ;
  assign n105 = n104 ^ x16 ;
  assign n106 = n102 & ~n105 ;
  assign n107 = x6 & x13 ;
  assign n108 = ~n106 & ~n107 ;
  assign n109 = ~n101 & n108 ;
  assign n110 = ~x17 & n109 ;
  assign n111 = ~x1 & ~n110 ;
  assign n112 = x16 & n48 ;
  assign n113 = n112 ^ x10 ;
  assign n114 = n113 ^ n112 ;
  assign n115 = ~x1 & ~x15 ;
  assign n116 = n115 ^ n112 ;
  assign n117 = n116 ^ n112 ;
  assign n118 = n114 & n117 ;
  assign n119 = n118 ^ n112 ;
  assign n120 = x13 & n119 ;
  assign n121 = n120 ^ n112 ;
  assign n122 = x12 & n121 ;
  assign n123 = ~x8 & n44 ;
  assign n124 = x7 & x13 ;
  assign n125 = ~x12 & n124 ;
  assign n126 = n125 ^ n102 ;
  assign n127 = n123 & n126 ;
  assign n128 = n127 ^ n102 ;
  assign n129 = x11 & n128 ;
  assign n130 = ~x12 & ~x13 ;
  assign n131 = ~x9 & n130 ;
  assign n132 = ~x6 & x8 ;
  assign n133 = n131 & n132 ;
  assign n134 = n65 & n133 ;
  assign n135 = ~x1 & ~n134 ;
  assign n136 = ~n129 & n135 ;
  assign n137 = x16 & ~n136 ;
  assign n138 = ~n122 & ~n137 ;
  assign n139 = ~n111 & n138 ;
  assign n140 = x5 & ~n139 ;
  assign n141 = ~n43 & ~n140 ;
  assign n142 = n42 & ~n141 ;
  assign n143 = x0 & x2 ;
  assign n144 = ~x4 & x5 ;
  assign n145 = ~x21 & n144 ;
  assign n146 = x8 & n54 ;
  assign n147 = n48 & ~n65 ;
  assign n148 = x11 ^ x8 ;
  assign n149 = n147 & ~n148 ;
  assign n150 = ~n146 & ~n149 ;
  assign n151 = x9 & ~n150 ;
  assign n152 = n54 & n60 ;
  assign n153 = ~n151 & ~n152 ;
  assign n154 = n130 & ~n153 ;
  assign n155 = ~x1 & n154 ;
  assign n156 = ~n145 & ~n155 ;
  assign n157 = n143 & ~n156 ;
  assign n158 = ~x21 & x22 ;
  assign n159 = ~x2 & n158 ;
  assign n160 = x9 & ~x12 ;
  assign n161 = ~x13 & n160 ;
  assign n162 = x1 & n161 ;
  assign n163 = ~n150 & n162 ;
  assign n164 = ~n159 & ~n163 ;
  assign n165 = ~x4 & ~x5 ;
  assign n166 = ~x0 & n165 ;
  assign n167 = ~n164 & n166 ;
  assign n168 = n65 & n160 ;
  assign n169 = x0 & ~x13 ;
  assign n170 = ~n168 & n169 ;
  assign n171 = x1 & x5 ;
  assign n172 = ~n143 & n171 ;
  assign n173 = ~n170 & n172 ;
  assign n174 = ~n144 & ~n173 ;
  assign n175 = n43 ^ x15 ;
  assign n176 = n175 ^ x4 ;
  assign n183 = n176 ^ n175 ;
  assign n177 = n176 ^ x0 ;
  assign n178 = n177 ^ n175 ;
  assign n179 = n176 ^ n43 ;
  assign n180 = n179 ^ x0 ;
  assign n181 = n180 ^ n178 ;
  assign n182 = ~n178 & n181 ;
  assign n184 = n183 ^ n182 ;
  assign n185 = n184 ^ n178 ;
  assign n186 = n175 ^ x12 ;
  assign n187 = n182 ^ n178 ;
  assign n188 = n186 & ~n187 ;
  assign n189 = n188 ^ n175 ;
  assign n190 = n185 & n189 ;
  assign n191 = n190 ^ n175 ;
  assign n192 = n191 ^ x15 ;
  assign n193 = n192 ^ n175 ;
  assign n194 = ~n174 & n193 ;
  assign n195 = ~n167 & ~n194 ;
  assign n196 = ~n157 & n195 ;
  assign n197 = ~x3 & n196 ;
  assign n198 = ~n142 & n197 ;
  assign n199 = ~x22 & n143 ;
  assign n200 = ~n43 & ~n199 ;
  assign n201 = n149 & n161 ;
  assign n202 = ~x2 & n201 ;
  assign n203 = ~x4 & ~n202 ;
  assign n204 = ~n200 & ~n203 ;
  assign n205 = n204 ^ x5 ;
  assign n206 = n205 ^ n204 ;
  assign n207 = n206 ^ x3 ;
  assign n208 = x4 & ~n115 ;
  assign n209 = n131 ^ n60 ;
  assign n210 = x11 ^ x10 ;
  assign n211 = n210 ^ x11 ;
  assign n212 = x11 & x15 ;
  assign n213 = n212 ^ x11 ;
  assign n214 = ~n211 & ~n213 ;
  assign n215 = n214 ^ x11 ;
  assign n216 = n215 ^ n131 ;
  assign n217 = n209 & ~n216 ;
  assign n218 = n217 ^ n214 ;
  assign n219 = n218 ^ x11 ;
  assign n220 = n219 ^ n60 ;
  assign n221 = n131 & ~n220 ;
  assign n222 = n221 ^ n131 ;
  assign n223 = n222 ^ x0 ;
  assign n224 = n222 ^ x2 ;
  assign n225 = n222 & ~n224 ;
  assign n226 = n225 ^ n222 ;
  assign n227 = n223 & n226 ;
  assign n228 = n227 ^ n225 ;
  assign n229 = n228 ^ n222 ;
  assign n230 = n229 ^ x2 ;
  assign n231 = ~n25 & ~n230 ;
  assign n232 = n231 ^ x1 ;
  assign n233 = n232 ^ n208 ;
  assign n234 = ~n208 & ~n233 ;
  assign n235 = n234 ^ n204 ;
  assign n236 = n235 ^ n208 ;
  assign n237 = n207 & ~n236 ;
  assign n238 = n237 ^ n234 ;
  assign n239 = n238 ^ n208 ;
  assign n240 = x3 & ~n239 ;
  assign n241 = n240 ^ x3 ;
  assign n242 = ~n198 & ~n241 ;
  assign n243 = n42 & n171 ;
  assign n244 = ~x0 & n243 ;
  assign n245 = ~n242 & ~n244 ;
  assign n246 = n245 ^ x20 ;
  assign n247 = ~x20 & n246 ;
  assign n248 = n247 ^ x18 ;
  assign n249 = n248 ^ x20 ;
  assign n250 = n41 & n249 ;
  assign n251 = n250 ^ n247 ;
  assign n252 = n251 ^ x20 ;
  assign n253 = ~n38 & ~n252 ;
  assign n254 = n253 ^ n38 ;
  assign n255 = x14 & n254 ;
  assign y0 = n255 ;
endmodule
