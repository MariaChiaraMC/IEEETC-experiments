module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 ;
  assign n9 = ~x3 & ~x4 ;
  assign n8 = x2 ^ x1 ;
  assign n10 = n9 ^ n8 ;
  assign n12 = n10 ^ n9 ;
  assign n11 = n10 ^ x2 ;
  assign n13 = n12 ^ n11 ;
  assign n20 = n13 ^ n10 ;
  assign n21 = n20 ^ n12 ;
  assign n22 = n21 ^ n12 ;
  assign n14 = ~x5 & ~x6 ;
  assign n23 = x0 & n14 ;
  assign n24 = ~x3 & ~n23 ;
  assign n25 = n24 ^ n10 ;
  assign n26 = n25 ^ n12 ;
  assign n27 = ~n22 & n26 ;
  assign n15 = n14 ^ n10 ;
  assign n16 = n15 ^ n10 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n17 ^ n12 ;
  assign n19 = n13 & ~n18 ;
  assign n28 = n27 ^ n19 ;
  assign n29 = n28 ^ n13 ;
  assign n30 = n19 ^ n12 ;
  assign n31 = n30 ^ n21 ;
  assign n32 = n12 & ~n31 ;
  assign n33 = n32 ^ n19 ;
  assign n34 = n29 & n33 ;
  assign n35 = n34 ^ n27 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ n13 ;
  assign n38 = n37 ^ n12 ;
  assign n39 = n38 ^ n21 ;
  assign n40 = n39 ^ x1 ;
  assign y0 = ~n40 ;
endmodule
