module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ;
  assign n15 = x10 & ~x12 ;
  assign n16 = ~x9 & ~n15 ;
  assign n17 = x11 & ~n16 ;
  assign n18 = x10 ^ x9 ;
  assign n19 = n18 ^ x13 ;
  assign n20 = n19 ^ x9 ;
  assign n21 = n20 ^ x7 ;
  assign n22 = x13 ^ x12 ;
  assign n23 = ~x11 & ~n22 ;
  assign n24 = n23 ^ x13 ;
  assign n25 = n24 ^ n20 ;
  assign n26 = ~x9 & n25 ;
  assign n27 = n26 ^ x13 ;
  assign n28 = n27 ^ x9 ;
  assign n29 = n28 ^ n20 ;
  assign n30 = n29 ^ x7 ;
  assign n31 = ~n21 & ~n30 ;
  assign n32 = n31 ^ n26 ;
  assign n33 = n32 ^ x13 ;
  assign n34 = n33 ^ n20 ;
  assign n35 = x7 & n34 ;
  assign n36 = n35 ^ x7 ;
  assign n37 = n36 ^ x7 ;
  assign n38 = n37 ^ x7 ;
  assign n39 = ~n17 & n38 ;
  assign y0 = n39 ;
endmodule
