module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 ;
  assign n84 = x3 & ~x5 ;
  assign n103 = ~x1 & x8 ;
  assign n104 = x6 & ~x13 ;
  assign n105 = n103 & n104 ;
  assign n106 = n84 & n105 ;
  assign n53 = ~x13 & ~x14 ;
  assign n54 = x3 & n53 ;
  assign n55 = ~x7 & ~x10 ;
  assign n56 = ~x2 & ~x4 ;
  assign n57 = n55 & n56 ;
  assign n58 = n54 & n57 ;
  assign n59 = ~x6 & n58 ;
  assign n60 = x2 & x4 ;
  assign n61 = x10 & n60 ;
  assign n62 = x14 ^ x13 ;
  assign n63 = x13 ^ x3 ;
  assign n64 = n63 ^ n62 ;
  assign n65 = x6 & ~x7 ;
  assign n66 = n65 ^ x14 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = ~x6 & x11 ;
  assign n69 = n68 ^ n65 ;
  assign n70 = n67 & n69 ;
  assign n71 = n70 ^ n65 ;
  assign n72 = n71 ^ n62 ;
  assign n73 = ~n64 & ~n72 ;
  assign n74 = n73 ^ n70 ;
  assign n75 = n74 ^ n65 ;
  assign n76 = n75 ^ n63 ;
  assign n77 = ~n62 & n76 ;
  assign n78 = n77 ^ n62 ;
  assign n79 = n61 & ~n78 ;
  assign n80 = ~n59 & ~n79 ;
  assign n81 = ~x8 & ~x15 ;
  assign n82 = x5 & n81 ;
  assign n83 = ~n80 & n82 ;
  assign n85 = x15 & ~n84 ;
  assign n86 = x8 & n56 ;
  assign n87 = n53 & n65 ;
  assign n88 = n86 & n87 ;
  assign n89 = n85 & n88 ;
  assign n90 = x10 & n89 ;
  assign n91 = ~n83 & ~n90 ;
  assign n17 = ~x14 & ~x15 ;
  assign n18 = x6 & n17 ;
  assign n19 = ~x5 & n18 ;
  assign n20 = x8 ^ x1 ;
  assign n21 = ~x2 & ~n20 ;
  assign n22 = n19 & n21 ;
  assign n23 = x4 & ~x13 ;
  assign n24 = x7 & x10 ;
  assign n25 = n23 & n24 ;
  assign n26 = x3 & n25 ;
  assign n27 = n22 & n26 ;
  assign n92 = n91 ^ n27 ;
  assign n28 = ~x8 & n23 ;
  assign n29 = x5 & x7 ;
  assign n30 = x14 & ~n29 ;
  assign n31 = x10 ^ x7 ;
  assign n32 = x6 & n31 ;
  assign n33 = n30 & ~n32 ;
  assign n36 = n33 ^ n19 ;
  assign n37 = n36 ^ n33 ;
  assign n34 = n33 ^ x10 ;
  assign n35 = n34 ^ n33 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = n33 ^ x7 ;
  assign n40 = n39 ^ n33 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n37 & n41 ;
  assign n43 = n42 ^ n37 ;
  assign n44 = ~n38 & n43 ;
  assign n45 = n44 ^ n42 ;
  assign n46 = n45 ^ n33 ;
  assign n47 = n46 ^ n37 ;
  assign n48 = ~x2 & n47 ;
  assign n49 = n48 ^ n33 ;
  assign n50 = x3 & n49 ;
  assign n51 = n28 & n50 ;
  assign n52 = n51 ^ n27 ;
  assign n93 = n92 ^ n52 ;
  assign n94 = n92 ^ x1 ;
  assign n95 = n94 ^ n92 ;
  assign n96 = ~n93 & n95 ;
  assign n97 = n96 ^ n92 ;
  assign n98 = x9 & ~n97 ;
  assign n99 = n98 ^ n27 ;
  assign n107 = n106 ^ n99 ;
  assign n108 = n107 ^ n99 ;
  assign n100 = x7 & x9 ;
  assign n101 = n100 ^ n99 ;
  assign n102 = n101 ^ n99 ;
  assign n109 = n108 ^ n102 ;
  assign n110 = n17 & n60 ;
  assign n111 = n110 ^ n99 ;
  assign n112 = n111 ^ n99 ;
  assign n113 = n112 ^ n108 ;
  assign n114 = n108 & n113 ;
  assign n115 = n114 ^ n108 ;
  assign n116 = n109 & n115 ;
  assign n117 = n116 ^ n114 ;
  assign n118 = n117 ^ n99 ;
  assign n119 = n118 ^ n108 ;
  assign n120 = x0 & n119 ;
  assign n121 = n120 ^ n99 ;
  assign n122 = ~x12 & n121 ;
  assign y0 = n122 ;
endmodule
