module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n8 = x1 & ~x4 ;
  assign n7 = ~x0 & x2 ;
  assign n9 = n8 ^ n7 ;
  assign n10 = n9 ^ x5 ;
  assign n11 = n10 ^ n7 ;
  assign n12 = n11 ^ x3 ;
  assign n13 = ~x1 & x4 ;
  assign n14 = x0 & ~x2 ;
  assign n15 = ~n13 & n14 ;
  assign n16 = n15 ^ x5 ;
  assign n17 = n15 & ~n16 ;
  assign n18 = n17 ^ n7 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n12 & n19 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n21 ^ n15 ;
  assign n23 = ~x3 & n22 ;
  assign n24 = ~x4 & ~x5 ;
  assign n25 = x3 & ~n24 ;
  assign n26 = ~x1 & ~x5 ;
  assign n27 = x1 ^ x0 ;
  assign n28 = x2 ^ x1 ;
  assign n29 = ~n27 & ~n28 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = n26 & n30 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = n25 & n32 ;
  assign n34 = ~n23 & ~n33 ;
  assign y0 = ~n34 ;
endmodule
