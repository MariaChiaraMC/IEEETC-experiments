module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 ;
  assign n13 = x8 & x9 ;
  assign n14 = ~x5 & n13 ;
  assign n15 = x3 & x4 ;
  assign n16 = x2 & n15 ;
  assign n17 = n14 & n16 ;
  assign n18 = x10 & ~x11 ;
  assign n19 = x6 & n18 ;
  assign n20 = n17 & n19 ;
  assign n21 = x7 & n20 ;
  assign n22 = x5 & ~x6 ;
  assign n23 = ~x3 & ~x4 ;
  assign n24 = ~x2 & x7 ;
  assign n25 = n13 & n24 ;
  assign n26 = n23 & n25 ;
  assign n27 = x10 & n26 ;
  assign n28 = n27 ^ x11 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ n22 ;
  assign n31 = n15 ^ x9 ;
  assign n32 = n31 ^ n15 ;
  assign n33 = x3 & ~x4 ;
  assign n34 = n33 ^ n15 ;
  assign n35 = n34 ^ n15 ;
  assign n36 = n32 & n35 ;
  assign n37 = n36 ^ n15 ;
  assign n38 = x8 & n37 ;
  assign n39 = n38 ^ n15 ;
  assign n40 = n39 ^ x2 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = n41 ^ x7 ;
  assign n43 = ~x10 & n13 ;
  assign n44 = n43 ^ n33 ;
  assign n45 = ~n33 & ~n44 ;
  assign n46 = n45 ^ n39 ;
  assign n47 = n46 ^ n33 ;
  assign n48 = ~n42 & ~n47 ;
  assign n49 = n48 ^ n45 ;
  assign n50 = n49 ^ n33 ;
  assign n51 = x7 & ~n50 ;
  assign n52 = ~x2 & n15 ;
  assign n53 = ~n23 & ~n52 ;
  assign n54 = ~x7 & ~x8 ;
  assign n55 = x9 & n54 ;
  assign n56 = ~n53 & n55 ;
  assign n57 = n56 ^ n51 ;
  assign n58 = ~n51 & n57 ;
  assign n59 = n58 ^ n27 ;
  assign n60 = n59 ^ n51 ;
  assign n61 = ~n30 & n60 ;
  assign n62 = n61 ^ n58 ;
  assign n63 = n62 ^ n51 ;
  assign n64 = n22 & ~n63 ;
  assign n65 = n64 ^ n22 ;
  assign n66 = ~n21 & ~n65 ;
  assign n67 = x0 & ~n66 ;
  assign n68 = x1 & n67 ;
  assign y0 = n68 ;
endmodule
