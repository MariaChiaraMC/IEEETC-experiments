module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n9 = x7 ^ x5 ;
  assign n10 = x5 ^ x3 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = x1 & ~x2 ;
  assign n13 = x0 & x6 ;
  assign n14 = n12 & n13 ;
  assign n15 = n14 ^ x7 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = ~x1 & x2 ;
  assign n18 = ~x0 & ~x6 ;
  assign n19 = n17 & n18 ;
  assign n20 = n19 ^ n14 ;
  assign n21 = n16 & n20 ;
  assign n22 = n21 ^ n14 ;
  assign n23 = n22 ^ n9 ;
  assign n24 = n11 & ~n23 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ n14 ;
  assign n27 = n26 ^ n10 ;
  assign n28 = ~n9 & ~n27 ;
  assign n29 = n28 ^ n9 ;
  assign n30 = ~x4 & ~n29 ;
  assign y0 = n30 ;
endmodule
