module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 ;
  assign n11 = x1 & x7 ;
  assign n12 = x2 & n11 ;
  assign n13 = ~x3 & x7 ;
  assign n14 = ~x0 & n13 ;
  assign n15 = x1 & ~x3 ;
  assign n16 = ~n14 & ~n15 ;
  assign n17 = ~n12 & n16 ;
  assign n18 = x6 & ~n17 ;
  assign n19 = ~x1 & ~x7 ;
  assign n20 = x3 & n19 ;
  assign n21 = x5 ^ x2 ;
  assign n22 = x5 ^ x1 ;
  assign n23 = x8 & x9 ;
  assign n24 = n23 ^ x1 ;
  assign n25 = ~x1 & ~n24 ;
  assign n26 = n25 ^ x1 ;
  assign n27 = n22 & ~n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n28 ^ x1 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = ~n21 & ~n30 ;
  assign n32 = ~n20 & n31 ;
  assign n33 = ~n18 & n32 ;
  assign n34 = x4 ^ x1 ;
  assign n35 = n34 ^ x7 ;
  assign n36 = x6 ^ x0 ;
  assign n37 = n13 ^ x6 ;
  assign n38 = n37 ^ n13 ;
  assign n39 = ~x3 & ~n19 ;
  assign n40 = n39 ^ n13 ;
  assign n41 = ~n38 & ~n40 ;
  assign n42 = n41 ^ n13 ;
  assign n43 = ~n36 & n42 ;
  assign n44 = n43 ^ x0 ;
  assign n45 = n35 & ~n44 ;
  assign n46 = n33 & n45 ;
  assign y0 = n46 ;
endmodule
