module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n8 = x2 & ~x3 ;
  assign n9 = ~x4 & ~n8 ;
  assign n11 = x5 ^ x3 ;
  assign n12 = n11 ^ x5 ;
  assign n21 = n12 ^ x5 ;
  assign n10 = x5 ^ x0 ;
  assign n13 = n12 ^ n10 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n14 ^ x5 ;
  assign n16 = ~x1 & x2 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n15 & ~n19 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n22 ^ n15 ;
  assign n24 = x1 & ~x4 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = n20 ^ n15 ;
  assign n27 = ~n25 & n26 ;
  assign n28 = n27 ^ x5 ;
  assign n29 = n23 & ~n28 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = n30 ^ n11 ;
  assign n32 = n31 ^ x5 ;
  assign n33 = ~n9 & ~n32 ;
  assign n34 = x6 & ~n33 ;
  assign y0 = n34 ;
endmodule
