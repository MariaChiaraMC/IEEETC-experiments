module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 ;
  assign n12 = x2 & x3 ;
  assign n8 = ~x3 & x6 ;
  assign n9 = ~x5 & ~x6 ;
  assign n10 = ~x2 & n9 ;
  assign n11 = ~n8 & ~n10 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = ~x2 & ~x3 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = n16 ^ n12 ;
  assign n18 = ~n14 & ~n17 ;
  assign n19 = n18 ^ n12 ;
  assign n20 = x1 & n19 ;
  assign n21 = n20 ^ n12 ;
  assign n22 = ~x4 & n21 ;
  assign n23 = ~x1 & x5 ;
  assign n24 = n15 & n23 ;
  assign n25 = ~x3 & x5 ;
  assign n26 = x6 & n25 ;
  assign n27 = x5 & x6 ;
  assign n28 = x3 & ~n27 ;
  assign n29 = x2 & ~n28 ;
  assign n30 = ~n26 & n29 ;
  assign n31 = ~n24 & ~n30 ;
  assign n32 = n31 ^ x4 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = n33 ^ x0 ;
  assign n35 = n12 & ~n23 ;
  assign n36 = ~n8 & ~n28 ;
  assign n37 = x6 ^ x5 ;
  assign n38 = ~x1 & n37 ;
  assign n39 = ~n36 & ~n38 ;
  assign n40 = ~x2 & ~n39 ;
  assign n41 = n40 ^ n35 ;
  assign n42 = ~n35 & n41 ;
  assign n43 = n42 ^ n31 ;
  assign n44 = n43 ^ n35 ;
  assign n45 = ~n34 & ~n44 ;
  assign n46 = n45 ^ n42 ;
  assign n47 = n46 ^ n35 ;
  assign n48 = ~x0 & ~n47 ;
  assign n49 = n48 ^ x0 ;
  assign n50 = ~n22 & n49 ;
  assign n51 = x3 & ~x4 ;
  assign n52 = n51 ^ n25 ;
  assign n53 = ~x1 & n52 ;
  assign n54 = n53 ^ n25 ;
  assign n55 = ~x3 & x4 ;
  assign n56 = ~x2 & ~n55 ;
  assign n57 = n56 ^ n51 ;
  assign n58 = n57 ^ x5 ;
  assign n59 = x6 ^ x1 ;
  assign n60 = n51 & ~n59 ;
  assign n61 = n60 ^ x1 ;
  assign n62 = ~n58 & ~n61 ;
  assign n63 = n62 ^ n60 ;
  assign n64 = n63 ^ x1 ;
  assign n65 = n64 ^ n51 ;
  assign n66 = ~x5 & ~n65 ;
  assign n67 = ~n54 & ~n66 ;
  assign n69 = n67 ^ x0 ;
  assign n68 = n67 ^ n55 ;
  assign n70 = n69 ^ n68 ;
  assign n71 = n70 ^ n69 ;
  assign n72 = n71 ^ n67 ;
  assign n73 = x2 & ~n9 ;
  assign n74 = n70 ^ x1 ;
  assign n75 = ~n73 & ~n74 ;
  assign n76 = n69 ^ n67 ;
  assign n77 = n71 & n76 ;
  assign n78 = n77 ^ n72 ;
  assign n79 = n75 & n78 ;
  assign n80 = n79 ^ n77 ;
  assign n81 = n72 & n80 ;
  assign n82 = n81 ^ n77 ;
  assign n83 = n82 ^ x0 ;
  assign n84 = n50 & ~n83 ;
  assign y0 = ~n84 ;
endmodule
