module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 ;
  assign n9 = ~x5 & x7 ;
  assign n10 = ~x4 & n9 ;
  assign n11 = x3 & ~x6 ;
  assign n12 = ~x0 & n11 ;
  assign n13 = n10 & n12 ;
  assign n14 = x4 & x6 ;
  assign n15 = x5 & ~x7 ;
  assign n16 = ~x0 & ~x3 ;
  assign n17 = n15 & n16 ;
  assign n18 = n14 & n17 ;
  assign n19 = ~x1 & n18 ;
  assign n20 = ~n13 & ~n19 ;
  assign n21 = x7 ^ x5 ;
  assign n22 = x6 ^ x3 ;
  assign n30 = n22 ^ x3 ;
  assign n31 = n30 ^ x3 ;
  assign n32 = ~n30 & n31 ;
  assign n23 = n22 ^ x7 ;
  assign n24 = n23 ^ x0 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n23 ^ n22 ;
  assign n27 = n26 ^ x3 ;
  assign n28 = n25 & n27 ;
  assign n35 = n32 ^ n28 ;
  assign n29 = n28 ^ n21 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = ~n29 & ~n33 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = ~n21 & n36 ;
  assign n38 = n37 ^ n28 ;
  assign n39 = n38 ^ n32 ;
  assign n40 = n39 ^ n34 ;
  assign n41 = ~x1 & n40 ;
  assign n42 = x1 & x6 ;
  assign n43 = n9 & n16 ;
  assign n44 = n42 & n43 ;
  assign n45 = ~x4 & ~n44 ;
  assign n46 = ~n41 & n45 ;
  assign n47 = x1 & ~x6 ;
  assign n48 = n43 & n47 ;
  assign n49 = ~x3 & x6 ;
  assign n50 = x1 & ~n49 ;
  assign n51 = n50 ^ x0 ;
  assign n52 = n11 ^ x7 ;
  assign n53 = n52 ^ n11 ;
  assign n54 = n53 ^ n21 ;
  assign n55 = x3 ^ x1 ;
  assign n56 = ~x1 & ~n55 ;
  assign n57 = n56 ^ n11 ;
  assign n58 = n57 ^ x1 ;
  assign n59 = n54 & n58 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = n60 ^ x1 ;
  assign n62 = ~n21 & ~n61 ;
  assign n63 = n62 ^ n50 ;
  assign n64 = n63 ^ n62 ;
  assign n65 = n64 ^ n51 ;
  assign n66 = x5 & ~x6 ;
  assign n67 = x3 & ~x5 ;
  assign n68 = ~n66 & ~n67 ;
  assign n69 = n68 ^ x7 ;
  assign n70 = n68 & ~n69 ;
  assign n71 = n70 ^ n62 ;
  assign n72 = n71 ^ n68 ;
  assign n73 = ~n65 & n72 ;
  assign n74 = n73 ^ n70 ;
  assign n75 = n74 ^ n68 ;
  assign n76 = ~n51 & n75 ;
  assign n77 = x4 & ~n76 ;
  assign n78 = ~n48 & n77 ;
  assign n79 = ~n46 & ~n78 ;
  assign n80 = n79 ^ x2 ;
  assign n81 = n80 ^ n79 ;
  assign n82 = n81 ^ n20 ;
  assign n83 = x5 & x7 ;
  assign n84 = ~n14 & ~n47 ;
  assign n85 = n83 & n84 ;
  assign n86 = n85 ^ x0 ;
  assign n87 = n86 ^ n85 ;
  assign n88 = n15 ^ x6 ;
  assign n89 = n88 ^ n15 ;
  assign n90 = n15 ^ n10 ;
  assign n91 = n89 & n90 ;
  assign n92 = n91 ^ n15 ;
  assign n93 = x1 & n92 ;
  assign n94 = n93 ^ n85 ;
  assign n95 = n87 & n94 ;
  assign n96 = n95 ^ n85 ;
  assign n97 = x3 & ~n96 ;
  assign n98 = ~x4 & ~x6 ;
  assign n99 = x0 & ~n98 ;
  assign n100 = x6 ^ x4 ;
  assign n101 = ~x5 & n100 ;
  assign n102 = ~x0 & ~n101 ;
  assign n103 = ~x1 & ~n102 ;
  assign n104 = n103 ^ x7 ;
  assign n105 = n104 ^ n103 ;
  assign n106 = n42 ^ x6 ;
  assign n107 = ~x5 & ~n106 ;
  assign n108 = n107 ^ x6 ;
  assign n109 = x4 & ~n108 ;
  assign n110 = n109 ^ n103 ;
  assign n111 = ~n105 & n110 ;
  assign n112 = n111 ^ n103 ;
  assign n113 = ~n99 & n112 ;
  assign n114 = ~x3 & ~n113 ;
  assign n115 = n114 ^ n97 ;
  assign n116 = ~n97 & n115 ;
  assign n117 = n116 ^ n79 ;
  assign n118 = n117 ^ n97 ;
  assign n119 = n82 & ~n118 ;
  assign n120 = n119 ^ n116 ;
  assign n121 = n120 ^ n97 ;
  assign n122 = n20 & ~n121 ;
  assign n123 = n122 ^ n20 ;
  assign y0 = ~n123 ;
endmodule
