module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 ;
  assign n17 = x7 & ~x14 ;
  assign n18 = ~x5 & x6 ;
  assign n19 = n17 & n18 ;
  assign n20 = x3 & x4 ;
  assign n21 = ~x2 & x15 ;
  assign n22 = n20 & n21 ;
  assign n23 = x0 & x1 ;
  assign n24 = n22 & n23 ;
  assign n25 = n19 & n24 ;
  assign n26 = x6 & ~x9 ;
  assign n27 = x8 & ~x15 ;
  assign n28 = x5 & n27 ;
  assign n29 = n26 & n28 ;
  assign n30 = x4 & ~n29 ;
  assign n31 = ~x0 & ~x1 ;
  assign n32 = x10 & n31 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = x9 & x14 ;
  assign n35 = n18 & n34 ;
  assign n36 = ~x3 & x11 ;
  assign n37 = n27 & n36 ;
  assign n38 = n35 & n37 ;
  assign n39 = ~x7 & n38 ;
  assign n40 = n39 ^ x2 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = ~x6 & ~x8 ;
  assign n43 = x15 & n42 ;
  assign n44 = x3 & ~x5 ;
  assign n45 = n43 & n44 ;
  assign n46 = ~n20 & ~n45 ;
  assign n47 = n17 & ~n46 ;
  assign n48 = n47 ^ n39 ;
  assign n49 = n41 & n48 ;
  assign n50 = n49 ^ n39 ;
  assign n51 = n50 ^ n30 ;
  assign n52 = ~n33 & ~n51 ;
  assign n53 = n52 ^ n49 ;
  assign n54 = n53 ^ n39 ;
  assign n55 = n54 ^ n32 ;
  assign n56 = ~n30 & n55 ;
  assign n57 = n56 ^ n30 ;
  assign n58 = ~n25 & n57 ;
  assign n59 = ~x12 & ~x13 ;
  assign n60 = ~n58 & n59 ;
  assign y0 = n60 ;
endmodule
