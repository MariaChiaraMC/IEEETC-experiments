module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 ;
  assign n19 = x5 ^ x3 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = n20 ^ x7 ;
  assign n22 = n21 ^ x7 ;
  assign n24 = x4 ^ x3 ;
  assign n23 = x6 ^ x3 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ x7 ;
  assign n27 = n26 ^ n22 ;
  assign n31 = n22 ^ n21 ;
  assign n32 = ~x3 & n31 ;
  assign n28 = n24 ^ x3 ;
  assign n29 = n28 ^ x3 ;
  assign n30 = ~n21 & ~n29 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ x3 ;
  assign n35 = n34 ^ n28 ;
  assign n36 = n27 & ~n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = ~n22 & n37 ;
  assign n39 = n38 ^ n30 ;
  assign n40 = n39 ^ n36 ;
  assign n41 = n40 ^ x3 ;
  assign n17 = x3 ^ x0 ;
  assign n18 = n17 ^ x3 ;
  assign n42 = n41 ^ n18 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = n43 ^ n17 ;
  assign n45 = n44 ^ n43 ;
  assign n46 = x7 & n45 ;
  assign n47 = n46 ^ n41 ;
  assign n48 = ~x10 & ~x11 ;
  assign n49 = x9 & n48 ;
  assign n50 = ~x8 & n49 ;
  assign n51 = x14 & x15 ;
  assign n52 = x14 ^ x13 ;
  assign n53 = n52 ^ x15 ;
  assign n54 = n51 & n53 ;
  assign n55 = n54 ^ n53 ;
  assign n56 = n50 & n55 ;
  assign n57 = ~x12 & n56 ;
  assign n58 = n57 ^ n41 ;
  assign n59 = ~n44 & n58 ;
  assign n60 = n59 ^ n43 ;
  assign n61 = n60 ^ n44 ;
  assign n62 = ~n47 & n61 ;
  assign n63 = ~n43 & n62 ;
  assign n64 = n63 ^ n46 ;
  assign y0 = n64 ;
endmodule
