module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 ;
  assign n9 = x1 ^ x0 ;
  assign n10 = x2 & x3 ;
  assign n11 = n10 ^ x1 ;
  assign n12 = n11 ^ x1 ;
  assign n13 = n12 ^ n9 ;
  assign n14 = ~x5 & ~x7 ;
  assign n15 = ~x6 & n14 ;
  assign n16 = n15 ^ x1 ;
  assign n17 = x4 ^ x1 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = ~n16 & ~n18 ;
  assign n20 = n19 ^ x1 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = ~n13 & ~n21 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n23 ^ n16 ;
  assign n25 = ~n9 & ~n24 ;
  assign n26 = n25 ^ n9 ;
  assign y0 = n26 ;
endmodule
