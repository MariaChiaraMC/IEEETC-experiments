module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 ;
  output y0 ;
  wire n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 ;
  assign n26 = ~x4 & ~x5 ;
  assign n27 = x24 & n26 ;
  assign n28 = x10 & n27 ;
  assign n29 = ~x1 & ~x2 ;
  assign n30 = ~x0 & ~x3 ;
  assign n31 = n29 & n30 ;
  assign n32 = x11 & n31 ;
  assign n33 = n28 & n32 ;
  assign n34 = x20 & x21 ;
  assign n35 = x19 & n34 ;
  assign n36 = n35 ^ x22 ;
  assign n37 = n36 ^ x22 ;
  assign n38 = x22 ^ x18 ;
  assign n39 = n38 ^ x22 ;
  assign n40 = n37 & n39 ;
  assign n41 = n40 ^ x22 ;
  assign n42 = ~x13 & n41 ;
  assign n43 = n42 ^ x22 ;
  assign n44 = n33 & n43 ;
  assign n45 = x10 & ~x11 ;
  assign n46 = n29 & n45 ;
  assign n47 = ~x24 & n30 ;
  assign n48 = n46 & ~n47 ;
  assign n49 = ~x13 & ~x14 ;
  assign n50 = ~x16 & ~n49 ;
  assign n51 = x15 & ~x17 ;
  assign n52 = ~n50 & n51 ;
  assign n53 = n48 & n52 ;
  assign n54 = n26 & n53 ;
  assign n55 = x16 ^ x3 ;
  assign n56 = x14 ^ x13 ;
  assign n57 = n56 ^ x16 ;
  assign n58 = x3 ^ x0 ;
  assign n59 = n58 ^ n56 ;
  assign n60 = ~n56 & n59 ;
  assign n61 = n60 ^ n56 ;
  assign n62 = ~n57 & ~n61 ;
  assign n63 = n62 ^ n60 ;
  assign n64 = n63 ^ n56 ;
  assign n65 = n64 ^ n58 ;
  assign n66 = n55 & n65 ;
  assign n67 = n66 ^ x16 ;
  assign n68 = n54 & ~n67 ;
  assign n69 = ~x12 & ~n68 ;
  assign n70 = ~n44 & n69 ;
  assign n71 = ~x10 & x11 ;
  assign n72 = n29 ^ x0 ;
  assign n79 = x4 & x5 ;
  assign n80 = ~x3 & ~n79 ;
  assign n81 = ~n26 & ~n80 ;
  assign n82 = ~n30 & ~n81 ;
  assign n73 = x0 & ~x16 ;
  assign n74 = ~x3 & n26 ;
  assign n75 = x13 & ~x14 ;
  assign n76 = ~x15 & n75 ;
  assign n77 = n74 & n76 ;
  assign n78 = n73 & n77 ;
  assign n83 = n82 ^ n78 ;
  assign n84 = n83 ^ x17 ;
  assign n95 = n84 ^ n83 ;
  assign n85 = ~x13 & x14 ;
  assign n86 = x15 & x17 ;
  assign n87 = x16 & n86 ;
  assign n88 = n85 & n87 ;
  assign n89 = n88 ^ n84 ;
  assign n90 = n89 ^ n83 ;
  assign n91 = n84 ^ n78 ;
  assign n92 = n91 ^ n88 ;
  assign n93 = n92 ^ n90 ;
  assign n94 = ~n90 & ~n93 ;
  assign n96 = n95 ^ n94 ;
  assign n97 = n96 ^ n90 ;
  assign n98 = ~x15 & ~x16 ;
  assign n99 = x13 & n98 ;
  assign n100 = x14 & n99 ;
  assign n101 = n100 ^ n83 ;
  assign n102 = n94 ^ n90 ;
  assign n103 = ~n101 & ~n102 ;
  assign n104 = n103 ^ n83 ;
  assign n105 = ~n97 & n104 ;
  assign n106 = n105 ^ n83 ;
  assign n107 = n106 ^ n82 ;
  assign n108 = n107 ^ n83 ;
  assign n109 = n108 ^ n72 ;
  assign n110 = n109 ^ n29 ;
  assign n111 = n110 ^ n109 ;
  assign n112 = ~x1 & ~n27 ;
  assign n113 = x17 ^ x14 ;
  assign n114 = n99 & n113 ;
  assign n115 = ~n88 & ~n114 ;
  assign n116 = ~n112 & ~n115 ;
  assign n117 = x14 & x17 ;
  assign n118 = x5 & ~n117 ;
  assign n119 = ~x4 & ~n118 ;
  assign n121 = ~x1 & ~x5 ;
  assign n122 = ~x3 & ~n121 ;
  assign n123 = ~x2 & n122 ;
  assign n120 = ~x1 & ~n113 ;
  assign n124 = n123 ^ n120 ;
  assign n125 = ~n119 & n124 ;
  assign n126 = n125 ^ n123 ;
  assign n127 = n99 & n126 ;
  assign n128 = ~x1 & n99 ;
  assign n129 = ~n88 & ~n128 ;
  assign n130 = ~x2 & n80 ;
  assign n131 = ~n129 & ~n130 ;
  assign n132 = ~n127 & ~n131 ;
  assign n133 = ~n116 & n132 ;
  assign n134 = n133 ^ n109 ;
  assign n135 = n134 ^ n72 ;
  assign n136 = n111 & n135 ;
  assign n137 = n136 ^ n133 ;
  assign n138 = n85 & n98 ;
  assign n139 = n75 & n87 ;
  assign n140 = ~n138 & ~n139 ;
  assign n141 = ~x3 & n27 ;
  assign n142 = ~n140 & n141 ;
  assign n143 = n133 & ~n142 ;
  assign n144 = n143 ^ n72 ;
  assign n145 = n137 & n144 ;
  assign n146 = n145 ^ n143 ;
  assign n147 = n72 & n146 ;
  assign n148 = n147 ^ n136 ;
  assign n149 = n148 ^ x0 ;
  assign n150 = n149 ^ n133 ;
  assign n151 = n71 & ~n150 ;
  assign n152 = n70 & ~n151 ;
  assign n153 = n33 & n76 ;
  assign n154 = x12 & ~n153 ;
  assign n155 = ~x8 & ~x9 ;
  assign n156 = ~x6 & ~x23 ;
  assign n157 = n155 & n156 ;
  assign n158 = ~x7 & n157 ;
  assign n159 = ~n154 & n158 ;
  assign n160 = ~n152 & n159 ;
  assign y0 = n160 ;
endmodule
