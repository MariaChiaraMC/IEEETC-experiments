module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 ;
  assign n9 = x3 ^ x2 ;
  assign n10 = n9 ^ x1 ;
  assign n18 = x4 & ~x5 ;
  assign n11 = x6 ^ x5 ;
  assign n12 = x7 ^ x4 ;
  assign n13 = x6 ^ x4 ;
  assign n14 = ~n12 & ~n13 ;
  assign n15 = n14 ^ x4 ;
  assign n16 = ~n11 & n15 ;
  assign n17 = n16 ^ x4 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = ~x2 & n19 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n10 & ~n21 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n23 ^ n18 ;
  assign n25 = n24 ^ x2 ;
  assign n26 = ~x1 & n25 ;
  assign y0 = ~n26 ;
endmodule
