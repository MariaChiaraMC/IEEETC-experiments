module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 ;
  assign n59 = ~x0 & ~x3 ;
  assign n60 = x5 & ~x6 ;
  assign n61 = n60 ^ x7 ;
  assign n62 = x8 ^ x1 ;
  assign n63 = n62 ^ x8 ;
  assign n64 = ~x8 & x9 ;
  assign n65 = n64 ^ x8 ;
  assign n66 = ~n63 & n65 ;
  assign n67 = n66 ^ x8 ;
  assign n68 = n67 ^ n60 ;
  assign n69 = n61 & n68 ;
  assign n70 = n69 ^ n66 ;
  assign n71 = n70 ^ x8 ;
  assign n72 = n71 ^ x7 ;
  assign n73 = n60 & n72 ;
  assign n74 = n73 ^ n60 ;
  assign n75 = n59 & n74 ;
  assign n76 = ~x6 & ~x8 ;
  assign n77 = ~x1 & ~n76 ;
  assign n78 = ~x7 & x9 ;
  assign n79 = n59 & n78 ;
  assign n80 = n77 & n79 ;
  assign n81 = x1 & ~x7 ;
  assign n82 = x0 & ~x6 ;
  assign n83 = n81 & n82 ;
  assign n84 = n64 & n83 ;
  assign n85 = ~n80 & ~n84 ;
  assign n86 = n85 ^ x5 ;
  assign n87 = n86 ^ n85 ;
  assign n88 = n87 ^ n75 ;
  assign n89 = ~x1 & x3 ;
  assign n90 = ~x6 & ~x9 ;
  assign n91 = x7 & x8 ;
  assign n92 = n90 & n91 ;
  assign n93 = x6 & x8 ;
  assign n94 = n78 & n93 ;
  assign n95 = ~n92 & ~n94 ;
  assign n96 = n89 & ~n95 ;
  assign n97 = ~x3 & ~x7 ;
  assign n98 = x6 ^ x1 ;
  assign n99 = n98 ^ x9 ;
  assign n100 = n99 ^ n98 ;
  assign n101 = n100 ^ n97 ;
  assign n50 = x1 & ~x8 ;
  assign n102 = n98 ^ n50 ;
  assign n103 = n101 & n102 ;
  assign n104 = n103 ^ n50 ;
  assign n105 = n97 & n104 ;
  assign n106 = ~n96 & ~n105 ;
  assign n107 = ~x0 & n106 ;
  assign n108 = ~x8 & n89 ;
  assign n109 = n90 & n108 ;
  assign n25 = x3 & x8 ;
  assign n11 = ~x3 & ~x8 ;
  assign n110 = n25 ^ n11 ;
  assign n111 = x6 & n110 ;
  assign n112 = n111 ^ n25 ;
  assign n113 = x9 & n112 ;
  assign n114 = x1 & n113 ;
  assign n115 = ~n109 & ~n114 ;
  assign n116 = n115 ^ x7 ;
  assign n117 = n116 ^ n115 ;
  assign n118 = n117 ^ x0 ;
  assign n119 = ~x3 & x8 ;
  assign n120 = x9 & n119 ;
  assign n121 = n120 ^ x1 ;
  assign n122 = x1 & n121 ;
  assign n123 = n122 ^ n115 ;
  assign n124 = n123 ^ x1 ;
  assign n125 = ~n118 & ~n124 ;
  assign n126 = n125 ^ n122 ;
  assign n127 = n126 ^ x1 ;
  assign n128 = x0 & n127 ;
  assign n129 = n128 ^ x0 ;
  assign n130 = n129 ^ n107 ;
  assign n131 = ~n107 & n130 ;
  assign n132 = n131 ^ n85 ;
  assign n133 = n132 ^ n107 ;
  assign n134 = n88 & n133 ;
  assign n135 = n134 ^ n131 ;
  assign n136 = n135 ^ n107 ;
  assign n137 = ~n75 & ~n136 ;
  assign n138 = n137 ^ n75 ;
  assign n24 = ~x5 & x9 ;
  assign n26 = ~x6 & n25 ;
  assign n27 = n24 & n26 ;
  assign n15 = ~x3 & ~x6 ;
  assign n28 = ~n15 & ~n25 ;
  assign n29 = ~x5 & ~x9 ;
  assign n30 = x6 & ~x8 ;
  assign n31 = n29 & ~n30 ;
  assign n32 = n28 & n31 ;
  assign n33 = ~n27 & ~n32 ;
  assign n12 = n11 ^ x5 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n13 ^ x9 ;
  assign n16 = n15 ^ x8 ;
  assign n17 = x8 & n16 ;
  assign n18 = n17 ^ n11 ;
  assign n19 = n18 ^ x8 ;
  assign n20 = ~n14 & n19 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n21 ^ x8 ;
  assign n23 = ~x9 & n22 ;
  assign n34 = n33 ^ n23 ;
  assign n35 = x1 & ~n34 ;
  assign n36 = n35 ^ n23 ;
  assign n37 = n36 ^ x0 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = x6 & ~x9 ;
  assign n40 = x5 & n11 ;
  assign n41 = n39 & n40 ;
  assign n42 = ~n27 & ~n41 ;
  assign n43 = ~x1 & ~n42 ;
  assign n44 = x6 & x9 ;
  assign n45 = ~x3 & ~x5 ;
  assign n46 = n44 & n45 ;
  assign n47 = x8 & n46 ;
  assign n48 = x3 & x5 ;
  assign n49 = ~x6 & x9 ;
  assign n51 = n49 & n50 ;
  assign n52 = n48 & n51 ;
  assign n53 = ~n47 & ~n52 ;
  assign n54 = ~n43 & n53 ;
  assign n55 = n54 ^ n36 ;
  assign n56 = n38 & ~n55 ;
  assign n57 = n56 ^ n36 ;
  assign n58 = x7 & ~n57 ;
  assign n139 = n138 ^ n58 ;
  assign n140 = n139 ^ n138 ;
  assign n141 = ~n11 & ~n25 ;
  assign n142 = x0 & x5 ;
  assign n143 = n39 & n142 ;
  assign n144 = n141 & n143 ;
  assign n145 = ~x5 & x6 ;
  assign n146 = ~n119 & n145 ;
  assign n147 = ~x0 & x3 ;
  assign n148 = ~x9 & n147 ;
  assign n149 = x8 & ~x9 ;
  assign n150 = x0 & ~n149 ;
  assign n151 = ~n148 & ~n150 ;
  assign n152 = n146 & n151 ;
  assign n153 = n25 ^ x5 ;
  assign n154 = n153 ^ n25 ;
  assign n155 = n110 & ~n154 ;
  assign n156 = n155 ^ n25 ;
  assign n157 = x9 & n156 ;
  assign n158 = n82 & n157 ;
  assign n159 = ~n152 & ~n158 ;
  assign n160 = ~n144 & n159 ;
  assign n161 = x1 & ~n160 ;
  assign n162 = x5 & x9 ;
  assign n163 = ~n90 & ~n162 ;
  assign n164 = x0 & ~n60 ;
  assign n165 = n108 & n164 ;
  assign n166 = ~n163 & n165 ;
  assign n167 = ~x7 & ~n166 ;
  assign n168 = ~n161 & n167 ;
  assign n169 = n168 ^ n138 ;
  assign n170 = n169 ^ n138 ;
  assign n171 = ~n140 & ~n170 ;
  assign n172 = n171 ^ n138 ;
  assign n173 = x4 & n172 ;
  assign n174 = n173 ^ n138 ;
  assign n175 = ~x2 & ~n174 ;
  assign n176 = ~x4 & ~x5 ;
  assign n177 = n59 & n176 ;
  assign n178 = n92 & n177 ;
  assign n179 = n178 ^ x2 ;
  assign n180 = x4 & ~x8 ;
  assign n181 = ~x4 & n93 ;
  assign n182 = ~n180 & ~n181 ;
  assign n183 = x0 & x3 ;
  assign n184 = n29 & n183 ;
  assign n185 = ~n182 & n184 ;
  assign n193 = ~x5 & n90 ;
  assign n188 = ~n24 & n25 ;
  assign n189 = ~x5 & n39 ;
  assign n190 = ~n49 & ~n189 ;
  assign n191 = n188 & ~n190 ;
  assign n194 = n193 ^ n191 ;
  assign n186 = x8 ^ x6 ;
  assign n187 = n162 & ~n186 ;
  assign n192 = n191 ^ n187 ;
  assign n195 = n194 ^ n192 ;
  assign n196 = n194 ^ x3 ;
  assign n197 = n196 ^ n194 ;
  assign n198 = n195 & ~n197 ;
  assign n199 = n198 ^ n194 ;
  assign n200 = ~x4 & n199 ;
  assign n201 = n200 ^ n191 ;
  assign n202 = n201 ^ x0 ;
  assign n203 = n202 ^ n201 ;
  assign n204 = n203 ^ n185 ;
  assign n205 = x8 ^ x4 ;
  assign n206 = n44 ^ x8 ;
  assign n207 = n206 ^ x3 ;
  assign n208 = n207 ^ n44 ;
  assign n209 = n208 ^ n205 ;
  assign n210 = n90 ^ x3 ;
  assign n211 = n90 & ~n210 ;
  assign n212 = n211 ^ n44 ;
  assign n213 = n212 ^ n90 ;
  assign n214 = ~n209 & n213 ;
  assign n215 = n214 ^ n211 ;
  assign n216 = n215 ^ n90 ;
  assign n217 = ~n205 & n216 ;
  assign n218 = n217 ^ x5 ;
  assign n219 = n217 & n218 ;
  assign n220 = n219 ^ n201 ;
  assign n221 = n220 ^ n217 ;
  assign n222 = ~n204 & n221 ;
  assign n223 = n222 ^ n219 ;
  assign n224 = n223 ^ n217 ;
  assign n225 = ~n185 & n224 ;
  assign n226 = n225 ^ n185 ;
  assign n227 = x7 & n226 ;
  assign n234 = n78 & ~n147 ;
  assign n235 = ~n141 & n176 ;
  assign n236 = n234 & n235 ;
  assign n237 = ~x0 & ~x9 ;
  assign n238 = n48 & n237 ;
  assign n239 = n180 & n238 ;
  assign n240 = ~n236 & ~n239 ;
  assign n228 = x4 & ~x7 ;
  assign n241 = n228 ^ n119 ;
  assign n242 = n24 ^ x0 ;
  assign n243 = n242 ^ n24 ;
  assign n229 = ~n29 & ~n162 ;
  assign n244 = n229 ^ n24 ;
  assign n245 = n243 & ~n244 ;
  assign n246 = n245 ^ n24 ;
  assign n247 = n246 ^ n119 ;
  assign n248 = n241 & n247 ;
  assign n249 = n248 ^ n245 ;
  assign n250 = n249 ^ n24 ;
  assign n251 = n250 ^ n228 ;
  assign n252 = n119 & n251 ;
  assign n253 = n252 ^ n119 ;
  assign n254 = n240 & ~n253 ;
  assign n230 = ~x0 & x5 ;
  assign n231 = x8 & ~n230 ;
  assign n232 = ~n229 & ~n231 ;
  assign n233 = n228 & n232 ;
  assign n255 = n254 ^ n233 ;
  assign n256 = n255 ^ n254 ;
  assign n257 = n254 ^ x3 ;
  assign n258 = n257 ^ n254 ;
  assign n259 = n256 & ~n258 ;
  assign n260 = n259 ^ n254 ;
  assign n261 = ~x6 & ~n260 ;
  assign n262 = n261 ^ n254 ;
  assign n263 = ~n227 & n262 ;
  assign n264 = n263 ^ x1 ;
  assign n265 = n264 ^ n263 ;
  assign n272 = ~x5 & n119 ;
  assign n302 = ~x7 & ~n272 ;
  assign n303 = x5 ^ x0 ;
  assign n304 = n49 & ~n303 ;
  assign n305 = ~n91 & n304 ;
  assign n306 = ~n302 & n305 ;
  assign n266 = n44 & n183 ;
  assign n267 = ~x5 & n266 ;
  assign n268 = x6 ^ x5 ;
  assign n269 = n148 & n268 ;
  assign n270 = ~n267 & ~n269 ;
  assign n271 = ~x8 & ~n270 ;
  assign n273 = ~n40 & ~n272 ;
  assign n274 = n90 & ~n273 ;
  assign n275 = x0 & n274 ;
  assign n276 = ~n271 & ~n275 ;
  assign n277 = n276 ^ x8 ;
  assign n278 = n277 ^ n276 ;
  assign n279 = x3 ^ x0 ;
  assign n280 = n279 ^ x5 ;
  assign n281 = n44 ^ x5 ;
  assign n282 = n281 ^ n44 ;
  assign n283 = n282 ^ n280 ;
  assign n284 = n90 & n210 ;
  assign n285 = n284 ^ n44 ;
  assign n286 = n285 ^ n90 ;
  assign n287 = ~n283 & n286 ;
  assign n288 = n287 ^ n284 ;
  assign n289 = n288 ^ n90 ;
  assign n290 = ~n280 & n289 ;
  assign n291 = n290 ^ n276 ;
  assign n292 = n291 ^ n276 ;
  assign n293 = n278 & n292 ;
  assign n294 = n293 ^ n276 ;
  assign n295 = x7 & ~n294 ;
  assign n296 = n295 ^ n276 ;
  assign n307 = n306 ^ n296 ;
  assign n308 = n307 ^ n296 ;
  assign n297 = n60 & n237 ;
  assign n298 = ~n91 & n297 ;
  assign n299 = ~n141 & n298 ;
  assign n300 = n299 ^ n296 ;
  assign n301 = n300 ^ n296 ;
  assign n309 = n308 ^ n301 ;
  assign n310 = n28 ^ x3 ;
  assign n311 = n310 ^ n28 ;
  assign n312 = n93 ^ n28 ;
  assign n313 = n312 ^ n28 ;
  assign n314 = ~n311 & n313 ;
  assign n315 = n314 ^ n28 ;
  assign n316 = ~x0 & ~n315 ;
  assign n317 = n316 ^ n28 ;
  assign n318 = n29 & ~n317 ;
  assign n319 = x7 & n318 ;
  assign n320 = n319 ^ n296 ;
  assign n321 = n320 ^ n296 ;
  assign n322 = n321 ^ n308 ;
  assign n323 = ~n308 & n322 ;
  assign n324 = n323 ^ n308 ;
  assign n325 = n309 & ~n324 ;
  assign n326 = n325 ^ n323 ;
  assign n327 = n326 ^ n296 ;
  assign n328 = n327 ^ n308 ;
  assign n329 = x4 & ~n328 ;
  assign n330 = n329 ^ n296 ;
  assign n331 = n330 ^ n263 ;
  assign n332 = ~n265 & n331 ;
  assign n333 = n332 ^ n263 ;
  assign n334 = n333 ^ n178 ;
  assign n335 = ~n179 & ~n334 ;
  assign n336 = n335 ^ n332 ;
  assign n337 = n336 ^ n263 ;
  assign n338 = n337 ^ x2 ;
  assign n339 = ~n178 & n338 ;
  assign n340 = n339 ^ n178 ;
  assign n341 = ~n175 & n340 ;
  assign y0 = n341 ;
endmodule
