module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 ;
  assign n9 = ~x5 & ~x7 ;
  assign n10 = ~x2 & x3 ;
  assign n11 = n9 & n10 ;
  assign n12 = ~x6 & n11 ;
  assign n13 = x4 & n12 ;
  assign n19 = x3 & ~x5 ;
  assign n20 = x7 & n19 ;
  assign n33 = ~x2 & n20 ;
  assign n36 = n33 ^ n9 ;
  assign n34 = x5 & x7 ;
  assign n35 = n34 ^ n33 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = n36 ^ x3 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n37 & n39 ;
  assign n41 = n40 ^ n36 ;
  assign n42 = x0 & n41 ;
  assign n43 = n42 ^ n33 ;
  assign n44 = ~x4 & n43 ;
  assign n45 = ~x0 & x4 ;
  assign n46 = ~n19 & n45 ;
  assign n16 = ~x3 & x5 ;
  assign n47 = n16 ^ x7 ;
  assign n48 = n47 ^ x7 ;
  assign n49 = x7 ^ x2 ;
  assign n50 = ~n48 & n49 ;
  assign n51 = n50 ^ x7 ;
  assign n52 = n46 & ~n51 ;
  assign n53 = ~n44 & ~n52 ;
  assign n14 = x6 ^ x4 ;
  assign n15 = n14 ^ x0 ;
  assign n17 = n16 ^ x6 ;
  assign n18 = n17 ^ n16 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = ~n18 & n21 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = n23 ^ n14 ;
  assign n25 = ~n15 & ~n24 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = n26 ^ n16 ;
  assign n28 = n27 ^ x0 ;
  assign n29 = ~n14 & n28 ;
  assign n30 = n29 ^ n14 ;
  assign n31 = n30 ^ x0 ;
  assign n32 = x2 & n31 ;
  assign n54 = n53 ^ n32 ;
  assign n55 = n54 ^ x6 ;
  assign n66 = n55 ^ n54 ;
  assign n56 = x5 & x6 ;
  assign n57 = ~x7 & n56 ;
  assign n58 = ~x3 & n57 ;
  assign n59 = ~x0 & ~n58 ;
  assign n60 = n59 ^ n55 ;
  assign n61 = n60 ^ n54 ;
  assign n62 = n59 ^ n32 ;
  assign n63 = n62 ^ n59 ;
  assign n64 = n63 ^ n61 ;
  assign n65 = n61 & n64 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = n67 ^ n61 ;
  assign n69 = n34 ^ x7 ;
  assign n70 = x4 ^ x3 ;
  assign n71 = n70 ^ x3 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = n34 ^ n19 ;
  assign n74 = ~n19 & n73 ;
  assign n75 = n74 ^ x3 ;
  assign n76 = n75 ^ n19 ;
  assign n77 = n72 & ~n76 ;
  assign n78 = n77 ^ n74 ;
  assign n79 = n78 ^ n19 ;
  assign n80 = ~n69 & ~n79 ;
  assign n81 = n80 ^ x7 ;
  assign n82 = n81 ^ n54 ;
  assign n83 = n65 ^ n61 ;
  assign n84 = ~n82 & n83 ;
  assign n85 = n84 ^ n54 ;
  assign n86 = n68 & ~n85 ;
  assign n87 = n86 ^ n54 ;
  assign n88 = n87 ^ n32 ;
  assign n89 = n88 ^ n54 ;
  assign n90 = ~n13 & ~n89 ;
  assign n91 = ~x1 & ~n90 ;
  assign n92 = n45 & n57 ;
  assign n93 = x0 & x7 ;
  assign n94 = n93 ^ x6 ;
  assign n95 = n93 ^ x5 ;
  assign n96 = n94 & ~n95 ;
  assign n97 = n96 ^ n93 ;
  assign n98 = ~x4 & ~n93 ;
  assign n99 = n98 ^ x1 ;
  assign n100 = ~n97 & n99 ;
  assign n101 = n100 ^ n98 ;
  assign n102 = x1 & n101 ;
  assign n103 = n102 ^ x1 ;
  assign n104 = ~n92 & ~n103 ;
  assign n105 = n10 & ~n104 ;
  assign n106 = ~x3 & n45 ;
  assign n107 = x2 & x6 ;
  assign n108 = x1 & x5 ;
  assign n109 = n108 ^ n9 ;
  assign n110 = n107 & n109 ;
  assign n111 = n110 ^ n9 ;
  assign n112 = n106 & n111 ;
  assign n113 = n107 & n108 ;
  assign n114 = ~x3 & n107 ;
  assign n115 = ~x5 & n114 ;
  assign n116 = x0 & ~n115 ;
  assign n117 = ~n113 & n116 ;
  assign n118 = ~n93 & ~n117 ;
  assign n119 = ~x2 & ~x3 ;
  assign n120 = ~x5 & x6 ;
  assign n121 = ~n34 & ~n120 ;
  assign n122 = n119 & n121 ;
  assign n123 = x1 & n122 ;
  assign n124 = ~n118 & ~n123 ;
  assign n125 = x7 & n16 ;
  assign n126 = ~n11 & ~n125 ;
  assign n127 = x1 & ~x6 ;
  assign n128 = ~n126 & n127 ;
  assign n129 = n56 & n119 ;
  assign n130 = x7 & n129 ;
  assign n131 = ~x0 & ~n130 ;
  assign n132 = ~n128 & n131 ;
  assign n133 = ~x4 & ~n132 ;
  assign n134 = ~n124 & n133 ;
  assign n135 = ~n112 & ~n134 ;
  assign n136 = ~n105 & n135 ;
  assign n137 = ~n91 & n136 ;
  assign y0 = ~n137 ;
endmodule
