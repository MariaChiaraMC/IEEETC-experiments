// Benchmark "./p3.pla" written by ABC on Thu Apr 23 10:59:59 2020

module \./p3.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z0  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z0;
  assign z0 = 1'b1;
endmodule


