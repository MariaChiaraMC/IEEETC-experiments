module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n9 = x5 ^ x4 ;
  assign n10 = n9 ^ x6 ;
  assign n11 = x5 ^ x2 ;
  assign n12 = n11 ^ x6 ;
  assign n13 = n12 ^ n10 ;
  assign n14 = x7 ^ x6 ;
  assign n15 = n14 ^ x2 ;
  assign n16 = ~x2 & n15 ;
  assign n17 = n16 ^ x6 ;
  assign n18 = n17 ^ x2 ;
  assign n19 = n13 & n18 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = n10 & ~n21 ;
  assign n23 = n22 ^ x2 ;
  assign n24 = ~x3 & n23 ;
  assign n25 = x4 & ~x5 ;
  assign n26 = x2 & n25 ;
  assign n27 = ~x1 & ~n26 ;
  assign n28 = ~n24 & n27 ;
  assign n29 = ~x0 & ~n28 ;
  assign y0 = n29 ;
endmodule
