module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 ;
  assign n13 = ~x5 & x11 ;
  assign n14 = ~x9 & x10 ;
  assign n29 = x4 & x8 ;
  assign n30 = ~x6 & n29 ;
  assign n15 = x7 ^ x4 ;
  assign n16 = x8 ^ x7 ;
  assign n17 = n16 ^ x8 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = n16 ^ x2 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = ~n18 & n20 ;
  assign n22 = n21 ^ n16 ;
  assign n23 = ~x1 & ~n16 ;
  assign n24 = n23 ^ n15 ;
  assign n25 = ~n22 & ~n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = ~n15 & n26 ;
  assign n28 = n27 ^ n15 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = n30 ^ x6 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = ~n32 & n34 ;
  assign n36 = n35 ^ n30 ;
  assign n37 = n14 & n36 ;
  assign n38 = n37 ^ n30 ;
  assign n39 = n13 & n38 ;
  assign n40 = ~x11 & n30 ;
  assign n41 = x7 ^ x5 ;
  assign n42 = n40 & ~n41 ;
  assign n43 = ~n39 & ~n42 ;
  assign n44 = ~x0 & ~n43 ;
  assign y0 = n44 ;
endmodule
