module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 ;
  assign n9 = ~x5 & x7 ;
  assign n10 = x0 & x3 ;
  assign n11 = x4 & n10 ;
  assign n12 = n9 & n11 ;
  assign n13 = x2 ^ x1 ;
  assign n14 = n12 & n13 ;
  assign n15 = ~x1 & x2 ;
  assign n16 = n9 & n15 ;
  assign n17 = x5 ^ x2 ;
  assign n18 = n17 ^ x1 ;
  assign n19 = x7 ^ x0 ;
  assign n20 = x5 ^ x0 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = n21 ^ x0 ;
  assign n23 = n22 ^ n17 ;
  assign n24 = ~n18 & ~n23 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ x0 ;
  assign n27 = n26 ^ x1 ;
  assign n28 = ~n17 & n27 ;
  assign n29 = n28 ^ n17 ;
  assign n30 = ~n16 & n29 ;
  assign n31 = ~x3 & ~n30 ;
  assign n33 = x5 & ~x7 ;
  assign n34 = x3 & n33 ;
  assign n32 = ~x0 & ~x1 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = n32 ^ n9 ;
  assign n37 = n34 ^ x2 ;
  assign n38 = n37 ^ n32 ;
  assign n39 = n32 & ~n38 ;
  assign n40 = n39 ^ n32 ;
  assign n41 = ~n36 & n40 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = n42 ^ n32 ;
  assign n44 = n43 ^ n37 ;
  assign n45 = n35 & ~n44 ;
  assign n46 = n45 ^ n34 ;
  assign n47 = ~x4 & ~n46 ;
  assign n48 = ~n31 & n47 ;
  assign n49 = ~n9 & ~n33 ;
  assign n50 = n10 ^ x3 ;
  assign n51 = n49 & ~n50 ;
  assign n52 = n51 ^ x3 ;
  assign n53 = ~x2 & ~n52 ;
  assign n54 = ~x1 & n53 ;
  assign n67 = ~x0 & x1 ;
  assign n65 = x2 & x5 ;
  assign n55 = x7 ^ x1 ;
  assign n56 = x7 ^ x3 ;
  assign n57 = x7 & n19 ;
  assign n58 = n57 ^ x7 ;
  assign n59 = n56 & n58 ;
  assign n60 = n59 ^ n57 ;
  assign n61 = n60 ^ x7 ;
  assign n62 = n61 ^ x0 ;
  assign n63 = ~n55 & n62 ;
  assign n64 = x5 & ~n63 ;
  assign n66 = n65 ^ n64 ;
  assign n68 = n67 ^ n66 ;
  assign n69 = n68 ^ n64 ;
  assign n75 = n69 ^ n66 ;
  assign n76 = n75 ^ n64 ;
  assign n77 = n76 ^ n64 ;
  assign n78 = ~x3 & ~x7 ;
  assign n79 = n78 ^ n66 ;
  assign n80 = n79 ^ n66 ;
  assign n81 = n80 ^ n64 ;
  assign n82 = ~n77 & ~n81 ;
  assign n70 = x2 & x3 ;
  assign n71 = n70 ^ n66 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = n72 ^ n64 ;
  assign n74 = n69 & n73 ;
  assign n83 = n82 ^ n74 ;
  assign n84 = n83 ^ n69 ;
  assign n85 = n74 ^ n64 ;
  assign n86 = n85 ^ n76 ;
  assign n87 = ~n64 & ~n86 ;
  assign n88 = n87 ^ n74 ;
  assign n89 = n84 & n88 ;
  assign n90 = n89 ^ n82 ;
  assign n91 = n90 ^ n87 ;
  assign n92 = n91 ^ n69 ;
  assign n93 = n92 ^ n64 ;
  assign n94 = n93 ^ n76 ;
  assign n95 = n94 ^ n65 ;
  assign n96 = x4 & n95 ;
  assign n97 = ~n54 & n96 ;
  assign n98 = ~n48 & ~n97 ;
  assign n99 = n98 ^ x6 ;
  assign n100 = n99 ^ n98 ;
  assign n126 = n56 ^ x2 ;
  assign n127 = n126 ^ x1 ;
  assign n128 = n127 ^ x7 ;
  assign n135 = n128 ^ n56 ;
  assign n129 = n128 ^ x5 ;
  assign n130 = n129 ^ n56 ;
  assign n131 = x5 ^ x1 ;
  assign n132 = n131 ^ x5 ;
  assign n133 = n132 ^ n130 ;
  assign n134 = ~n130 & ~n133 ;
  assign n136 = n135 ^ n134 ;
  assign n137 = n136 ^ n130 ;
  assign n138 = n56 ^ x7 ;
  assign n139 = n134 ^ n130 ;
  assign n140 = n138 & ~n139 ;
  assign n141 = n140 ^ n56 ;
  assign n142 = n137 & ~n141 ;
  assign n143 = n142 ^ n56 ;
  assign n144 = n143 ^ n56 ;
  assign n109 = x1 & ~x2 ;
  assign n110 = ~n78 & n109 ;
  assign n111 = ~n9 & n110 ;
  assign n101 = x1 & ~x7 ;
  assign n112 = ~x4 & ~n101 ;
  assign n113 = n112 ^ x3 ;
  assign n114 = n113 ^ n112 ;
  assign n115 = ~x1 & x5 ;
  assign n116 = n115 ^ n112 ;
  assign n117 = n114 & ~n116 ;
  assign n118 = n117 ^ n112 ;
  assign n119 = x2 & ~n118 ;
  assign n120 = ~n111 & ~n119 ;
  assign n121 = n78 & n115 ;
  assign n122 = x4 & ~n121 ;
  assign n123 = ~n120 & ~n122 ;
  assign n102 = ~x2 & ~x5 ;
  assign n103 = ~n70 & ~n102 ;
  assign n104 = n101 & ~n103 ;
  assign n105 = x3 & x5 ;
  assign n106 = ~x2 & n105 ;
  assign n107 = x7 & n106 ;
  assign n108 = ~n104 & ~n107 ;
  assign n124 = n123 ^ n108 ;
  assign n125 = n124 ^ n108 ;
  assign n145 = n144 ^ n125 ;
  assign n146 = n145 ^ n124 ;
  assign n147 = n124 ^ x4 ;
  assign n148 = n147 ^ n124 ;
  assign n149 = ~n146 & n148 ;
  assign n150 = n149 ^ n124 ;
  assign n151 = x0 & ~n150 ;
  assign n152 = n151 ^ n123 ;
  assign n153 = n70 ^ x4 ;
  assign n154 = n9 & n153 ;
  assign n155 = x1 & n154 ;
  assign n156 = ~n152 & ~n155 ;
  assign n157 = n156 ^ n98 ;
  assign n158 = ~n100 & ~n157 ;
  assign n159 = n158 ^ n98 ;
  assign n160 = ~n14 & ~n159 ;
  assign y0 = ~n160 ;
endmodule
