module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n9 = x5 ^ x3 ;
  assign n11 = n9 ^ x5 ;
  assign n12 = n11 ^ n9 ;
  assign n10 = n9 ^ x6 ;
  assign n13 = n12 ^ n10 ;
  assign n14 = n9 ^ x7 ;
  assign n15 = n14 ^ n9 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = ~n12 & ~n16 ;
  assign n18 = n17 ^ n12 ;
  assign n19 = n13 & ~n18 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n20 ^ n9 ;
  assign n22 = n21 ^ n12 ;
  assign n23 = ~x4 & ~n22 ;
  assign n24 = n23 ^ x3 ;
  assign y0 = ~n24 ;
endmodule
