module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 ;
  assign n9 = x4 & x6 ;
  assign n10 = x2 & x6 ;
  assign n11 = x5 & n10 ;
  assign n12 = ~n9 & ~n11 ;
  assign n13 = x2 & x4 ;
  assign n14 = x3 & ~n13 ;
  assign n15 = ~n12 & n14 ;
  assign n16 = ~x1 & n15 ;
  assign n17 = ~x3 & ~x4 ;
  assign n18 = n11 & n17 ;
  assign n19 = x5 & x7 ;
  assign n20 = ~x5 & ~x7 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = x2 & n21 ;
  assign n23 = ~x3 & ~x7 ;
  assign n24 = x3 & x7 ;
  assign n25 = x4 & ~n24 ;
  assign n26 = ~n23 & n25 ;
  assign n27 = ~n22 & ~n26 ;
  assign n28 = ~x6 & ~n27 ;
  assign n30 = x5 ^ x3 ;
  assign n29 = x4 ^ x2 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n29 ^ x4 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = ~n31 & ~n33 ;
  assign n35 = n34 ^ x4 ;
  assign n36 = n35 ^ n29 ;
  assign n37 = n36 ^ n31 ;
  assign n38 = n37 ^ x6 ;
  assign n39 = n29 ^ x6 ;
  assign n43 = x5 ^ x4 ;
  assign n44 = n43 ^ x4 ;
  assign n45 = n44 ^ n31 ;
  assign n46 = n44 & ~n45 ;
  assign n40 = n31 ^ x4 ;
  assign n41 = n20 ^ x4 ;
  assign n42 = n40 & n41 ;
  assign n47 = n46 ^ n42 ;
  assign n48 = n47 ^ n43 ;
  assign n49 = n48 ^ n20 ;
  assign n50 = n49 ^ x4 ;
  assign n51 = n50 ^ n31 ;
  assign n52 = n51 ^ x6 ;
  assign n53 = n39 & ~n52 ;
  assign n54 = n53 ^ n46 ;
  assign n55 = n54 ^ n43 ;
  assign n56 = n55 ^ n29 ;
  assign n57 = n56 ^ x6 ;
  assign n58 = n38 & ~n57 ;
  assign n59 = n58 ^ n46 ;
  assign n60 = n59 ^ n53 ;
  assign n61 = n60 ^ n43 ;
  assign n62 = n61 ^ n29 ;
  assign n63 = n62 ^ x6 ;
  assign n64 = ~n28 & n63 ;
  assign n65 = ~x3 & ~x5 ;
  assign n66 = n65 ^ x4 ;
  assign n67 = n29 & ~n66 ;
  assign n68 = n67 ^ x2 ;
  assign n69 = n64 & ~n68 ;
  assign n70 = n69 ^ x1 ;
  assign n71 = n70 ^ n69 ;
  assign n72 = n71 ^ n18 ;
  assign n73 = n17 & ~n21 ;
  assign n74 = ~x6 & n73 ;
  assign n75 = x3 & ~n19 ;
  assign n76 = ~x6 & x7 ;
  assign n77 = ~x4 & x5 ;
  assign n78 = ~n76 & ~n77 ;
  assign n79 = n75 & ~n78 ;
  assign n80 = x6 ^ x4 ;
  assign n81 = ~x5 & n23 ;
  assign n82 = n81 ^ x6 ;
  assign n83 = n80 & n82 ;
  assign n84 = n83 ^ x4 ;
  assign n85 = ~n79 & n84 ;
  assign n86 = ~x2 & ~n85 ;
  assign n87 = n86 ^ n74 ;
  assign n88 = ~n74 & n87 ;
  assign n89 = n88 ^ n69 ;
  assign n90 = n89 ^ n74 ;
  assign n91 = ~n72 & n90 ;
  assign n92 = n91 ^ n88 ;
  assign n93 = n92 ^ n74 ;
  assign n94 = ~n18 & ~n93 ;
  assign n95 = n94 ^ n18 ;
  assign n96 = n95 ^ x0 ;
  assign n97 = n96 ^ n95 ;
  assign n98 = ~x5 & ~x6 ;
  assign n99 = x3 & ~n98 ;
  assign n100 = x7 ^ x1 ;
  assign n101 = n100 ^ x7 ;
  assign n102 = ~n65 & ~n76 ;
  assign n103 = n102 ^ x7 ;
  assign n104 = ~n101 & n103 ;
  assign n105 = n104 ^ x7 ;
  assign n106 = ~n99 & n105 ;
  assign n107 = n13 & ~n106 ;
  assign n108 = ~x2 & ~x3 ;
  assign n109 = n19 & n108 ;
  assign n110 = ~x1 & ~n109 ;
  assign n111 = ~n20 & n110 ;
  assign n112 = n9 & ~n75 ;
  assign n113 = ~n111 & n112 ;
  assign n114 = x5 ^ x1 ;
  assign n115 = n114 ^ x4 ;
  assign n116 = n115 ^ x4 ;
  assign n121 = x7 ^ x5 ;
  assign n117 = x4 ^ x3 ;
  assign n118 = n117 ^ x1 ;
  assign n122 = n121 ^ n118 ;
  assign n123 = n122 ^ x4 ;
  assign n124 = ~x4 & n123 ;
  assign n119 = x5 & n118 ;
  assign n127 = n124 ^ n119 ;
  assign n120 = n119 ^ n116 ;
  assign n125 = n124 ^ x4 ;
  assign n126 = n120 & ~n125 ;
  assign n128 = n127 ^ n126 ;
  assign n129 = n116 & n128 ;
  assign n130 = n129 ^ n124 ;
  assign n131 = n130 ^ n126 ;
  assign n132 = n131 ^ x4 ;
  assign n133 = n10 & ~n132 ;
  assign n134 = ~n113 & ~n133 ;
  assign n135 = ~n107 & n134 ;
  assign n136 = n135 ^ n95 ;
  assign n137 = ~n97 & ~n136 ;
  assign n138 = n137 ^ n95 ;
  assign n139 = ~n16 & ~n138 ;
  assign y0 = ~n139 ;
endmodule
