// Benchmark "./newcwp.pla" written by ABC on Thu Apr 23 10:59:58 2020

module \./newcwp.pla  ( 
    x0, x1, x2, x3,
    z1  );
  input  x0, x1, x2, x3;
  output z1;
  assign z1 = 1'b1;
endmodule


