module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 ;
  assign n9 = x0 & ~x1 ;
  assign n10 = x3 & x4 ;
  assign n11 = x5 & x7 ;
  assign n12 = x2 & ~n11 ;
  assign n13 = n10 & ~n12 ;
  assign n15 = x7 ^ x6 ;
  assign n14 = x7 ^ x5 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n14 ^ x7 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = x2 & n19 ;
  assign n21 = n20 ^ n14 ;
  assign n22 = n21 ^ x2 ;
  assign n23 = ~n17 & n22 ;
  assign n24 = n23 ^ n20 ;
  assign n25 = n24 ^ x2 ;
  assign n26 = n13 & n25 ;
  assign n27 = n9 & ~n26 ;
  assign n28 = x7 ^ x3 ;
  assign n29 = ~x1 & x6 ;
  assign n30 = n29 ^ x7 ;
  assign n31 = n30 ^ x2 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = n32 ^ n28 ;
  assign n34 = ~x0 & x1 ;
  assign n35 = n34 ^ x2 ;
  assign n36 = ~x2 & ~n35 ;
  assign n37 = n36 ^ n29 ;
  assign n38 = n37 ^ x2 ;
  assign n39 = ~n33 & ~n38 ;
  assign n40 = n39 ^ n36 ;
  assign n41 = n40 ^ x2 ;
  assign n42 = ~n28 & ~n41 ;
  assign n43 = ~x4 & n42 ;
  assign n44 = n10 & n34 ;
  assign n45 = ~x2 & x6 ;
  assign n46 = ~x2 & ~x7 ;
  assign n47 = ~n45 & ~n46 ;
  assign n48 = n44 & n47 ;
  assign n49 = ~x3 & n46 ;
  assign n50 = ~x4 & ~x6 ;
  assign n51 = x0 & n50 ;
  assign n52 = n49 & n51 ;
  assign n53 = ~n48 & ~n52 ;
  assign n54 = ~n43 & n53 ;
  assign n55 = x5 & ~n54 ;
  assign n56 = x2 & n34 ;
  assign n57 = x4 ^ x3 ;
  assign n58 = n57 ^ x6 ;
  assign n59 = x6 ^ x4 ;
  assign n60 = ~x5 & x7 ;
  assign n61 = n60 ^ x4 ;
  assign n62 = n59 & n61 ;
  assign n63 = n62 ^ x4 ;
  assign n64 = n58 & n63 ;
  assign n65 = n56 & n64 ;
  assign n66 = ~n55 & ~n65 ;
  assign n67 = ~n27 & n66 ;
  assign y0 = ~n67 ;
endmodule
