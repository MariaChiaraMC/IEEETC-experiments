// Benchmark "./pla/max128.pla_dbb_orig_18NonExact" written by ABC on Fri Nov 20 10:25:27 2020

module \./pla/max128.pla_dbb_orig_18NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = 1'b1;
endmodule


