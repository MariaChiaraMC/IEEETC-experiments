module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 ;
  assign n10 = x5 ^ x0 ;
  assign n11 = n10 ^ x1 ;
  assign n12 = n11 ^ x3 ;
  assign n13 = n12 ^ x5 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n14 ^ n10 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = ~x3 & ~n16 ;
  assign n18 = n17 ^ n12 ;
  assign n19 = ~x6 & ~x7 ;
  assign n20 = n19 ^ n12 ;
  assign n21 = n15 & n20 ;
  assign n22 = n21 ^ n14 ;
  assign n23 = n22 ^ n15 ;
  assign n24 = ~n18 & ~n23 ;
  assign n25 = ~n14 & n24 ;
  assign n26 = n25 ^ n17 ;
  assign n27 = n26 ^ x0 ;
  assign n28 = x2 & n27 ;
  assign n29 = ~x1 & x3 ;
  assign n30 = n29 ^ x0 ;
  assign n31 = x6 & x7 ;
  assign n32 = x2 & n31 ;
  assign n33 = x3 & x5 ;
  assign n34 = ~n32 & n33 ;
  assign n35 = x1 & n34 ;
  assign n36 = n35 ^ n30 ;
  assign n37 = x2 ^ x0 ;
  assign n38 = n37 ^ x2 ;
  assign n39 = x3 & x6 ;
  assign n40 = x6 ^ x2 ;
  assign n41 = ~x5 & ~n40 ;
  assign n42 = n41 ^ x2 ;
  assign n43 = ~x1 & ~n42 ;
  assign n44 = ~n39 & ~n43 ;
  assign n45 = n44 ^ x2 ;
  assign n46 = n38 & n45 ;
  assign n47 = n46 ^ x2 ;
  assign n48 = n47 ^ n30 ;
  assign n49 = ~n36 & ~n48 ;
  assign n50 = n49 ^ n46 ;
  assign n51 = n50 ^ x2 ;
  assign n52 = n51 ^ n35 ;
  assign n53 = n30 & n52 ;
  assign n54 = n53 ^ n30 ;
  assign n55 = n54 ^ n35 ;
  assign n56 = ~n28 & ~n55 ;
  assign n57 = x4 & ~n56 ;
  assign n58 = ~x0 & ~x2 ;
  assign n59 = x1 & ~x3 ;
  assign n60 = x5 & n31 ;
  assign n61 = n59 & ~n60 ;
  assign n62 = x5 & x6 ;
  assign n63 = n29 & n62 ;
  assign n64 = ~n61 & ~n63 ;
  assign n65 = n58 & ~n64 ;
  assign n66 = ~n57 & ~n65 ;
  assign n67 = x4 ^ x0 ;
  assign n68 = ~x1 & ~x6 ;
  assign n69 = n68 ^ x0 ;
  assign n70 = ~x5 & ~x6 ;
  assign n71 = ~x7 & ~x8 ;
  assign n72 = n70 & n71 ;
  assign n73 = n72 ^ x0 ;
  assign n74 = ~x0 & n73 ;
  assign n75 = n74 ^ x0 ;
  assign n76 = ~n69 & ~n75 ;
  assign n77 = n76 ^ n74 ;
  assign n78 = n77 ^ x0 ;
  assign n79 = n78 ^ n72 ;
  assign n80 = n67 & n79 ;
  assign n81 = n80 ^ x0 ;
  assign n82 = ~x3 & ~n81 ;
  assign n83 = ~x4 & x5 ;
  assign n84 = ~x0 & ~n83 ;
  assign n85 = x1 & ~n84 ;
  assign n86 = ~n82 & ~n85 ;
  assign n87 = x2 & ~n86 ;
  assign n88 = n29 & n58 ;
  assign n89 = x5 & x7 ;
  assign n90 = n88 & n89 ;
  assign n91 = n90 ^ x4 ;
  assign n92 = n91 ^ x8 ;
  assign n106 = n92 ^ n59 ;
  assign n93 = n92 ^ n90 ;
  assign n94 = n93 ^ n92 ;
  assign n105 = n94 ^ n59 ;
  assign n107 = n106 ^ n105 ;
  assign n96 = x0 & ~x2 ;
  assign n97 = n29 & n96 ;
  assign n98 = ~n62 & ~n89 ;
  assign n99 = n97 & n98 ;
  assign n100 = n99 ^ n93 ;
  assign n95 = n94 ^ n91 ;
  assign n101 = n100 ^ n95 ;
  assign n102 = n95 ^ n59 ;
  assign n103 = ~n101 & n102 ;
  assign n104 = n103 ^ n59 ;
  assign n108 = n107 ^ n104 ;
  assign n109 = n108 ^ n100 ;
  assign n110 = n107 ^ n106 ;
  assign n111 = n110 ^ n95 ;
  assign n112 = ~n106 & n111 ;
  assign n113 = x0 & x5 ;
  assign n114 = n31 & n113 ;
  assign n115 = n106 ^ n100 ;
  assign n116 = ~n114 & ~n115 ;
  assign n117 = n116 ^ n114 ;
  assign n118 = n117 ^ n100 ;
  assign n119 = n118 ^ n95 ;
  assign n120 = n112 & n119 ;
  assign n121 = n120 ^ n59 ;
  assign n122 = ~n109 & ~n121 ;
  assign n123 = n122 ^ n112 ;
  assign n124 = n123 ^ n120 ;
  assign n125 = n124 ^ n59 ;
  assign n126 = n125 ^ n106 ;
  assign n127 = n126 ^ n107 ;
  assign n128 = n127 ^ x4 ;
  assign n129 = n128 ^ n94 ;
  assign n130 = ~n87 & n129 ;
  assign n131 = n66 & n130 ;
  assign y0 = ~n131 ;
endmodule
