module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 ;
  assign n72 = x9 & ~x13 ;
  assign n73 = x10 & n72 ;
  assign n16 = x10 ^ x9 ;
  assign n17 = n16 ^ x10 ;
  assign n18 = n17 ^ x13 ;
  assign n19 = n18 ^ n16 ;
  assign n27 = n19 ^ n16 ;
  assign n28 = n27 ^ n17 ;
  assign n20 = ~x3 & x4 ;
  assign n21 = ~x2 & x13 ;
  assign n22 = ~n20 & n21 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = n23 ^ n19 ;
  assign n25 = n24 ^ n16 ;
  assign n26 = n25 ^ n17 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = ~n17 & ~n29 ;
  assign n31 = n30 ^ n19 ;
  assign n32 = n31 ^ n28 ;
  assign n48 = ~x2 & ~x3 ;
  assign n49 = x0 & ~x1 ;
  assign n54 = ~n48 & n49 ;
  assign n55 = x14 & ~n54 ;
  assign n59 = n55 ^ n16 ;
  assign n33 = x0 & x3 ;
  assign n34 = x4 & ~x5 ;
  assign n35 = x2 & n34 ;
  assign n36 = x0 & ~n35 ;
  assign n37 = ~n33 & ~n36 ;
  assign n38 = x6 ^ x2 ;
  assign n39 = ~x1 & n38 ;
  assign n40 = n39 ^ x2 ;
  assign n41 = n37 & ~n40 ;
  assign n42 = x1 & x2 ;
  assign n43 = n33 & n42 ;
  assign n44 = x6 ^ x4 ;
  assign n45 = x5 & ~n44 ;
  assign n46 = n45 ^ x4 ;
  assign n47 = n43 & n46 ;
  assign n50 = n48 & n49 ;
  assign n51 = x5 & n50 ;
  assign n52 = ~n47 & ~n51 ;
  assign n53 = ~n41 & n52 ;
  assign n56 = n55 ^ n53 ;
  assign n57 = n28 ^ n19 ;
  assign n58 = ~n56 & n57 ;
  assign n60 = n59 ^ n58 ;
  assign n61 = n60 ^ n56 ;
  assign n62 = n61 ^ n17 ;
  assign n63 = n31 & ~n62 ;
  assign n64 = n63 ^ n19 ;
  assign n65 = n64 ^ n17 ;
  assign n66 = n65 ^ n28 ;
  assign n67 = n32 & ~n66 ;
  assign n68 = n67 ^ n19 ;
  assign n69 = n68 ^ n17 ;
  assign n70 = n69 ^ n28 ;
  assign n71 = n70 ^ x10 ;
  assign n74 = n73 ^ n71 ;
  assign n75 = ~x11 & ~n74 ;
  assign n76 = n75 ^ n73 ;
  assign y0 = n76 ;
endmodule
