module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 ;
  assign n9 = x6 ^ x4 ;
  assign n10 = n9 ^ x5 ;
  assign n11 = x2 & x7 ;
  assign n12 = ~x1 & ~n11 ;
  assign n13 = n12 ^ x2 ;
  assign n14 = x4 & n13 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n10 & ~n15 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = n17 ^ n12 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = x5 & ~n19 ;
  assign n21 = x2 ^ x1 ;
  assign n22 = n21 ^ x2 ;
  assign n23 = n22 ^ x5 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n24 ^ n23 ;
  assign n28 = n21 ^ x6 ;
  assign n26 = n23 ^ x7 ;
  assign n27 = n26 ^ n24 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = ~n25 & n29 ;
  assign n31 = n30 ^ n25 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = n25 ^ n21 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = n33 ^ n23 ;
  assign n36 = n34 & ~n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ n27 ;
  assign n39 = n38 ^ n23 ;
  assign n40 = n34 ^ n23 ;
  assign n41 = n21 ^ x4 ;
  assign n42 = n41 ^ n25 ;
  assign n43 = n42 ^ n33 ;
  assign n44 = ~n40 & n43 ;
  assign n45 = n44 ^ n41 ;
  assign n46 = n45 ^ n33 ;
  assign n47 = n46 ^ n27 ;
  assign n48 = n47 ^ n23 ;
  assign n49 = ~n39 & n48 ;
  assign n50 = n49 ^ n23 ;
  assign n51 = ~n32 & ~n50 ;
  assign n52 = n51 ^ n36 ;
  assign n53 = n52 ^ n33 ;
  assign n54 = n53 ^ n27 ;
  assign n55 = n54 ^ n23 ;
  assign n56 = n55 ^ x1 ;
  assign n57 = n56 ^ n23 ;
  assign n58 = ~n20 & ~n57 ;
  assign y0 = n58 ;
endmodule
