module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n7 = ~x3 & x4 ;
  assign n8 = ~x2 & ~n7 ;
  assign n9 = x2 ^ x1 ;
  assign n10 = x5 ^ x3 ;
  assign n11 = x3 ^ x2 ;
  assign n12 = n11 ^ x3 ;
  assign n13 = ~n10 & ~n12 ;
  assign n14 = n13 ^ x3 ;
  assign n15 = ~n9 & ~n14 ;
  assign n16 = n15 ^ x1 ;
  assign n17 = x0 & n16 ;
  assign n18 = ~n8 & n17 ;
  assign n19 = ~x0 & ~x2 ;
  assign n20 = x5 ^ x4 ;
  assign n21 = n20 ^ n10 ;
  assign n22 = n10 ^ x1 ;
  assign n23 = n10 & ~n22 ;
  assign n24 = n23 ^ n10 ;
  assign n25 = ~n21 & n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n26 ^ n10 ;
  assign n28 = n27 ^ x1 ;
  assign n29 = n19 & ~n28 ;
  assign n30 = ~n18 & ~n29 ;
  assign y0 = ~n30 ;
endmodule
