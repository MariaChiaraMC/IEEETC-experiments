module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 ;
  assign n31 = x7 & x8 ;
  assign n32 = x3 & ~n31 ;
  assign n33 = x5 & ~n32 ;
  assign n34 = x12 & ~x13 ;
  assign n35 = ~x9 & n34 ;
  assign n36 = ~x6 & n35 ;
  assign n37 = ~n33 & n36 ;
  assign n38 = ~x2 & x3 ;
  assign n39 = ~x5 & ~n38 ;
  assign n40 = ~x4 & ~n39 ;
  assign n41 = ~x7 & ~x8 ;
  assign n42 = ~x10 & ~x11 ;
  assign n43 = ~n41 & n42 ;
  assign n44 = ~x0 & n43 ;
  assign n45 = ~n40 & n44 ;
  assign n46 = n37 & n45 ;
  assign n17 = x4 ^ x2 ;
  assign n18 = n17 ^ x4 ;
  assign n15 = x4 ^ x3 ;
  assign n16 = n15 ^ x4 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = x5 ^ x4 ;
  assign n21 = n20 ^ x4 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = n18 & n22 ;
  assign n24 = n23 ^ n18 ;
  assign n25 = n19 & n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n26 ^ x4 ;
  assign n28 = n27 ^ n18 ;
  assign n29 = ~x0 & n28 ;
  assign n30 = n29 ^ x4 ;
  assign n47 = n46 ^ n30 ;
  assign n48 = x1 & n47 ;
  assign n49 = n48 ^ n30 ;
  assign y0 = n49 ;
endmodule
