module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n24 = x8 ^ x4 ;
  assign n25 = ~x0 & n24 ;
  assign n26 = n25 ^ x4 ;
  assign n28 = n26 ^ x3 ;
  assign n27 = n26 ^ x7 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n28 ^ x0 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n29 & ~n31 ;
  assign n33 = n32 ^ n28 ;
  assign n34 = x2 & n33 ;
  assign n35 = n34 ^ n26 ;
  assign n12 = x10 ^ x6 ;
  assign n13 = ~x0 & n12 ;
  assign n14 = n13 ^ x6 ;
  assign n16 = n14 ^ x5 ;
  assign n15 = n14 ^ x9 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n16 ^ x0 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n17 & ~n19 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = x2 & n21 ;
  assign n23 = n22 ^ n14 ;
  assign n36 = n35 ^ n23 ;
  assign n37 = ~x1 & n36 ;
  assign n38 = n37 ^ n35 ;
  assign y0 = n38 ;
endmodule
