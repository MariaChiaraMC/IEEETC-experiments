// Benchmark "./pla/ryy6.pla_dbb_orig_0NonExact" written by ABC on Fri Nov 20 10:28:15 2020

module \./pla/ryy6.pla_dbb_orig_0NonExact  ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15,
    z0  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15;
  output z0;
  wire new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_, new_n24_,
    new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_, new_n31_,
    new_n32_;
  assign new_n18_ = x10 & x11;
  assign new_n19_ = x07 & x08;
  assign new_n20_ = ~new_n18_ & ~new_n19_;
  assign new_n21_ = x02 & x09;
  assign new_n22_ = ~new_n20_ & new_n21_;
  assign new_n23_ = x05 & x06;
  assign new_n24_ = x03 & x04;
  assign new_n25_ = ~new_n23_ & ~new_n24_;
  assign new_n26_ = ~new_n22_ & new_n25_;
  assign new_n27_ = ~x00 & ~x02;
  assign new_n28_ = x01 & ~new_n27_;
  assign new_n29_ = x14 & x15;
  assign new_n30_ = x13 & new_n29_;
  assign new_n31_ = x12 & new_n30_;
  assign new_n32_ = ~new_n28_ & ~new_n31_;
  assign z0 = new_n26_ & new_n32_;
endmodule


