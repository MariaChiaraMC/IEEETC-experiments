module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 ;
  assign n16 = ~x4 & ~x6 ;
  assign n17 = x4 & x6 ;
  assign n18 = ~n16 & ~n17 ;
  assign n19 = ~x0 & x14 ;
  assign n20 = x9 & ~x11 ;
  assign n21 = ~x9 & x11 ;
  assign n22 = ~n20 & ~n21 ;
  assign n23 = x8 & ~x10 ;
  assign n24 = x2 & ~x12 ;
  assign n25 = x3 & ~x7 ;
  assign n26 = x5 & n25 ;
  assign n29 = x7 & ~x13 ;
  assign n27 = ~x1 & ~x3 ;
  assign n28 = ~x5 & n27 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n31 ^ n26 ;
  assign n33 = ~x7 & x13 ;
  assign n34 = x1 & ~x5 ;
  assign n35 = ~x3 & n34 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = ~n33 & ~n36 ;
  assign n38 = n37 ^ n28 ;
  assign n39 = n38 ^ n33 ;
  assign n40 = n32 & ~n39 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n41 ^ n33 ;
  assign n43 = ~n26 & ~n42 ;
  assign n44 = n43 ^ n26 ;
  assign n45 = n24 & n44 ;
  assign n46 = n23 & n45 ;
  assign n47 = x5 & x13 ;
  assign n48 = x1 & ~x7 ;
  assign n49 = ~n47 & n48 ;
  assign n50 = ~x3 & ~n49 ;
  assign n51 = x7 & x13 ;
  assign n52 = ~x1 & x5 ;
  assign n53 = n51 & n52 ;
  assign n54 = ~x3 & ~n47 ;
  assign n55 = ~x5 & ~x13 ;
  assign n56 = ~n54 & ~n55 ;
  assign n57 = n48 & ~n56 ;
  assign n58 = ~n53 & ~n57 ;
  assign n59 = x10 & x12 ;
  assign n60 = x2 & ~x8 ;
  assign n61 = n59 & n60 ;
  assign n62 = ~n58 & n61 ;
  assign n63 = ~n50 & n62 ;
  assign n64 = x3 & x12 ;
  assign n65 = ~x2 & x10 ;
  assign n66 = n64 & n65 ;
  assign n67 = n48 & n66 ;
  assign n68 = n47 & n67 ;
  assign n69 = ~x1 & ~x2 ;
  assign n70 = x7 & x10 ;
  assign n71 = x12 & n70 ;
  assign n72 = n69 & n71 ;
  assign n73 = ~n56 & n72 ;
  assign n74 = ~n68 & ~n73 ;
  assign n75 = x8 & ~n74 ;
  assign n76 = ~n63 & ~n75 ;
  assign n77 = ~n46 & n76 ;
  assign n78 = ~n22 & ~n77 ;
  assign n79 = ~x10 & x12 ;
  assign n80 = x10 & ~x12 ;
  assign n81 = ~n79 & ~n80 ;
  assign n82 = x8 & ~x9 ;
  assign n83 = ~x11 & n82 ;
  assign n84 = x3 & x5 ;
  assign n85 = n51 & n69 ;
  assign n86 = ~x7 & ~x13 ;
  assign n87 = x1 & x2 ;
  assign n88 = n86 & n87 ;
  assign n89 = ~n85 & ~n88 ;
  assign n90 = n84 & ~n89 ;
  assign n91 = ~x3 & ~x5 ;
  assign n92 = n87 & n91 ;
  assign n93 = ~n33 & n92 ;
  assign n94 = ~n90 & ~n93 ;
  assign n95 = n83 & ~n94 ;
  assign n96 = x9 & ~n95 ;
  assign n97 = x11 & n84 ;
  assign n98 = ~x8 & x13 ;
  assign n99 = ~x2 & ~x7 ;
  assign n100 = x2 & x7 ;
  assign n101 = ~n99 & ~n100 ;
  assign n102 = n98 & ~n101 ;
  assign n103 = n97 & n102 ;
  assign n104 = n103 ^ n95 ;
  assign n105 = x8 & x11 ;
  assign n106 = ~x2 & x3 ;
  assign n107 = n47 & n106 ;
  assign n108 = x2 & ~x3 ;
  assign n109 = n55 & n108 ;
  assign n110 = ~n107 & ~n109 ;
  assign n111 = n48 & ~n110 ;
  assign n112 = ~x1 & x7 ;
  assign n113 = x13 ^ x2 ;
  assign n114 = n112 & n113 ;
  assign n115 = n91 & n114 ;
  assign n116 = ~n111 & ~n115 ;
  assign n117 = n105 & ~n116 ;
  assign n118 = n117 ^ n96 ;
  assign n119 = n104 & n118 ;
  assign n120 = n119 ^ n117 ;
  assign n121 = n96 & n120 ;
  assign n122 = n121 ^ n95 ;
  assign n123 = ~n81 & n122 ;
  assign n124 = ~x8 & x10 ;
  assign n125 = ~x5 & ~x7 ;
  assign n126 = n124 & n125 ;
  assign n127 = x12 & ~x13 ;
  assign n128 = ~x2 & ~x3 ;
  assign n129 = x1 & ~x11 ;
  assign n130 = n128 & n129 ;
  assign n131 = n127 & n130 ;
  assign n132 = n126 & n131 ;
  assign n133 = ~n123 & ~n132 ;
  assign n134 = x1 & ~x12 ;
  assign n148 = x8 & ~x11 ;
  assign n135 = ~x8 & x11 ;
  assign n136 = n70 & n91 ;
  assign n137 = ~x10 & x13 ;
  assign n138 = n26 & n137 ;
  assign n139 = ~n136 & ~n138 ;
  assign n140 = n135 & ~n139 ;
  assign n149 = n148 ^ n140 ;
  assign n150 = n149 ^ n140 ;
  assign n141 = ~x3 & x5 ;
  assign n142 = x3 & ~x5 ;
  assign n143 = ~n141 & ~n142 ;
  assign n144 = ~x5 & x13 ;
  assign n145 = n143 & ~n144 ;
  assign n146 = n145 ^ n140 ;
  assign n147 = n146 ^ n140 ;
  assign n151 = n150 ^ n147 ;
  assign n152 = ~x7 & x10 ;
  assign n153 = n152 ^ n140 ;
  assign n154 = n153 ^ n140 ;
  assign n155 = n154 ^ n150 ;
  assign n156 = n150 & n155 ;
  assign n157 = n156 ^ n150 ;
  assign n158 = n151 & n157 ;
  assign n159 = n158 ^ n156 ;
  assign n160 = n159 ^ n140 ;
  assign n161 = n160 ^ n150 ;
  assign n162 = ~x2 & n161 ;
  assign n163 = n162 ^ n140 ;
  assign n164 = n134 & n163 ;
  assign n165 = ~n48 & ~n112 ;
  assign n166 = ~x2 & x12 ;
  assign n167 = ~x9 & x10 ;
  assign n168 = ~x8 & n167 ;
  assign n169 = n166 & n168 ;
  assign n170 = x9 & x12 ;
  assign n171 = ~x9 & ~x12 ;
  assign n172 = ~n170 & ~n171 ;
  assign n173 = ~x11 & x13 ;
  assign n174 = x2 & x8 ;
  assign n175 = ~x10 & n174 ;
  assign n176 = n173 & n175 ;
  assign n177 = ~n172 & n176 ;
  assign n178 = ~n169 & ~n177 ;
  assign n179 = n84 & ~n178 ;
  assign n180 = ~x3 & ~x13 ;
  assign n181 = ~x2 & ~x9 ;
  assign n182 = ~x5 & x11 ;
  assign n183 = n181 & n182 ;
  assign n184 = n180 & n183 ;
  assign n185 = n124 & n184 ;
  assign n186 = ~n179 & ~n185 ;
  assign n187 = ~n165 & ~n186 ;
  assign n188 = ~n164 & ~n187 ;
  assign n189 = n52 & n106 ;
  assign n190 = ~x7 & x8 ;
  assign n191 = x10 & x11 ;
  assign n192 = ~x12 & n191 ;
  assign n193 = n190 & n192 ;
  assign n194 = n189 & n193 ;
  assign n195 = n188 & ~n194 ;
  assign n196 = n133 & n195 ;
  assign n218 = x2 & x3 ;
  assign n219 = x5 & n218 ;
  assign n300 = ~x11 & ~x12 ;
  assign n301 = n124 & n300 ;
  assign n302 = n219 & n301 ;
  assign n303 = ~n24 & ~n166 ;
  assign n304 = ~x1 & ~n303 ;
  assign n305 = x10 & ~x11 ;
  assign n306 = ~x13 & n305 ;
  assign n307 = ~x5 & x8 ;
  assign n308 = ~x3 & n307 ;
  assign n309 = n306 & n308 ;
  assign n310 = n304 & n309 ;
  assign n311 = ~n302 & ~n310 ;
  assign n312 = x5 & x8 ;
  assign n313 = ~x5 & ~x8 ;
  assign n314 = ~n312 & ~n313 ;
  assign n315 = ~x3 & ~n314 ;
  assign n316 = x3 & x8 ;
  assign n317 = ~x5 & n316 ;
  assign n318 = ~n315 & ~n317 ;
  assign n319 = n127 & ~n318 ;
  assign n265 = x8 & ~x12 ;
  assign n320 = n47 ^ x3 ;
  assign n321 = n320 ^ n47 ;
  assign n322 = x5 & ~x13 ;
  assign n323 = ~n144 & ~n322 ;
  assign n324 = n323 ^ n47 ;
  assign n325 = n321 & ~n324 ;
  assign n326 = n325 ^ n47 ;
  assign n327 = n265 & n326 ;
  assign n328 = ~n319 & ~n327 ;
  assign n329 = ~x10 & ~x11 ;
  assign n330 = n87 & n329 ;
  assign n331 = ~n328 & n330 ;
  assign n332 = n311 & ~n331 ;
  assign n333 = x1 & ~x2 ;
  assign n334 = ~x8 & n91 ;
  assign n335 = x10 & ~x13 ;
  assign n336 = n334 & n335 ;
  assign n337 = n23 & n84 ;
  assign n338 = n173 & n337 ;
  assign n339 = ~n336 & ~n338 ;
  assign n340 = n339 ^ x12 ;
  assign n341 = n340 ^ n339 ;
  assign n342 = n341 ^ n333 ;
  assign n343 = ~x10 & x11 ;
  assign n344 = x11 & ~x13 ;
  assign n345 = ~n343 & ~n344 ;
  assign n346 = ~x8 & ~x11 ;
  assign n281 = x8 & x10 ;
  assign n347 = n84 & ~n281 ;
  assign n348 = ~n346 & n347 ;
  assign n349 = n345 & n348 ;
  assign n350 = n191 & n334 ;
  assign n351 = n350 ^ n349 ;
  assign n352 = ~n349 & n351 ;
  assign n353 = n352 ^ n339 ;
  assign n354 = n353 ^ n349 ;
  assign n355 = n342 & ~n354 ;
  assign n356 = n355 ^ n352 ;
  assign n357 = n356 ^ n349 ;
  assign n358 = n333 & ~n357 ;
  assign n359 = n358 ^ n333 ;
  assign n360 = n332 & ~n359 ;
  assign n361 = x7 & ~n360 ;
  assign n362 = x11 & x13 ;
  assign n363 = ~x2 & ~n362 ;
  assign n364 = ~n87 & ~n363 ;
  assign n249 = x5 & ~x12 ;
  assign n365 = ~n105 & n249 ;
  assign n366 = x7 & ~x10 ;
  assign n367 = ~n300 & n366 ;
  assign n368 = ~n365 & n367 ;
  assign n253 = ~x2 & ~x12 ;
  assign n369 = x8 & ~n253 ;
  assign n370 = ~x11 & n127 ;
  assign n371 = n369 & ~n370 ;
  assign n372 = n145 & ~n371 ;
  assign n373 = n368 & n372 ;
  assign n374 = n364 & n373 ;
  assign n375 = ~n361 & ~n374 ;
  assign n376 = n60 & n192 ;
  assign n377 = ~x12 & x13 ;
  assign n378 = n191 & n377 ;
  assign n379 = ~x2 & ~x10 ;
  assign n380 = ~n378 & ~n379 ;
  assign n381 = n369 & ~n380 ;
  assign n382 = x1 & n381 ;
  assign n383 = ~n376 & ~n382 ;
  assign n384 = n26 & ~n383 ;
  assign n385 = ~x11 & ~x13 ;
  assign n386 = n91 & n385 ;
  assign n387 = n124 & n304 ;
  assign n288 = ~x2 & n23 ;
  assign n388 = x1 & x12 ;
  assign n389 = n288 & n388 ;
  assign n390 = ~n387 & ~n389 ;
  assign n391 = n386 & ~n390 ;
  assign n392 = ~n384 & ~n391 ;
  assign n393 = n375 & n392 ;
  assign n197 = x5 & ~x7 ;
  assign n198 = n106 & n197 ;
  assign n199 = x8 & ~x13 ;
  assign n200 = n79 & n199 ;
  assign n201 = n198 & n200 ;
  assign n202 = ~x7 & ~x8 ;
  assign n203 = x2 & ~x10 ;
  assign n204 = n145 & n203 ;
  assign n205 = x5 & x10 ;
  assign n206 = x3 & n205 ;
  assign n207 = ~x2 & n206 ;
  assign n208 = ~n204 & ~n207 ;
  assign n209 = n202 & ~n208 ;
  assign n210 = x12 & n209 ;
  assign n211 = n107 & n124 ;
  assign n212 = ~x5 & n108 ;
  assign n213 = n200 & n212 ;
  assign n214 = ~n211 & ~n213 ;
  assign n215 = x7 & ~n214 ;
  assign n216 = n55 & n128 ;
  assign n217 = n79 & n216 ;
  assign n220 = ~x7 & ~x12 ;
  assign n221 = x13 ^ x10 ;
  assign n222 = n220 & n221 ;
  assign n223 = n219 & n222 ;
  assign n224 = ~n217 & ~n223 ;
  assign n225 = ~x8 & ~n224 ;
  assign n226 = ~n215 & ~n225 ;
  assign n227 = ~n210 & n226 ;
  assign n228 = ~n201 & n227 ;
  assign n229 = n129 & ~n228 ;
  assign n230 = ~x8 & ~x10 ;
  assign n231 = ~x12 & ~x13 ;
  assign n232 = n230 & n231 ;
  assign n233 = n112 & n232 ;
  assign n234 = n233 ^ x1 ;
  assign n235 = n234 ^ n233 ;
  assign n236 = ~x10 & ~x12 ;
  assign n237 = ~x13 & n236 ;
  assign n238 = n190 & n237 ;
  assign n239 = ~x8 & n71 ;
  assign n240 = ~n238 & ~n239 ;
  assign n241 = n240 ^ n233 ;
  assign n242 = n241 ^ n233 ;
  assign n243 = n235 & ~n242 ;
  assign n244 = n243 ^ n233 ;
  assign n245 = ~x2 & n244 ;
  assign n246 = n245 ^ n233 ;
  assign n247 = n91 & n246 ;
  assign n248 = ~n29 & ~n33 ;
  assign n250 = n218 & n249 ;
  assign n251 = n248 & n250 ;
  assign n252 = ~n48 & n251 ;
  assign n254 = x2 & x12 ;
  assign n255 = ~n253 & ~n254 ;
  assign n256 = ~x2 & x7 ;
  assign n257 = n35 & ~n256 ;
  assign n258 = n255 & n257 ;
  assign n259 = ~n252 & ~n258 ;
  assign n260 = n23 & ~n259 ;
  assign n261 = ~x8 & x12 ;
  assign n262 = n203 & n261 ;
  assign n263 = n91 & n112 ;
  assign n264 = n262 & n263 ;
  assign n266 = n35 & n265 ;
  assign n267 = ~x1 & n84 ;
  assign n268 = n127 & n202 ;
  assign n269 = n267 & n268 ;
  assign n270 = ~n266 & ~n269 ;
  assign n271 = n65 & ~n270 ;
  assign n272 = ~n264 & ~n271 ;
  assign n273 = ~n260 & n272 ;
  assign n274 = n273 ^ x1 ;
  assign n275 = n274 ^ n273 ;
  assign n276 = ~x13 & n91 ;
  assign n277 = x7 & x8 ;
  assign n278 = n24 & ~n277 ;
  assign n279 = ~n202 & ~n230 ;
  assign n280 = n278 & n279 ;
  assign n282 = n256 & ~n281 ;
  assign n283 = x12 & n282 ;
  assign n284 = ~n280 & ~n283 ;
  assign n285 = n276 & ~n284 ;
  assign n286 = x5 & x7 ;
  assign n287 = x3 & n286 ;
  assign n289 = ~n231 & n288 ;
  assign n290 = n287 & n289 ;
  assign n291 = ~n285 & ~n290 ;
  assign n292 = n291 ^ n273 ;
  assign n293 = n292 ^ n273 ;
  assign n294 = ~n275 & ~n293 ;
  assign n295 = n294 ^ n273 ;
  assign n296 = ~x11 & ~n295 ;
  assign n297 = n296 ^ n273 ;
  assign n298 = ~n247 & n297 ;
  assign n299 = ~n229 & n298 ;
  assign n394 = n393 ^ n299 ;
  assign n395 = n394 ^ n299 ;
  assign n396 = ~x1 & x2 ;
  assign n397 = ~x3 & n182 ;
  assign n398 = n84 & n300 ;
  assign n399 = ~n397 & ~n398 ;
  assign n400 = n23 & ~n399 ;
  assign n401 = n396 & n400 ;
  assign n402 = n87 & n124 ;
  assign n403 = n143 & n402 ;
  assign n404 = ~x11 & x12 ;
  assign n405 = x11 & ~x12 ;
  assign n406 = ~x5 & n405 ;
  assign n407 = ~n404 & ~n406 ;
  assign n408 = n403 & ~n407 ;
  assign n409 = n59 & n267 ;
  assign n410 = x1 & x11 ;
  assign n411 = ~x10 & n91 ;
  assign n412 = ~x12 & n206 ;
  assign n413 = ~n411 & ~n412 ;
  assign n414 = n410 & ~n413 ;
  assign n415 = ~n409 & ~n414 ;
  assign n416 = ~n135 & ~n148 ;
  assign n417 = ~x2 & n416 ;
  assign n418 = ~n415 & n417 ;
  assign n419 = ~n408 & ~n418 ;
  assign n420 = ~n401 & n419 ;
  assign n421 = n86 & ~n420 ;
  assign n422 = n421 ^ n299 ;
  assign n423 = n422 ^ n299 ;
  assign n424 = n395 & ~n423 ;
  assign n425 = n424 ^ n299 ;
  assign n426 = ~x9 & n425 ;
  assign n427 = n426 ^ n299 ;
  assign n428 = n196 & n427 ;
  assign n429 = ~n78 & n428 ;
  assign n430 = n19 & ~n429 ;
  assign n431 = x11 & x12 ;
  assign n432 = ~x9 & ~x10 ;
  assign n433 = n431 & n432 ;
  assign n434 = x9 & x10 ;
  assign n435 = n300 & n434 ;
  assign n436 = ~n433 & ~n435 ;
  assign n437 = x0 & x1 ;
  assign n438 = ~x2 & n437 ;
  assign n439 = n190 & n438 ;
  assign n440 = n322 & n439 ;
  assign n441 = n144 ^ x0 ;
  assign n442 = ~x0 & x2 ;
  assign n443 = x8 & n442 ;
  assign n444 = n443 ^ n441 ;
  assign n445 = n444 ^ n144 ;
  assign n446 = n445 ^ n444 ;
  assign n447 = n60 & n322 ;
  assign n448 = n447 ^ n444 ;
  assign n449 = n448 ^ n441 ;
  assign n450 = n446 & ~n449 ;
  assign n451 = n450 ^ n447 ;
  assign n452 = ~x2 & x8 ;
  assign n453 = ~n447 & ~n452 ;
  assign n454 = n453 ^ n441 ;
  assign n455 = ~n451 & ~n454 ;
  assign n456 = n455 ^ n453 ;
  assign n457 = ~n441 & n456 ;
  assign n458 = n457 ^ n450 ;
  assign n459 = n458 ^ x0 ;
  assign n460 = n459 ^ n447 ;
  assign n461 = n112 & ~n460 ;
  assign n462 = n47 & n333 ;
  assign n463 = x7 ^ x0 ;
  assign n464 = n463 ^ x8 ;
  assign n465 = n277 & ~n464 ;
  assign n466 = n465 ^ n464 ;
  assign n467 = n462 & ~n466 ;
  assign n468 = ~n88 & ~n114 ;
  assign n469 = ~x0 & ~n468 ;
  assign n470 = x0 & ~x1 ;
  assign n471 = ~x2 & n470 ;
  assign n472 = n29 & n471 ;
  assign n473 = ~n469 & ~n472 ;
  assign n474 = n307 & ~n473 ;
  assign n475 = x8 ^ x2 ;
  assign n476 = n86 ^ n51 ;
  assign n477 = n51 ^ x8 ;
  assign n478 = n477 ^ n51 ;
  assign n479 = n476 & n478 ;
  assign n480 = n479 ^ n51 ;
  assign n481 = n475 & n480 ;
  assign n482 = x0 & n481 ;
  assign n483 = ~x0 & x8 ;
  assign n484 = n99 ^ x13 ;
  assign n485 = n484 ^ n99 ;
  assign n486 = n101 ^ n99 ;
  assign n487 = ~n485 & n486 ;
  assign n488 = n487 ^ n99 ;
  assign n489 = n483 & n488 ;
  assign n490 = ~n482 & ~n489 ;
  assign n491 = n52 & ~n490 ;
  assign n492 = ~n474 & ~n491 ;
  assign n493 = ~n467 & n492 ;
  assign n494 = x14 & ~n493 ;
  assign n495 = ~n461 & ~n494 ;
  assign n496 = ~n440 & n495 ;
  assign n497 = x3 & ~n496 ;
  assign n498 = ~x3 & x8 ;
  assign n499 = ~x0 & ~x2 ;
  assign n500 = x14 & ~n499 ;
  assign n501 = ~x1 & ~x5 ;
  assign n502 = x13 & ~n501 ;
  assign n503 = ~n500 & ~n502 ;
  assign n504 = n498 & ~n503 ;
  assign n505 = ~n47 & ~n286 ;
  assign n506 = x1 & ~n505 ;
  assign n507 = x14 & ~n51 ;
  assign n508 = n87 & ~n507 ;
  assign n509 = ~n506 & ~n508 ;
  assign n510 = ~x1 & ~x7 ;
  assign n511 = ~n99 & ~n510 ;
  assign n512 = x0 & ~x2 ;
  assign n513 = ~n442 & ~n512 ;
  assign n514 = ~n19 & n513 ;
  assign n515 = n511 & ~n514 ;
  assign n516 = n509 & n515 ;
  assign n517 = n504 & n516 ;
  assign n518 = ~x8 & x14 ;
  assign n519 = ~x7 & n518 ;
  assign n520 = n437 & n519 ;
  assign n521 = n212 & n520 ;
  assign n522 = ~n517 & ~n521 ;
  assign n523 = ~n497 & n522 ;
  assign n524 = ~n436 & ~n523 ;
  assign n525 = ~x8 & ~x9 ;
  assign n526 = ~x13 & ~x14 ;
  assign n527 = x12 & ~n526 ;
  assign n528 = n525 & n527 ;
  assign n529 = x9 & x14 ;
  assign n530 = x8 & n377 ;
  assign n531 = n529 & n530 ;
  assign n532 = ~n528 & ~n531 ;
  assign n533 = ~x1 & x11 ;
  assign n534 = x0 & x10 ;
  assign n535 = n533 & n534 ;
  assign n536 = n198 & n535 ;
  assign n537 = x0 & n343 ;
  assign n538 = n34 & n537 ;
  assign n539 = x5 & ~x10 ;
  assign n540 = ~x0 & ~x1 ;
  assign n541 = x5 & n540 ;
  assign n542 = ~n539 & ~n541 ;
  assign n543 = ~x0 & x1 ;
  assign n544 = ~n470 & ~n543 ;
  assign n545 = n544 ^ n437 ;
  assign n546 = n545 ^ n437 ;
  assign n547 = n437 ^ x10 ;
  assign n548 = n547 ^ n437 ;
  assign n549 = n546 & ~n548 ;
  assign n550 = n549 ^ n437 ;
  assign n551 = x11 & ~n550 ;
  assign n552 = n551 ^ n437 ;
  assign n553 = ~n542 & n552 ;
  assign n554 = ~n538 & ~n553 ;
  assign n555 = n25 & ~n554 ;
  assign n556 = ~x5 & x7 ;
  assign n557 = x1 & ~x3 ;
  assign n558 = n556 & n557 ;
  assign n559 = n537 & n558 ;
  assign n560 = x5 & x11 ;
  assign n561 = ~x10 & n560 ;
  assign n562 = ~x3 & ~x7 ;
  assign n563 = n437 & n562 ;
  assign n564 = n561 & n563 ;
  assign n565 = ~n559 & ~n564 ;
  assign n566 = ~n555 & n565 ;
  assign n567 = x2 & ~n566 ;
  assign n568 = ~n536 & ~n567 ;
  assign n569 = ~n532 & ~n568 ;
  assign n570 = ~x1 & n362 ;
  assign n571 = ~x7 & ~x10 ;
  assign n572 = ~n60 & ~n452 ;
  assign n573 = x0 & ~n572 ;
  assign n574 = ~n443 & ~n573 ;
  assign n575 = n571 & ~n574 ;
  assign n576 = n570 & n575 ;
  assign n577 = x7 & ~x11 ;
  assign n578 = n124 & n438 ;
  assign n579 = n577 & n578 ;
  assign n580 = ~n576 & ~n579 ;
  assign n581 = x5 & n64 ;
  assign n582 = n581 ^ n91 ;
  assign n583 = n582 ^ n91 ;
  assign n584 = n91 ^ x14 ;
  assign n585 = n584 ^ n91 ;
  assign n586 = n583 & n585 ;
  assign n587 = n586 ^ n91 ;
  assign n588 = x9 & n587 ;
  assign n589 = n588 ^ n91 ;
  assign n590 = ~n580 & n589 ;
  assign n591 = x9 & ~x13 ;
  assign n592 = n236 & n591 ;
  assign n593 = n87 & n592 ;
  assign n594 = n277 & n593 ;
  assign n595 = n202 & n434 ;
  assign n596 = n277 & n432 ;
  assign n597 = ~n595 & ~n596 ;
  assign n598 = ~n333 & ~n396 ;
  assign n599 = x12 & ~n598 ;
  assign n600 = ~n597 & n599 ;
  assign n601 = ~x8 & ~x13 ;
  assign n602 = n256 & n434 ;
  assign n603 = n601 & n602 ;
  assign n604 = x7 & ~x9 ;
  assign n605 = ~x7 & x9 ;
  assign n606 = ~n604 & ~n605 ;
  assign n607 = n175 & n606 ;
  assign n608 = ~n603 & ~n607 ;
  assign n609 = n388 & ~n608 ;
  assign n610 = ~n600 & ~n609 ;
  assign n611 = ~n594 & n610 ;
  assign n612 = n97 & ~n611 ;
  assign n613 = ~n590 & ~n612 ;
  assign n614 = x8 & x9 ;
  assign n615 = n84 & n614 ;
  assign n616 = ~n70 & ~n571 ;
  assign n617 = ~n343 & n616 ;
  assign n618 = n615 & n617 ;
  assign n619 = n87 & n618 ;
  assign n620 = n613 & ~n619 ;
  assign n621 = ~n569 & n620 ;
  assign n622 = ~n524 & n621 ;
  assign n623 = ~n300 & ~n431 ;
  assign n624 = ~x0 & x10 ;
  assign n625 = x1 & x3 ;
  assign n626 = x5 & n625 ;
  assign n627 = ~x9 & n51 ;
  assign n628 = n626 & n627 ;
  assign n629 = ~x3 & x9 ;
  assign n630 = n501 & n629 ;
  assign n631 = n86 & n630 ;
  assign n632 = ~n628 & ~n631 ;
  assign n633 = n624 & ~n632 ;
  assign n634 = n51 & n437 ;
  assign n635 = n84 & n634 ;
  assign n636 = n432 & n635 ;
  assign n637 = ~n633 & ~n636 ;
  assign n638 = n623 & ~n637 ;
  assign n639 = x1 & x5 ;
  assign n640 = n51 & n639 ;
  assign n641 = n22 & n80 ;
  assign n642 = x9 & ~x10 ;
  assign n643 = ~n623 & n642 ;
  assign n644 = ~n641 & ~n643 ;
  assign n645 = n640 & ~n644 ;
  assign n646 = n20 & n79 ;
  assign n647 = ~x9 & n192 ;
  assign n648 = ~n646 & ~n647 ;
  assign n649 = x13 ^ x7 ;
  assign n650 = n639 ^ x13 ;
  assign n651 = n649 & ~n650 ;
  assign n652 = n651 ^ x7 ;
  assign n653 = ~n648 & n652 ;
  assign n654 = ~n501 & n653 ;
  assign n655 = ~n645 & ~n654 ;
  assign n656 = n655 ^ x3 ;
  assign n657 = n656 ^ n655 ;
  assign n658 = ~x7 & ~x9 ;
  assign n659 = ~x13 & n658 ;
  assign n660 = n343 & n501 ;
  assign n661 = n659 & n660 ;
  assign n662 = n640 & ~n648 ;
  assign n663 = ~x5 & x9 ;
  assign n664 = ~x12 & n385 ;
  assign n665 = n510 & n664 ;
  assign n666 = n51 & n410 ;
  assign n667 = ~n81 & n666 ;
  assign n668 = ~n665 & ~n667 ;
  assign n669 = n663 & ~n668 ;
  assign n670 = ~n662 & ~n669 ;
  assign n671 = ~n661 & n670 ;
  assign n672 = n671 ^ n655 ;
  assign n673 = ~n657 & n672 ;
  assign n674 = n673 ^ n655 ;
  assign n675 = x0 & ~n674 ;
  assign n676 = ~n638 & ~n675 ;
  assign n677 = x14 & ~n676 ;
  assign n693 = ~x10 & n173 ;
  assign n694 = n287 & n693 ;
  assign n695 = ~x7 & x11 ;
  assign n696 = n59 & n695 ;
  assign n697 = n276 & n696 ;
  assign n698 = ~n694 & ~n697 ;
  assign n678 = ~n51 & n91 ;
  assign n679 = n678 ^ n59 ;
  assign n680 = ~x13 & n571 ;
  assign n681 = n680 ^ n678 ;
  assign n682 = n681 ^ n680 ;
  assign n683 = n682 ^ n679 ;
  assign n684 = n143 ^ n86 ;
  assign n685 = ~n143 & ~n684 ;
  assign n686 = n685 ^ n680 ;
  assign n687 = n686 ^ n143 ;
  assign n688 = ~n683 & n687 ;
  assign n689 = n688 ^ n685 ;
  assign n690 = n689 ^ n143 ;
  assign n691 = n679 & ~n690 ;
  assign n692 = n691 ^ n678 ;
  assign n699 = n698 ^ n692 ;
  assign n700 = n699 ^ n698 ;
  assign n701 = n698 ^ x11 ;
  assign n702 = n701 ^ n698 ;
  assign n703 = n700 & n702 ;
  assign n704 = n703 ^ n698 ;
  assign n705 = ~x1 & ~n704 ;
  assign n706 = n705 ^ n698 ;
  assign n707 = x9 & ~n706 ;
  assign n708 = ~x10 & n404 ;
  assign n709 = ~x9 & n191 ;
  assign n710 = ~n708 & ~n709 ;
  assign n711 = n510 & ~n710 ;
  assign n712 = n431 & n604 ;
  assign n713 = x1 & x10 ;
  assign n714 = n712 & n713 ;
  assign n715 = ~n711 & ~n714 ;
  assign n716 = n276 & ~n715 ;
  assign n717 = ~x1 & n26 ;
  assign n718 = ~n558 & ~n717 ;
  assign n719 = x12 ^ x9 ;
  assign n720 = x12 ^ x10 ;
  assign n721 = n720 ^ x12 ;
  assign n722 = n721 ^ n719 ;
  assign n723 = x13 ^ x11 ;
  assign n724 = ~x11 & n723 ;
  assign n725 = n724 ^ x12 ;
  assign n726 = n725 ^ x11 ;
  assign n727 = ~n722 & ~n726 ;
  assign n728 = n727 ^ n724 ;
  assign n729 = n728 ^ x11 ;
  assign n730 = ~n719 & ~n729 ;
  assign n731 = ~n718 & n730 ;
  assign n732 = ~n716 & ~n731 ;
  assign n733 = ~n707 & n732 ;
  assign n734 = n19 & ~n733 ;
  assign n735 = ~n362 & ~n431 ;
  assign n736 = x1 & x7 ;
  assign n737 = n735 & n736 ;
  assign n738 = ~x12 & n344 ;
  assign n739 = ~x7 & n470 ;
  assign n740 = n738 & n739 ;
  assign n741 = ~n737 & ~n740 ;
  assign n742 = n206 & ~n741 ;
  assign n743 = ~x0 & ~x7 ;
  assign n744 = n28 & n743 ;
  assign n745 = n173 & n744 ;
  assign n747 = ~x5 & ~x11 ;
  assign n746 = n322 & n343 ;
  assign n748 = n747 ^ n746 ;
  assign n749 = x3 & n748 ;
  assign n750 = n749 ^ n747 ;
  assign n751 = n739 & n750 ;
  assign n752 = n97 & ~n137 ;
  assign n753 = ~x0 & ~x3 ;
  assign n754 = x10 & x13 ;
  assign n755 = ~x11 & n754 ;
  assign n756 = n753 & n755 ;
  assign n757 = ~x5 & n756 ;
  assign n758 = ~n752 & ~n757 ;
  assign n759 = n736 & ~n758 ;
  assign n760 = ~n751 & ~n759 ;
  assign n761 = ~n745 & n760 ;
  assign n762 = x12 & ~n761 ;
  assign n763 = x0 & ~x3 ;
  assign n764 = ~x5 & n763 ;
  assign n765 = ~n385 & ~n404 ;
  assign n766 = n510 & n765 ;
  assign n767 = n764 & n766 ;
  assign n768 = ~n762 & ~n767 ;
  assign n769 = ~n742 & n768 ;
  assign n770 = n769 ^ x9 ;
  assign n771 = n770 ^ n769 ;
  assign n772 = n771 ^ n734 ;
  assign n773 = ~x5 & n362 ;
  assign n774 = ~n134 & n165 ;
  assign n775 = n753 & n774 ;
  assign n776 = n773 & n775 ;
  assign n777 = x0 & ~x7 ;
  assign n778 = n267 & n777 ;
  assign n779 = ~n776 & ~n778 ;
  assign n780 = n779 ^ x10 ;
  assign n781 = ~n779 & ~n780 ;
  assign n782 = n781 ^ n769 ;
  assign n783 = n782 ^ n779 ;
  assign n784 = n772 & n783 ;
  assign n785 = n784 ^ n781 ;
  assign n786 = n785 ^ n779 ;
  assign n787 = ~n734 & ~n786 ;
  assign n788 = n787 ^ n734 ;
  assign n789 = ~n677 & ~n788 ;
  assign n790 = ~n572 & ~n789 ;
  assign n791 = ~x8 & ~x14 ;
  assign n792 = ~x9 & n173 ;
  assign n793 = n26 & n792 ;
  assign n794 = x7 & x11 ;
  assign n795 = n91 & n794 ;
  assign n796 = n591 & n795 ;
  assign n797 = ~n793 & ~n796 ;
  assign n798 = n24 & ~n797 ;
  assign n799 = ~x9 & ~x11 ;
  assign n800 = n84 & n799 ;
  assign n801 = x5 & ~x11 ;
  assign n802 = ~n182 & ~n801 ;
  assign n803 = n629 & ~n802 ;
  assign n804 = ~n800 & ~n803 ;
  assign n805 = n29 & ~n804 ;
  assign n806 = n397 & n605 ;
  assign n807 = ~n805 & ~n806 ;
  assign n808 = n166 & ~n807 ;
  assign n809 = ~n798 & ~n808 ;
  assign n810 = ~x10 & ~n809 ;
  assign n811 = ~x13 & n80 ;
  assign n812 = x5 & ~x9 ;
  assign n813 = ~n663 & ~n812 ;
  assign n814 = ~x3 & x11 ;
  assign n815 = ~n813 & n814 ;
  assign n816 = ~n800 & ~n815 ;
  assign n817 = n811 & ~n816 ;
  assign n818 = n256 & n817 ;
  assign n819 = ~n810 & ~n818 ;
  assign n820 = n437 & ~n819 ;
  assign n821 = ~n197 & ~n556 ;
  assign n822 = n69 & n431 ;
  assign n823 = n87 & n300 ;
  assign n824 = ~n822 & ~n823 ;
  assign n825 = n753 & n754 ;
  assign n826 = ~n824 & n825 ;
  assign n827 = n396 & n405 ;
  assign n828 = n129 & n166 ;
  assign n829 = ~n827 & ~n828 ;
  assign n830 = ~x10 & ~x13 ;
  assign n831 = x0 & x3 ;
  assign n832 = n830 & n831 ;
  assign n833 = ~n829 & n832 ;
  assign n834 = ~n826 & ~n833 ;
  assign n835 = x9 & ~n834 ;
  assign n836 = ~n821 & n835 ;
  assign n837 = x3 & ~x11 ;
  assign n838 = n125 & n434 ;
  assign n839 = n616 & n812 ;
  assign n840 = ~n838 & ~n839 ;
  assign n841 = n837 & ~n840 ;
  assign n842 = ~x7 & n91 ;
  assign n843 = x11 & n434 ;
  assign n844 = n842 & n843 ;
  assign n845 = ~n841 & ~n844 ;
  assign n846 = ~x0 & n87 ;
  assign n847 = n377 & n846 ;
  assign n848 = ~n845 & n847 ;
  assign n849 = ~n836 & ~n848 ;
  assign n850 = x12 & n543 ;
  assign n851 = n605 & n773 ;
  assign n852 = ~x3 & n851 ;
  assign n853 = x10 ^ x2 ;
  assign n854 = n853 ^ n852 ;
  assign n855 = ~x13 & n799 ;
  assign n856 = n287 & n855 ;
  assign n857 = n856 ^ x10 ;
  assign n858 = n857 ^ n856 ;
  assign n859 = x3 & ~x9 ;
  assign n860 = ~n33 & ~n577 ;
  assign n861 = ~n802 & ~n860 ;
  assign n862 = n859 & n861 ;
  assign n863 = n862 ^ n856 ;
  assign n864 = ~n858 & n863 ;
  assign n865 = n864 ^ n856 ;
  assign n866 = n865 ^ n852 ;
  assign n867 = ~n854 & n866 ;
  assign n868 = n867 ^ n864 ;
  assign n869 = n868 ^ n856 ;
  assign n870 = n869 ^ n853 ;
  assign n871 = ~n852 & ~n870 ;
  assign n872 = n871 ^ n852 ;
  assign n873 = n872 ^ n853 ;
  assign n874 = n850 & ~n873 ;
  assign n875 = n849 & ~n874 ;
  assign n876 = n648 ^ x13 ;
  assign n877 = n876 ^ n648 ;
  assign n878 = n648 ^ n436 ;
  assign n879 = n877 & n878 ;
  assign n880 = n879 ^ n648 ;
  assign n881 = n649 & ~n880 ;
  assign n882 = ~n513 & n881 ;
  assign n886 = ~n173 & ~n404 ;
  assign n887 = n602 & ~n886 ;
  assign n883 = x7 & ~n22 ;
  assign n884 = x2 & n883 ;
  assign n885 = n237 & n884 ;
  assign n888 = n887 ^ n885 ;
  assign n889 = n888 ^ x0 ;
  assign n898 = n889 ^ n888 ;
  assign n890 = ~x0 & x7 ;
  assign n891 = ~n22 & ~n890 ;
  assign n892 = n891 ^ n889 ;
  assign n893 = n892 ^ n888 ;
  assign n894 = n889 ^ n885 ;
  assign n895 = n894 ^ n891 ;
  assign n896 = n895 ^ n893 ;
  assign n897 = n893 & n896 ;
  assign n899 = n898 ^ n897 ;
  assign n900 = n899 ^ n893 ;
  assign n901 = n166 & n754 ;
  assign n902 = n901 ^ n888 ;
  assign n903 = n897 ^ n893 ;
  assign n904 = n902 & n903 ;
  assign n905 = n904 ^ n888 ;
  assign n906 = n900 & n905 ;
  assign n907 = n906 ^ n888 ;
  assign n908 = n907 ^ n887 ;
  assign n909 = n908 ^ n888 ;
  assign n910 = ~n882 & ~n909 ;
  assign n911 = n84 & ~n910 ;
  assign n920 = x0 & x2 ;
  assign n921 = n344 & n920 ;
  assign n912 = ~x2 & x13 ;
  assign n913 = ~x0 & x11 ;
  assign n914 = x12 & n913 ;
  assign n915 = n912 & n914 ;
  assign n916 = n838 & n915 ;
  assign n922 = n921 ^ n916 ;
  assign n923 = n922 ^ n916 ;
  assign n917 = ~x12 & n642 ;
  assign n918 = n917 ^ n916 ;
  assign n919 = n918 ^ n916 ;
  assign n924 = n923 ^ n919 ;
  assign n925 = n916 ^ n286 ;
  assign n926 = n925 ^ n916 ;
  assign n927 = n926 ^ n923 ;
  assign n928 = n923 & n927 ;
  assign n929 = n928 ^ n923 ;
  assign n930 = n924 & n929 ;
  assign n931 = n930 ^ n928 ;
  assign n932 = n931 ^ n916 ;
  assign n933 = n932 ^ n923 ;
  assign n934 = ~x3 & n933 ;
  assign n935 = n934 ^ n916 ;
  assign n936 = ~n911 & ~n935 ;
  assign n937 = n936 ^ x1 ;
  assign n938 = n937 ^ n936 ;
  assign n939 = n938 ^ n875 ;
  assign n940 = ~x0 & n108 ;
  assign n941 = x12 & x13 ;
  assign n942 = ~x10 & n941 ;
  assign n943 = n940 & n942 ;
  assign n944 = ~x2 & n831 ;
  assign n945 = n811 & n944 ;
  assign n946 = ~n943 & ~n945 ;
  assign n947 = n21 & ~n946 ;
  assign n948 = n947 ^ n821 ;
  assign n949 = n947 & ~n948 ;
  assign n950 = n949 ^ n936 ;
  assign n951 = n950 ^ n947 ;
  assign n952 = n939 & ~n951 ;
  assign n953 = n952 ^ n949 ;
  assign n954 = n953 ^ n947 ;
  assign n955 = n875 & n954 ;
  assign n956 = n955 ^ n875 ;
  assign n957 = ~n820 & n956 ;
  assign n958 = ~n791 & ~n957 ;
  assign n959 = x0 & ~n597 ;
  assign n960 = ~x9 & n281 ;
  assign n961 = n890 & n960 ;
  assign n962 = ~n959 & ~n961 ;
  assign n963 = x2 & ~x11 ;
  assign n964 = ~x12 & n963 ;
  assign n965 = n143 ^ n84 ;
  assign n966 = x1 & ~n965 ;
  assign n967 = n966 ^ n84 ;
  assign n968 = n964 & n967 ;
  assign n969 = ~x2 & ~x11 ;
  assign n970 = ~x1 & n969 ;
  assign n971 = n581 & n970 ;
  assign n972 = n92 & n405 ;
  assign n973 = ~n971 & ~n972 ;
  assign n974 = ~n968 & n973 ;
  assign n975 = ~n526 & ~n974 ;
  assign n976 = n47 & n218 ;
  assign n977 = ~n216 & ~n976 ;
  assign n978 = x11 & x14 ;
  assign n979 = ~x12 & n978 ;
  assign n980 = ~x1 & n979 ;
  assign n981 = ~n977 & n980 ;
  assign n982 = ~n975 & ~n981 ;
  assign n983 = ~n962 & ~n982 ;
  assign n984 = ~n958 & ~n983 ;
  assign n985 = ~n790 & n984 ;
  assign n986 = n622 & n985 ;
  assign n987 = ~n430 & n986 ;
  assign n988 = ~x10 & x14 ;
  assign n989 = ~x9 & n988 ;
  assign n990 = n405 & n989 ;
  assign n991 = n202 & n990 ;
  assign n992 = ~x12 & x14 ;
  assign n993 = n329 & n992 ;
  assign n994 = ~x8 & n993 ;
  assign n995 = ~n606 & n994 ;
  assign n996 = ~n991 & ~n995 ;
  assign n997 = n995 ^ n431 ;
  assign n998 = n190 & n642 ;
  assign n999 = n124 & n604 ;
  assign n1000 = ~n998 & ~n999 ;
  assign n1001 = n1000 ^ n996 ;
  assign n1002 = ~n997 & n1001 ;
  assign n1003 = n1002 ^ n1000 ;
  assign n1004 = n996 & n1003 ;
  assign n1005 = n219 & ~n1004 ;
  assign n1006 = x5 ^ x3 ;
  assign n1007 = x10 & n277 ;
  assign n1008 = n300 & n1007 ;
  assign n1009 = n1008 ^ x5 ;
  assign n1010 = n1009 ^ n1008 ;
  assign n1011 = ~x8 & n152 ;
  assign n1012 = x11 & n1011 ;
  assign n1013 = n79 & n577 ;
  assign n1014 = n230 & n794 ;
  assign n1015 = ~n1008 & ~n1014 ;
  assign n1016 = ~n301 & n1015 ;
  assign n1017 = ~x13 & ~n1016 ;
  assign n1018 = ~n1013 & ~n1017 ;
  assign n1019 = ~n1012 & n1018 ;
  assign n1020 = n1019 ^ n1008 ;
  assign n1021 = ~n1010 & ~n1020 ;
  assign n1022 = n1021 ^ n1008 ;
  assign n1023 = ~n1006 & n1022 ;
  assign n1024 = ~n526 & n1023 ;
  assign n1025 = x11 & ~n29 ;
  assign n1026 = ~x3 & n747 ;
  assign n1027 = ~n97 & ~n1026 ;
  assign n1028 = n261 & ~n1027 ;
  assign n1029 = ~n1025 & n1028 ;
  assign n1030 = x10 & n1029 ;
  assign n1031 = x8 & x12 ;
  assign n1032 = ~x13 & n277 ;
  assign n1033 = ~n1031 & ~n1032 ;
  assign n1034 = ~x7 & ~n405 ;
  assign n1035 = ~n231 & n1034 ;
  assign n1036 = x14 & n84 ;
  assign n1037 = ~n281 & n1036 ;
  assign n1038 = ~n1035 & n1037 ;
  assign n1039 = ~n230 & ~n794 ;
  assign n1040 = ~x12 & ~n1039 ;
  assign n1041 = ~x11 & n59 ;
  assign n1042 = ~x13 & n59 ;
  assign n1043 = ~n1041 & ~n1042 ;
  assign n1044 = ~n1040 & n1043 ;
  assign n1045 = n1038 & n1044 ;
  assign n1046 = n1033 & n1045 ;
  assign n1047 = n136 & n765 ;
  assign n1048 = ~n1046 & ~n1047 ;
  assign n1049 = ~n1030 & n1048 ;
  assign n1050 = ~n1024 & n1049 ;
  assign n1051 = n181 & ~n1050 ;
  assign n1052 = ~x10 & n992 ;
  assign n1053 = n363 & n1052 ;
  assign n1054 = x2 & x10 ;
  assign n1055 = ~n963 & ~n1054 ;
  assign n1056 = ~n1053 & n1055 ;
  assign n1057 = n26 & ~n1056 ;
  assign n1058 = ~x10 & n431 ;
  assign n1059 = x13 & n1058 ;
  assign n1060 = ~x2 & ~n1059 ;
  assign n1061 = n91 & ~n1060 ;
  assign n1062 = x2 & ~n143 ;
  assign n1063 = ~x5 & n128 ;
  assign n1064 = n405 & ~n526 ;
  assign n1065 = n1063 & n1064 ;
  assign n1066 = ~n84 & ~n1065 ;
  assign n1067 = ~n1062 & n1066 ;
  assign n1068 = n1067 ^ x14 ;
  assign n1069 = n1068 ^ n1067 ;
  assign n1070 = ~x13 & n431 ;
  assign n1071 = n1063 & n1070 ;
  assign n1072 = ~n91 & ~n385 ;
  assign n1073 = n24 & n1072 ;
  assign n1074 = n1073 ^ n253 ;
  assign n1075 = n1074 ^ n386 ;
  assign n1076 = n1074 ^ n1073 ;
  assign n1077 = n1076 ^ n1075 ;
  assign n1078 = ~n1075 & ~n1077 ;
  assign n1079 = n1078 ^ n1074 ;
  assign n1080 = n1079 ^ n1075 ;
  assign n1081 = n362 ^ n84 ;
  assign n1082 = n1073 ^ n84 ;
  assign n1083 = ~n1081 & n1082 ;
  assign n1084 = n1083 ^ n1074 ;
  assign n1085 = ~n1080 & n1084 ;
  assign n1086 = n1085 ^ n1074 ;
  assign n1087 = n1086 ^ n1073 ;
  assign n1088 = ~n1071 & ~n1087 ;
  assign n1089 = n1088 ^ n1067 ;
  assign n1090 = n1089 ^ n1067 ;
  assign n1091 = n1069 & ~n1090 ;
  assign n1092 = n1091 ^ n1067 ;
  assign n1093 = ~x10 & ~n1092 ;
  assign n1094 = n1093 ^ n1067 ;
  assign n1095 = ~n1061 & n1094 ;
  assign n1096 = x7 & ~n1095 ;
  assign n1097 = ~n1057 & ~n1096 ;
  assign n1098 = n614 & ~n1097 ;
  assign n1099 = ~x10 & n105 ;
  assign n1100 = n287 & n1099 ;
  assign n1101 = x7 & ~x8 ;
  assign n1102 = ~n152 & ~n1101 ;
  assign n1103 = ~n366 & n1102 ;
  assign n1104 = ~x13 & x14 ;
  assign n1105 = ~x8 & n1104 ;
  assign n1106 = ~x10 & ~n1105 ;
  assign n1107 = n1026 & ~n1106 ;
  assign n1108 = n1103 & n1107 ;
  assign n1109 = ~n1100 & ~n1108 ;
  assign n1110 = n166 & ~n1109 ;
  assign n1111 = ~x1 & ~n1110 ;
  assign n1112 = x2 & ~x9 ;
  assign n1113 = n300 & n1104 ;
  assign n1114 = n411 & n1113 ;
  assign n1115 = ~n206 & ~n1114 ;
  assign n1116 = n277 & ~n1115 ;
  assign n1117 = n84 & n190 ;
  assign n1118 = n236 & ~n1104 ;
  assign n1119 = n334 & ~n1118 ;
  assign n1120 = ~n343 & n1119 ;
  assign n1121 = ~n1117 & ~n1120 ;
  assign n1122 = n411 & n765 ;
  assign n1123 = ~n124 & ~n1122 ;
  assign n1124 = n84 & ~n735 ;
  assign n1125 = ~n1123 & ~n1124 ;
  assign n1126 = x7 & n1125 ;
  assign n1127 = n1121 & ~n1126 ;
  assign n1128 = ~n1116 & n1127 ;
  assign n1129 = n1112 & ~n1128 ;
  assign n1130 = n1111 & ~n1129 ;
  assign n1131 = ~n1098 & n1130 ;
  assign n1132 = ~x8 & x9 ;
  assign n1133 = x7 ^ x2 ;
  assign n1134 = ~x2 & x11 ;
  assign n1135 = x12 & n1134 ;
  assign n1136 = n206 & n1135 ;
  assign n1137 = n91 & n345 ;
  assign n1138 = n84 & n306 ;
  assign n1139 = ~n1137 & ~n1138 ;
  assign n1140 = x12 & ~n1139 ;
  assign n1141 = ~n231 & ~n431 ;
  assign n1142 = n91 & ~n1141 ;
  assign n1143 = n84 & n362 ;
  assign n1144 = x12 & n1143 ;
  assign n1145 = ~n1142 & ~n1144 ;
  assign n1146 = n988 & ~n1145 ;
  assign n1147 = x10 & x14 ;
  assign n1148 = n623 ^ n276 ;
  assign n1149 = n1148 ^ n276 ;
  assign n1150 = x3 & n47 ;
  assign n1151 = n1150 ^ n276 ;
  assign n1152 = n1149 & n1151 ;
  assign n1153 = n1152 ^ n276 ;
  assign n1154 = n1147 & n1153 ;
  assign n1155 = ~n1146 & ~n1154 ;
  assign n1156 = ~n1140 & n1155 ;
  assign n1157 = n256 & ~n1156 ;
  assign n1158 = ~n1136 & ~n1157 ;
  assign n1159 = n1158 ^ n1133 ;
  assign n1160 = n142 & n191 ;
  assign n1161 = ~n539 & n802 ;
  assign n1162 = ~x3 & n1161 ;
  assign n1163 = ~n1160 & ~n1162 ;
  assign n1164 = n941 & ~n1163 ;
  assign n1165 = n59 & n142 ;
  assign n1166 = ~n411 & ~n1165 ;
  assign n1167 = n344 & ~n1166 ;
  assign n1171 = n581 ^ n54 ;
  assign n1172 = n1171 ^ n581 ;
  assign n1168 = ~n173 & ~n801 ;
  assign n1169 = n1168 ^ n581 ;
  assign n1170 = n1169 ^ n581 ;
  assign n1173 = n1172 ^ n1170 ;
  assign n1174 = n581 ^ x12 ;
  assign n1175 = n1174 ^ n581 ;
  assign n1176 = n1175 ^ n1172 ;
  assign n1177 = n1172 & n1176 ;
  assign n1178 = n1177 ^ n1172 ;
  assign n1179 = n1173 & n1178 ;
  assign n1180 = n1179 ^ n1177 ;
  assign n1181 = n1180 ^ n581 ;
  assign n1182 = n1181 ^ n1172 ;
  assign n1183 = x10 & n1182 ;
  assign n1184 = n1183 ^ n581 ;
  assign n1185 = ~n1167 & ~n1184 ;
  assign n1186 = x14 & ~n1185 ;
  assign n1187 = ~n1164 & ~n1186 ;
  assign n1188 = n1187 ^ x2 ;
  assign n1189 = n1188 ^ n1187 ;
  assign n1190 = ~n231 & ~n992 ;
  assign n1191 = n91 & ~n1190 ;
  assign n1192 = x12 & x14 ;
  assign n1193 = ~n127 & ~n1192 ;
  assign n1194 = ~n143 & ~n1193 ;
  assign n1195 = ~n1191 & ~n1194 ;
  assign n1196 = n343 & ~n1195 ;
  assign n1197 = x13 & x14 ;
  assign n1198 = x13 & ~n1197 ;
  assign n1199 = ~n143 & ~n1198 ;
  assign n1200 = ~n1036 & ~n1199 ;
  assign n1201 = n192 & ~n1200 ;
  assign n1202 = ~n1196 & ~n1201 ;
  assign n1203 = ~n91 & ~n1036 ;
  assign n1204 = n1058 & ~n1203 ;
  assign n1205 = n84 & n127 ;
  assign n1206 = ~n91 & ~n1205 ;
  assign n1207 = ~x5 & x10 ;
  assign n1208 = ~x3 & n1207 ;
  assign n1209 = ~n329 & ~n1208 ;
  assign n1210 = ~n1206 & ~n1209 ;
  assign n1211 = ~n1204 & ~n1210 ;
  assign n1212 = n1202 & n1211 ;
  assign n1213 = n1212 ^ n1187 ;
  assign n1214 = n1189 & n1213 ;
  assign n1215 = n1214 ^ n1187 ;
  assign n1216 = n1215 ^ n1133 ;
  assign n1217 = ~n1159 & n1216 ;
  assign n1218 = n1217 ^ n1214 ;
  assign n1219 = n1218 ^ n1187 ;
  assign n1220 = n1219 ^ n1158 ;
  assign n1221 = ~n1133 & ~n1220 ;
  assign n1222 = n1221 ^ n1133 ;
  assign n1223 = n1222 ^ n1158 ;
  assign n1224 = n1132 & n1223 ;
  assign n1225 = n1131 & ~n1224 ;
  assign n1226 = ~n1051 & n1225 ;
  assign n1227 = x2 & n1104 ;
  assign n1228 = ~x13 & ~n1227 ;
  assign n1229 = n1026 & ~n1228 ;
  assign n1230 = x14 ^ x13 ;
  assign n1231 = n1230 ^ n84 ;
  assign n1233 = ~n963 & ~n1134 ;
  assign n1232 = x2 & x11 ;
  assign n1234 = n1233 ^ n1232 ;
  assign n1235 = x14 & ~n1234 ;
  assign n1236 = n1235 ^ n1232 ;
  assign n1237 = ~n1231 & n1236 ;
  assign n1238 = n1237 ^ n1235 ;
  assign n1239 = n1238 ^ n1232 ;
  assign n1240 = n1239 ^ x14 ;
  assign n1241 = n84 & n1240 ;
  assign n1242 = ~n1229 & ~n1241 ;
  assign n1243 = n236 & ~n1242 ;
  assign n1244 = x8 & ~n397 ;
  assign n1245 = ~n281 & ~n1244 ;
  assign n1246 = ~n1243 & ~n1245 ;
  assign n1247 = ~x5 & ~x12 ;
  assign n1248 = ~n1228 & n1247 ;
  assign n1249 = ~x3 & n1248 ;
  assign n1250 = x10 & ~n397 ;
  assign n1251 = ~n1249 & n1250 ;
  assign n1252 = n300 & ~n526 ;
  assign n1253 = ~n738 & ~n1252 ;
  assign n1254 = n219 & ~n1253 ;
  assign n1255 = ~x2 & x14 ;
  assign n1256 = ~x2 & n127 ;
  assign n1257 = ~n1255 & ~n1256 ;
  assign n1258 = n84 & ~n1257 ;
  assign n1259 = ~n623 & n1258 ;
  assign n1260 = ~n1254 & ~n1259 ;
  assign n1261 = n1251 & n1260 ;
  assign n1262 = n1104 ^ n941 ;
  assign n1263 = n1262 ^ x11 ;
  assign n1271 = n1263 ^ n1262 ;
  assign n1264 = x2 & n623 ;
  assign n1265 = n1264 ^ n1263 ;
  assign n1266 = n1265 ^ n1262 ;
  assign n1267 = n1263 ^ n941 ;
  assign n1268 = n1267 ^ n1264 ;
  assign n1269 = n1268 ^ n1266 ;
  assign n1270 = n1266 & ~n1269 ;
  assign n1272 = n1271 ^ n1270 ;
  assign n1273 = n1272 ^ n1266 ;
  assign n1274 = n1262 ^ x2 ;
  assign n1275 = n1270 ^ n1266 ;
  assign n1276 = n1274 & n1275 ;
  assign n1277 = n1276 ^ n1262 ;
  assign n1278 = ~n1273 & n1277 ;
  assign n1279 = n1278 ^ n1262 ;
  assign n1280 = n1279 ^ n1104 ;
  assign n1281 = n1280 ^ n1262 ;
  assign n1282 = n91 & n1281 ;
  assign n1283 = n581 & n1255 ;
  assign n1284 = n230 & ~n1283 ;
  assign n1285 = ~n1282 & n1284 ;
  assign n1286 = ~n1261 & ~n1285 ;
  assign n1287 = n219 & n431 ;
  assign n1288 = ~n1286 & ~n1287 ;
  assign n1289 = ~n1246 & ~n1288 ;
  assign n1290 = n143 ^ x2 ;
  assign n1291 = n1290 ^ n143 ;
  assign n1292 = n1291 ^ n281 ;
  assign n1293 = ~n84 & ~n91 ;
  assign n1294 = n1293 ^ n837 ;
  assign n1295 = ~n1293 & n1294 ;
  assign n1296 = n1295 ^ n143 ;
  assign n1297 = n1296 ^ n1293 ;
  assign n1298 = ~n1292 & n1297 ;
  assign n1299 = n1298 ^ n1295 ;
  assign n1300 = n1299 ^ n1293 ;
  assign n1301 = n281 & ~n1300 ;
  assign n1302 = n1301 ^ n281 ;
  assign n1303 = ~n1289 & ~n1302 ;
  assign n1304 = ~x9 & ~n1303 ;
  assign n1305 = ~x2 & n1104 ;
  assign n1306 = n300 & n1305 ;
  assign n1307 = ~x8 & ~n404 ;
  assign n1308 = ~n174 & ~n1307 ;
  assign n1309 = ~n1306 & ~n1308 ;
  assign n1310 = n1208 & ~n1309 ;
  assign n1311 = ~n1304 & ~n1310 ;
  assign n1312 = ~x7 & ~n1311 ;
  assign n1313 = ~n24 & n411 ;
  assign n1314 = ~x12 & ~x14 ;
  assign n1315 = ~n377 & ~n1314 ;
  assign n1316 = n83 & n1315 ;
  assign n1317 = n1313 & n1316 ;
  assign n1318 = ~x14 & n144 ;
  assign n1319 = ~n591 & n978 ;
  assign n1320 = x5 & ~n799 ;
  assign n1321 = ~n1198 & ~n1320 ;
  assign n1322 = ~n1319 & ~n1321 ;
  assign n1323 = ~x8 & n66 ;
  assign n1324 = ~x5 & n22 ;
  assign n1325 = n1323 & ~n1324 ;
  assign n1326 = ~n1322 & n1325 ;
  assign n1327 = ~n1318 & n1326 ;
  assign n1328 = ~x14 & n362 ;
  assign n1329 = x12 & n65 ;
  assign n1330 = ~n105 & n1329 ;
  assign n1331 = ~n1328 & n1330 ;
  assign n1332 = ~x14 & ~n127 ;
  assign n1333 = ~n765 & ~n1332 ;
  assign n1334 = ~x2 & n230 ;
  assign n1335 = n1333 & n1334 ;
  assign n1336 = ~x13 & n992 ;
  assign n1337 = n1134 & n1336 ;
  assign n1338 = ~n404 & ~n1337 ;
  assign n1339 = n23 & ~n1338 ;
  assign n1340 = ~n1335 & ~n1339 ;
  assign n1341 = ~n1331 & n1340 ;
  assign n1342 = n663 & ~n1341 ;
  assign n1343 = ~n237 & ~n378 ;
  assign n1344 = ~n1058 & n1343 ;
  assign n1345 = n1255 & ~n1344 ;
  assign n1346 = x11 & n65 ;
  assign n1347 = ~n377 & n1346 ;
  assign n1348 = ~x8 & ~n1347 ;
  assign n1349 = ~n708 & n1348 ;
  assign n1350 = ~n1345 & n1349 ;
  assign n1351 = ~x5 & ~x9 ;
  assign n1352 = ~n23 & n1351 ;
  assign n1353 = ~n1350 & n1352 ;
  assign n1354 = ~x2 & ~n22 ;
  assign n1355 = x5 & ~x8 ;
  assign n1356 = x10 & n1355 ;
  assign n1357 = n1354 & n1356 ;
  assign n1358 = ~n1193 & n1357 ;
  assign n1359 = ~n1353 & ~n1358 ;
  assign n1360 = ~n1342 & n1359 ;
  assign n1361 = n1360 ^ x3 ;
  assign n1362 = n1361 ^ n1360 ;
  assign n1363 = n1362 ^ n1327 ;
  assign n1364 = x5 & x12 ;
  assign n1365 = ~x8 & n1364 ;
  assign n1366 = n799 & n1365 ;
  assign n1367 = ~n137 & n1366 ;
  assign n1368 = n168 & n231 ;
  assign n1369 = ~n802 & n1368 ;
  assign n1370 = n404 & n591 ;
  assign n1371 = n230 & n1370 ;
  assign n1372 = ~n960 & ~n1371 ;
  assign n1373 = n1372 ^ x5 ;
  assign n1374 = n1373 ^ n1372 ;
  assign n1375 = n1374 ^ n1369 ;
  assign n1376 = n405 & n1197 ;
  assign n1377 = n642 & ~n1376 ;
  assign n1378 = n1377 ^ x8 ;
  assign n1379 = ~n1377 & ~n1378 ;
  assign n1380 = n1379 ^ n1372 ;
  assign n1381 = n1380 ^ n1377 ;
  assign n1382 = ~n1375 & n1381 ;
  assign n1383 = n1382 ^ n1379 ;
  assign n1384 = n1383 ^ n1377 ;
  assign n1385 = ~n1369 & ~n1384 ;
  assign n1386 = n1385 ^ n1369 ;
  assign n1387 = ~n1367 & ~n1386 ;
  assign n1388 = n1387 ^ x2 ;
  assign n1389 = x2 & ~n1388 ;
  assign n1390 = n1389 ^ n1360 ;
  assign n1391 = n1390 ^ x2 ;
  assign n1392 = ~n1363 & ~n1391 ;
  assign n1393 = n1392 ^ n1389 ;
  assign n1394 = n1393 ^ x2 ;
  assign n1395 = ~n1327 & n1394 ;
  assign n1396 = n1395 ^ n1327 ;
  assign n1397 = n1396 ^ x7 ;
  assign n1398 = ~x13 & ~n648 ;
  assign n1399 = n1355 & n1398 ;
  assign n1400 = x5 & n82 ;
  assign n1401 = x10 & n1400 ;
  assign n1402 = ~n993 & ~n1058 ;
  assign n1403 = n1402 ^ x8 ;
  assign n1404 = n1403 ^ n1402 ;
  assign n1405 = n1404 ^ n1351 ;
  assign n1406 = ~n173 & n992 ;
  assign n1407 = n1406 ^ x10 ;
  assign n1408 = ~n1406 & n1407 ;
  assign n1409 = n1408 ^ n1402 ;
  assign n1410 = n1409 ^ n1406 ;
  assign n1411 = ~n1405 & ~n1410 ;
  assign n1412 = n1411 ^ n1408 ;
  assign n1413 = n1412 ^ n1406 ;
  assign n1414 = n1351 & ~n1413 ;
  assign n1415 = n1414 ^ n1351 ;
  assign n1416 = ~n1401 & ~n1415 ;
  assign n1417 = n23 & ~n1252 ;
  assign n1418 = ~n993 & n1307 ;
  assign n1419 = n1070 ^ x10 ;
  assign n1420 = n1419 ^ n1070 ;
  assign n1421 = n1253 ^ n1070 ;
  assign n1422 = n1420 & ~n1421 ;
  assign n1423 = n1422 ^ n1070 ;
  assign n1424 = n1418 & ~n1423 ;
  assign n1425 = n663 & ~n1424 ;
  assign n1426 = ~n1417 & n1425 ;
  assign n1427 = n1416 & ~n1426 ;
  assign n1428 = ~n1399 & n1427 ;
  assign n1429 = n108 & ~n1428 ;
  assign n1430 = n1429 ^ n736 ;
  assign n1431 = ~n1397 & n1430 ;
  assign n1432 = n1431 ^ n1429 ;
  assign n1433 = n736 & n1432 ;
  assign n1434 = n1433 ^ x1 ;
  assign n1435 = ~n1317 & n1434 ;
  assign n1436 = n84 & n1336 ;
  assign n1437 = ~n91 & ~n1436 ;
  assign n1438 = n329 & ~n1437 ;
  assign n1439 = x14 & n343 ;
  assign n1440 = ~n143 & n231 ;
  assign n1441 = ~n581 & ~n1440 ;
  assign n1442 = n1439 & ~n1441 ;
  assign n1443 = n1202 & ~n1442 ;
  assign n1444 = ~n1438 & n1443 ;
  assign n1445 = n452 & ~n1444 ;
  assign n1446 = n334 & n708 ;
  assign n1447 = ~n1445 & ~n1446 ;
  assign n1448 = ~n199 & ~n1031 ;
  assign n1449 = n84 & ~n1448 ;
  assign n1450 = n334 & n1336 ;
  assign n1451 = ~n1205 & ~n1450 ;
  assign n1452 = ~n1449 & n1451 ;
  assign n1453 = n329 & ~n1452 ;
  assign n1454 = x3 & n314 ;
  assign n1455 = ~n312 & ~n431 ;
  assign n1456 = n315 & ~n1455 ;
  assign n1457 = ~n1454 & ~n1456 ;
  assign n1458 = x10 & ~n1457 ;
  assign n1459 = ~x8 & n343 ;
  assign n1460 = ~x12 & ~n1197 ;
  assign n1461 = n84 & ~n1460 ;
  assign n1462 = ~n526 & ~n1314 ;
  assign n1463 = n91 & n1462 ;
  assign n1464 = ~n1461 & ~n1463 ;
  assign n1465 = n1459 & ~n1464 ;
  assign n1466 = ~n1458 & ~n1465 ;
  assign n1467 = ~x13 & n1293 ;
  assign n1468 = ~n1036 & ~n1467 ;
  assign n1469 = ~x12 & n1099 ;
  assign n1470 = ~n1468 & n1469 ;
  assign n1471 = ~n308 & ~n1470 ;
  assign n1472 = n1466 & n1471 ;
  assign n1473 = ~n1453 & n1472 ;
  assign n1474 = n1473 ^ x2 ;
  assign n1475 = n1474 ^ n1473 ;
  assign n1476 = n1475 ^ n1447 ;
  assign n1477 = n623 ^ n431 ;
  assign n1478 = x10 & n1477 ;
  assign n1479 = n1478 ^ n431 ;
  assign n1480 = n1150 & n1479 ;
  assign n1481 = n81 & n276 ;
  assign n1482 = ~n305 & n1481 ;
  assign n1483 = ~n1480 & ~n1482 ;
  assign n1484 = x14 & ~n1483 ;
  assign n1485 = ~n84 & ~n362 ;
  assign n1486 = n59 & ~n1485 ;
  assign n1487 = ~n1072 & n1486 ;
  assign n1488 = ~n1484 & ~n1487 ;
  assign n1489 = n1488 ^ x8 ;
  assign n1490 = ~x8 & n1489 ;
  assign n1491 = n1490 ^ n1473 ;
  assign n1492 = n1491 ^ x8 ;
  assign n1493 = ~n1476 & n1492 ;
  assign n1494 = n1493 ^ n1490 ;
  assign n1495 = n1494 ^ x8 ;
  assign n1496 = n1447 & ~n1495 ;
  assign n1497 = n1496 ^ n1447 ;
  assign n1498 = n605 & ~n1497 ;
  assign n1499 = n1435 & ~n1498 ;
  assign n1500 = ~n1312 & n1499 ;
  assign n1501 = ~n1226 & ~n1500 ;
  assign n1502 = ~n1005 & ~n1501 ;
  assign n1503 = n1502 ^ x0 ;
  assign n1504 = n1503 ^ n1502 ;
  assign n1505 = ~x8 & n577 ;
  assign n1506 = n28 & n1505 ;
  assign n1507 = x1 & ~x10 ;
  assign n1508 = n84 & n1507 ;
  assign n1509 = n695 & n1508 ;
  assign n1510 = ~n1506 & ~n1509 ;
  assign n1511 = n254 & ~n1510 ;
  assign n1512 = x9 & n1511 ;
  assign n1513 = n51 & ~n1132 ;
  assign n1514 = ~x3 & n1513 ;
  assign n1515 = n1324 & n1514 ;
  assign n1516 = n86 & n615 ;
  assign n1517 = x11 & n1516 ;
  assign n1518 = ~n1515 & ~n1517 ;
  assign n1519 = n396 & ~n1518 ;
  assign n1520 = ~x3 & n190 ;
  assign n1521 = n34 & n1520 ;
  assign n1522 = n792 & n1521 ;
  assign n1523 = ~n1519 & ~n1522 ;
  assign n1524 = ~n81 & ~n1523 ;
  assign n1525 = n28 & n605 ;
  assign n1526 = ~n231 & n1525 ;
  assign n1527 = ~x3 & x12 ;
  assign n1528 = n137 & n1527 ;
  assign n1529 = n736 & n1528 ;
  assign n1530 = ~n813 & n1529 ;
  assign n1531 = ~n51 & ~n591 ;
  assign n1532 = ~x9 & n53 ;
  assign n1533 = x1 & ~n821 ;
  assign n1534 = ~n1532 & ~n1533 ;
  assign n1535 = x7 & x9 ;
  assign n1536 = ~x10 & ~n1535 ;
  assign n1537 = n64 & n1536 ;
  assign n1538 = ~n1534 & n1537 ;
  assign n1539 = ~n1531 & n1538 ;
  assign n1540 = ~n1530 & ~n1539 ;
  assign n1541 = ~n1526 & n1540 ;
  assign n1542 = n963 & ~n1541 ;
  assign n1543 = n48 & n1026 ;
  assign n1546 = n1543 ^ x9 ;
  assign n1555 = n1546 ^ n1543 ;
  assign n1544 = n97 & n112 ;
  assign n1545 = n1544 ^ n1543 ;
  assign n1547 = n1546 ^ n1545 ;
  assign n1548 = n1547 ^ n1546 ;
  assign n1549 = n1548 ^ n1543 ;
  assign n1550 = ~x9 & ~x13 ;
  assign n1551 = n1550 ^ n1547 ;
  assign n1552 = n1551 ^ n1547 ;
  assign n1553 = n1552 ^ n1549 ;
  assign n1554 = n1549 & ~n1553 ;
  assign n1556 = n1555 ^ n1554 ;
  assign n1557 = n1556 ^ n1549 ;
  assign n1558 = n1543 ^ x2 ;
  assign n1559 = n1554 ^ n1549 ;
  assign n1560 = n1558 & n1559 ;
  assign n1561 = n1560 ^ n1543 ;
  assign n1562 = n1557 & ~n1561 ;
  assign n1563 = n1562 ^ n1543 ;
  assign n1564 = n1563 ^ x9 ;
  assign n1565 = n1564 ^ n1543 ;
  assign n1566 = n79 & n1565 ;
  assign n1567 = ~x10 & n604 ;
  assign n1568 = n626 & n1567 ;
  assign n1569 = ~n1525 & ~n1568 ;
  assign n1570 = n1232 & ~n1569 ;
  assign n1571 = ~n1566 & ~n1570 ;
  assign n1572 = ~n1542 & n1571 ;
  assign n1573 = x8 & ~n1572 ;
  assign n1574 = ~n1524 & ~n1573 ;
  assign n1575 = ~n1512 & n1574 ;
  assign n1576 = ~x1 & x12 ;
  assign n1577 = x3 & ~x8 ;
  assign n1578 = ~n51 & ~n505 ;
  assign n1579 = x9 & x11 ;
  assign n1580 = ~x9 & ~n344 ;
  assign n1581 = ~n1579 & ~n1580 ;
  assign n1582 = n1578 & n1581 ;
  assign n1583 = ~n851 & ~n1582 ;
  assign n1584 = n1577 & ~n1583 ;
  assign n1585 = n525 & n1026 ;
  assign n1586 = x13 & n1579 ;
  assign n1587 = n202 & n1586 ;
  assign n1588 = n141 & n1587 ;
  assign n1589 = ~x3 & n556 ;
  assign n1590 = ~n346 & ~n601 ;
  assign n1591 = ~n21 & n1590 ;
  assign n1592 = n1589 & n1591 ;
  assign n1593 = ~n1588 & ~n1592 ;
  assign n1594 = ~n1585 & n1593 ;
  assign n1595 = ~n1584 & n1594 ;
  assign n1596 = n1576 & ~n1595 ;
  assign n1597 = ~x8 & n127 ;
  assign n1598 = n801 & n859 ;
  assign n1599 = n1597 & n1598 ;
  assign n1600 = x9 & ~n300 ;
  assign n1601 = n91 & ~n1600 ;
  assign n1602 = ~n143 & ~n404 ;
  assign n1603 = ~n82 & ~n308 ;
  assign n1604 = ~n1602 & ~n1603 ;
  assign n1605 = ~n1601 & n1604 ;
  assign n1606 = ~n1599 & ~n1605 ;
  assign n1607 = n736 & ~n1606 ;
  assign n1608 = ~x1 & ~x9 ;
  assign n1609 = ~n795 & ~n1117 ;
  assign n1610 = n1608 & ~n1609 ;
  assign n1611 = ~n1607 & ~n1610 ;
  assign n1612 = ~n1596 & n1611 ;
  assign n1613 = n615 ^ x7 ;
  assign n1614 = n1613 ^ n615 ;
  assign n1615 = n1614 ^ n1612 ;
  assign n1616 = ~x11 & n614 ;
  assign n1617 = x9 ^ x5 ;
  assign n1618 = n1617 ^ x9 ;
  assign n1619 = n22 ^ x9 ;
  assign n1620 = n1618 & ~n1619 ;
  assign n1621 = n1620 ^ x9 ;
  assign n1622 = n98 & n1621 ;
  assign n1623 = ~n1616 & ~n1622 ;
  assign n1624 = ~n747 & n1527 ;
  assign n1625 = ~n1623 & n1624 ;
  assign n1626 = ~x9 & n362 ;
  assign n1627 = ~x5 & x12 ;
  assign n1628 = n1626 & n1627 ;
  assign n1629 = ~n55 & ~n1550 ;
  assign n1630 = n404 & ~n1351 ;
  assign n1631 = n1629 & n1630 ;
  assign n1632 = x5 & x9 ;
  assign n1633 = n765 & n1632 ;
  assign n1634 = ~n1631 & ~n1633 ;
  assign n1635 = ~n1628 & n1634 ;
  assign n1636 = n1635 ^ x8 ;
  assign n1637 = n1636 ^ n1635 ;
  assign n1638 = n404 & n663 ;
  assign n1639 = n738 & n812 ;
  assign n1640 = ~n1638 & ~n1639 ;
  assign n1641 = n1640 ^ n1635 ;
  assign n1642 = n1637 & n1641 ;
  assign n1643 = n1642 ^ n1635 ;
  assign n1644 = x3 & ~n1643 ;
  assign n1645 = ~n1625 & ~n1644 ;
  assign n1646 = n1645 ^ x1 ;
  assign n1647 = ~n1645 & ~n1646 ;
  assign n1648 = n1647 ^ n615 ;
  assign n1649 = n1648 ^ n1645 ;
  assign n1650 = ~n1615 & ~n1649 ;
  assign n1651 = n1650 ^ n1647 ;
  assign n1652 = n1651 ^ n1645 ;
  assign n1653 = n1612 & ~n1652 ;
  assign n1654 = n1653 ^ n1612 ;
  assign n1655 = x2 & ~n1654 ;
  assign n1656 = n84 & ~n606 ;
  assign n1657 = n533 & n1656 ;
  assign n1658 = n86 & n626 ;
  assign n1659 = ~x1 & n51 ;
  assign n1660 = ~n143 & n1659 ;
  assign n1661 = ~n1658 & ~n1660 ;
  assign n1662 = n1354 & ~n1661 ;
  assign n1663 = ~n1543 & ~n1662 ;
  assign n1664 = ~n1657 & n1663 ;
  assign n1665 = x8 & ~n1664 ;
  assign n1666 = ~x7 & ~n912 ;
  assign n1667 = ~x8 & n1579 ;
  assign n1668 = n267 & n1667 ;
  assign n1669 = ~n1666 & n1668 ;
  assign n1670 = x1 & ~n190 ;
  assign n1671 = ~n86 & n1670 ;
  assign n1672 = ~n85 & ~n1671 ;
  assign n1673 = n91 & n799 ;
  assign n1674 = ~n1672 & n1673 ;
  assign n1675 = ~n1669 & ~n1674 ;
  assign n1676 = ~n1665 & n1675 ;
  assign n1677 = x12 & ~n1676 ;
  assign n1678 = ~n1655 & ~n1677 ;
  assign n1679 = x10 & ~n1678 ;
  assign n1680 = n189 & n1535 ;
  assign n1681 = ~x9 & n48 ;
  assign n1682 = n91 & n1681 ;
  assign n1683 = ~n1680 & ~n1682 ;
  assign n1684 = x11 & n281 ;
  assign n1685 = ~n1683 & n1684 ;
  assign n1686 = ~n1679 & ~n1685 ;
  assign n1687 = n1575 & n1686 ;
  assign n1688 = n1687 ^ n1502 ;
  assign n1689 = ~n1504 & n1688 ;
  assign n1690 = n1689 ^ n1502 ;
  assign n1691 = n987 & n1690 ;
  assign n1692 = n18 & ~n1691 ;
  assign n1693 = ~n23 & ~n124 ;
  assign n1694 = ~n129 & ~n533 ;
  assign n1711 = ~x4 & x5 ;
  assign n1712 = ~x6 & x12 ;
  assign n1713 = n1711 & n1712 ;
  assign n1714 = n218 & n1535 ;
  assign n1715 = n1713 & n1714 ;
  assign n1716 = ~x3 & x6 ;
  assign n1717 = ~x4 & n1716 ;
  assign n1718 = x4 & ~x5 ;
  assign n1719 = ~x6 & n1718 ;
  assign n1720 = ~n1717 & ~n1719 ;
  assign n1721 = n1535 & ~n1720 ;
  assign n1722 = x4 & ~x6 ;
  assign n1723 = n1535 & n1722 ;
  assign n1724 = ~x4 & n658 ;
  assign n1725 = x6 & n1724 ;
  assign n1726 = ~n1723 & ~n1725 ;
  assign n1727 = n141 & ~n1726 ;
  assign n1728 = x4 & ~x9 ;
  assign n1729 = x6 & x7 ;
  assign n1730 = ~n1728 & ~n1729 ;
  assign n1731 = ~x4 & x9 ;
  assign n1732 = ~x6 & ~x7 ;
  assign n1733 = ~n1731 & ~n1732 ;
  assign n1734 = n142 & ~n1733 ;
  assign n1735 = ~n1730 & n1734 ;
  assign n1736 = ~n1727 & ~n1735 ;
  assign n1737 = ~x13 & ~n1736 ;
  assign n1738 = ~n1721 & ~n1737 ;
  assign n1739 = n253 & ~n1738 ;
  assign n1740 = ~n1715 & ~n1739 ;
  assign n1695 = ~x4 & n254 ;
  assign n1696 = x6 & ~x9 ;
  assign n1697 = n197 & n1696 ;
  assign n1698 = ~x5 & n1535 ;
  assign n1699 = ~x6 & x13 ;
  assign n1700 = n1698 & n1699 ;
  assign n1701 = ~n1697 & ~n1700 ;
  assign n1702 = n1695 & ~n1701 ;
  assign n1703 = ~n322 & ~n1535 ;
  assign n1704 = ~n658 & ~n1535 ;
  assign n1705 = ~x2 & x4 ;
  assign n1706 = x6 & ~x12 ;
  assign n1707 = n1705 & n1706 ;
  assign n1708 = ~n1704 & n1707 ;
  assign n1709 = ~n1703 & n1708 ;
  assign n1710 = ~n1702 & ~n1709 ;
  assign n1741 = n1740 ^ n1710 ;
  assign n1742 = n1741 ^ n1740 ;
  assign n1743 = n1740 ^ x3 ;
  assign n1744 = n1743 ^ n1740 ;
  assign n1745 = ~n1742 & ~n1744 ;
  assign n1746 = n1745 ^ n1740 ;
  assign n1747 = ~x0 & ~n1746 ;
  assign n1748 = n1747 ^ n1740 ;
  assign n1749 = x14 & ~n1748 ;
  assign n1750 = n25 & n1728 ;
  assign n1751 = ~x2 & n1706 ;
  assign n1752 = n323 & n1751 ;
  assign n1753 = x2 & ~x6 ;
  assign n1754 = ~x5 & n1753 ;
  assign n1755 = x12 & n1754 ;
  assign n1756 = ~n1752 & ~n1755 ;
  assign n1757 = n19 & ~n1756 ;
  assign n1758 = n1750 & n1757 ;
  assign n1788 = ~x4 & n84 ;
  assign n1789 = n920 & n1788 ;
  assign n1759 = ~x0 & x5 ;
  assign n1760 = ~x3 & n1722 ;
  assign n1761 = n254 & n1760 ;
  assign n1762 = n1759 & n1761 ;
  assign n1763 = n1695 ^ n143 ;
  assign n1764 = ~x0 & x3 ;
  assign n1765 = ~x5 & x6 ;
  assign n1766 = n1764 & n1765 ;
  assign n1767 = n1766 ^ n1763 ;
  assign n1768 = n1767 ^ n1695 ;
  assign n1769 = n1768 ^ n1767 ;
  assign n1770 = ~x12 & n512 ;
  assign n1771 = n17 & n1770 ;
  assign n1772 = n1771 ^ n1767 ;
  assign n1773 = n1772 ^ n1763 ;
  assign n1774 = n1769 & ~n1773 ;
  assign n1775 = n1774 ^ n1771 ;
  assign n1776 = x0 & ~x6 ;
  assign n1777 = ~n1771 & ~n1776 ;
  assign n1778 = n1777 ^ n1763 ;
  assign n1779 = ~n1775 & n1778 ;
  assign n1780 = n1779 ^ n1777 ;
  assign n1781 = n1763 & n1780 ;
  assign n1782 = n1781 ^ n1774 ;
  assign n1783 = n1782 ^ n143 ;
  assign n1784 = n1783 ^ n1771 ;
  assign n1785 = ~n1762 & ~n1784 ;
  assign n1790 = n1789 ^ n1785 ;
  assign n1791 = n1790 ^ n1785 ;
  assign n1786 = n1785 ^ n1712 ;
  assign n1787 = n1786 ^ n1785 ;
  assign n1792 = n1791 ^ n1787 ;
  assign n1793 = n1785 ^ n658 ;
  assign n1794 = n1793 ^ n1785 ;
  assign n1795 = n1794 ^ n1791 ;
  assign n1796 = n1791 & ~n1795 ;
  assign n1797 = n1796 ^ n1791 ;
  assign n1798 = n1792 & n1797 ;
  assign n1799 = n1798 ^ n1796 ;
  assign n1800 = n1799 ^ n1785 ;
  assign n1801 = n1800 ^ n1791 ;
  assign n1802 = ~n1535 & ~n1801 ;
  assign n1803 = n1802 ^ n1785 ;
  assign n1804 = ~n1198 & ~n1803 ;
  assign n1805 = ~x2 & x5 ;
  assign n1806 = n1706 & n1805 ;
  assign n1807 = n1750 & n1806 ;
  assign n1808 = ~x4 & ~x5 ;
  assign n1809 = n1535 & n1808 ;
  assign n1810 = n1527 & n1753 ;
  assign n1811 = n1809 & n1810 ;
  assign n1812 = ~n1807 & ~n1811 ;
  assign n1813 = n1812 ^ x0 ;
  assign n1814 = n1813 ^ n1812 ;
  assign n1815 = n1814 ^ n526 ;
  assign n1816 = n197 & n1728 ;
  assign n1817 = x3 & x6 ;
  assign n1818 = n255 & n1817 ;
  assign n1819 = n1818 ^ n1816 ;
  assign n1820 = n1816 & n1819 ;
  assign n1821 = n1820 ^ n1812 ;
  assign n1822 = n1821 ^ n1816 ;
  assign n1823 = n1815 & ~n1822 ;
  assign n1824 = n1823 ^ n1820 ;
  assign n1825 = n1824 ^ n1816 ;
  assign n1826 = ~n526 & n1825 ;
  assign n1827 = ~n1804 & ~n1826 ;
  assign n1828 = ~n1758 & n1827 ;
  assign n1829 = ~n1749 & n1828 ;
  assign n1830 = ~n1694 & ~n1829 ;
  assign n1831 = x0 & x5 ;
  assign n1832 = x12 & n1535 ;
  assign n1833 = x6 & n27 ;
  assign n1834 = n1832 & n1833 ;
  assign n1835 = ~x3 & x4 ;
  assign n1836 = ~x7 & n1608 ;
  assign n1837 = n127 & n1535 ;
  assign n1838 = n1837 ^ x1 ;
  assign n1839 = n1838 ^ n1837 ;
  assign n1840 = ~n377 & n658 ;
  assign n1841 = n1840 ^ n1837 ;
  assign n1842 = n1839 & n1841 ;
  assign n1843 = n1842 ^ n1837 ;
  assign n1844 = ~x6 & n1843 ;
  assign n1845 = ~n1836 & ~n1844 ;
  assign n1846 = n1835 & ~n1845 ;
  assign n1847 = x6 & ~x13 ;
  assign n1848 = n134 & n1847 ;
  assign n1849 = n1750 & n1848 ;
  assign n1850 = ~n1846 & ~n1849 ;
  assign n1851 = ~n1834 & n1850 ;
  assign n1852 = n1134 & ~n1851 ;
  assign n1853 = ~x9 & x12 ;
  assign n1854 = n48 & n1853 ;
  assign n1855 = n1699 ^ x4 ;
  assign n1856 = n1855 ^ n1699 ;
  assign n1857 = n1699 ^ x2 ;
  assign n1858 = n1856 & n1857 ;
  assign n1859 = n1858 ^ n1699 ;
  assign n1860 = ~n1753 & n1859 ;
  assign n1861 = n1854 & ~n1860 ;
  assign n1862 = n17 & n69 ;
  assign n1863 = n377 & ~n606 ;
  assign n1864 = n1862 & n1863 ;
  assign n1865 = x2 & ~x4 ;
  assign n1866 = n1535 & n1865 ;
  assign n1867 = ~x6 & n127 ;
  assign n1868 = n1866 & n1867 ;
  assign n1869 = n1753 ^ n1724 ;
  assign n1870 = n1753 ^ n166 ;
  assign n1871 = n1870 ^ n166 ;
  assign n1872 = x4 & x7 ;
  assign n1873 = n170 & n1872 ;
  assign n1874 = n1873 ^ n166 ;
  assign n1875 = n1871 & ~n1874 ;
  assign n1876 = n1875 ^ n166 ;
  assign n1877 = n1869 & ~n1876 ;
  assign n1878 = n1877 ^ n1724 ;
  assign n1879 = ~n1868 & ~n1878 ;
  assign n1880 = ~x1 & ~n1879 ;
  assign n1881 = ~n1864 & ~n1880 ;
  assign n1882 = ~n1861 & n1881 ;
  assign n1883 = n837 & ~n1882 ;
  assign n1884 = n396 & n1535 ;
  assign n1885 = ~x9 & n99 ;
  assign n1886 = x9 & ~x12 ;
  assign n1887 = n100 & n1886 ;
  assign n1888 = ~n1885 & ~n1887 ;
  assign n1889 = x1 & ~n1888 ;
  assign n1890 = x13 & ~n99 ;
  assign n1891 = x9 & x13 ;
  assign n1892 = ~n1890 & ~n1891 ;
  assign n1893 = n1889 & n1892 ;
  assign n1894 = ~n1884 & ~n1893 ;
  assign n1895 = n1760 & ~n1894 ;
  assign n1896 = ~x1 & x6 ;
  assign n1897 = n1866 & n1896 ;
  assign n1898 = x2 & x4 ;
  assign n1899 = ~x6 & n1898 ;
  assign n1900 = n1535 & n1899 ;
  assign n1901 = ~x2 & n1724 ;
  assign n1902 = ~n1900 & ~n1901 ;
  assign n1903 = n557 & ~n1902 ;
  assign n1904 = ~n1897 & ~n1903 ;
  assign n1905 = x12 & ~n1904 ;
  assign n1906 = n377 & n1885 ;
  assign n1907 = n27 & n1906 ;
  assign n1908 = x4 & n1907 ;
  assign n1909 = ~n1905 & ~n1908 ;
  assign n1910 = ~n1895 & n1909 ;
  assign n1911 = n1910 ^ x11 ;
  assign n1912 = n1911 ^ n1910 ;
  assign n1913 = n1912 ^ n1883 ;
  assign n1914 = x3 & ~x6 ;
  assign n1915 = ~x1 & ~n377 ;
  assign n1916 = ~n127 & ~n1915 ;
  assign n1917 = n1914 & ~n1916 ;
  assign n1918 = ~n27 & ~n1917 ;
  assign n1919 = n1724 & ~n1918 ;
  assign n1920 = n1576 & n1723 ;
  assign n1921 = ~n1919 & ~n1920 ;
  assign n1922 = n1921 ^ x2 ;
  assign n1923 = ~n1921 & ~n1922 ;
  assign n1924 = n1923 ^ n1910 ;
  assign n1925 = n1924 ^ n1921 ;
  assign n1926 = ~n1913 & n1925 ;
  assign n1927 = n1926 ^ n1923 ;
  assign n1928 = n1927 ^ n1921 ;
  assign n1929 = ~n1883 & ~n1928 ;
  assign n1930 = n1929 ^ n1883 ;
  assign n1931 = ~n1852 & ~n1930 ;
  assign n1932 = n1831 & ~n1931 ;
  assign n1933 = x4 & n442 ;
  assign n1934 = n1896 & n1933 ;
  assign n1935 = ~x7 & n404 ;
  assign n1936 = x3 & n1935 ;
  assign n1937 = n1934 & n1936 ;
  assign n1938 = ~x1 & n1729 ;
  assign n1939 = x3 & x4 ;
  assign n1940 = n499 & n1939 ;
  assign n1941 = n1940 ^ x12 ;
  assign n1942 = n1940 ^ n385 ;
  assign n1943 = n1942 ^ n385 ;
  assign n1944 = ~x0 & x13 ;
  assign n1945 = ~n1232 & ~n1944 ;
  assign n1946 = ~x3 & ~x4 ;
  assign n1947 = ~n969 & n1946 ;
  assign n1948 = ~n1945 & n1947 ;
  assign n1949 = n1948 ^ n385 ;
  assign n1950 = ~n1943 & n1949 ;
  assign n1951 = n1950 ^ n385 ;
  assign n1952 = n1941 & ~n1951 ;
  assign n1953 = n1952 ^ x12 ;
  assign n1954 = n1938 & n1953 ;
  assign n1955 = x2 & x6 ;
  assign n1956 = ~n1817 & ~n1955 ;
  assign n1957 = ~n431 & n1956 ;
  assign n1958 = n736 & ~n1957 ;
  assign n1959 = ~x12 & n362 ;
  assign n1960 = x3 & ~x4 ;
  assign n1961 = x6 & ~n1960 ;
  assign n1962 = ~n1959 & n1961 ;
  assign n1963 = n1962 ^ x2 ;
  assign n1964 = n1963 ^ n1962 ;
  assign n1965 = ~n17 & ~n1817 ;
  assign n1966 = x3 & x13 ;
  assign n1967 = ~n1939 & ~n1966 ;
  assign n1968 = ~n664 & n1967 ;
  assign n1969 = n1965 & n1968 ;
  assign n1970 = ~n763 & n1969 ;
  assign n1971 = n1970 ^ n1962 ;
  assign n1972 = n1964 & n1971 ;
  assign n1973 = n1972 ^ n1962 ;
  assign n1974 = n1958 & n1973 ;
  assign n1975 = ~n1954 & ~n1974 ;
  assign n1976 = ~n1937 & n1975 ;
  assign n1977 = n1632 & ~n1976 ;
  assign n1978 = n1232 & n1832 ;
  assign n1979 = ~n1760 & ~n1960 ;
  assign n1980 = n1978 & ~n1979 ;
  assign n1981 = ~x6 & n64 ;
  assign n1982 = ~x7 & n799 ;
  assign n1983 = n1579 & n1872 ;
  assign n1984 = ~n1982 & ~n1983 ;
  assign n1985 = n1981 & ~n1984 ;
  assign n1986 = n512 & n1985 ;
  assign n1987 = ~n1980 & ~n1986 ;
  assign n1988 = n792 & n1732 ;
  assign n1989 = ~n1535 & ~n1699 ;
  assign n1990 = ~n658 & n1232 ;
  assign n1991 = ~n1989 & n1990 ;
  assign n1992 = ~n1988 & ~n1991 ;
  assign n1993 = n1527 & ~n1992 ;
  assign n1994 = x2 & ~x13 ;
  assign n1995 = x3 & x9 ;
  assign n1996 = n1706 & n1995 ;
  assign n1997 = n1994 & n1996 ;
  assign n1998 = n577 & n1997 ;
  assign n1999 = ~n1993 & ~n1998 ;
  assign n2000 = ~x4 & ~n1999 ;
  assign n2001 = ~x2 & x6 ;
  assign n2002 = n658 & n1960 ;
  assign n2003 = x9 & n1872 ;
  assign n2004 = ~n2002 & ~n2003 ;
  assign n2005 = n2004 ^ n362 ;
  assign n2006 = n2005 ^ n2004 ;
  assign n2007 = n1535 & n1835 ;
  assign n2008 = ~n2002 & ~n2007 ;
  assign n2009 = n2008 ^ n2004 ;
  assign n2010 = n2009 ^ n2004 ;
  assign n2011 = ~n2006 & ~n2010 ;
  assign n2012 = n2011 ^ n2004 ;
  assign n2013 = ~n431 & ~n2012 ;
  assign n2014 = n2013 ^ n2004 ;
  assign n2015 = n2001 & ~n2014 ;
  assign n2016 = ~n2000 & ~n2015 ;
  assign n2017 = n2016 ^ x0 ;
  assign n2018 = n2017 ^ n2016 ;
  assign n2019 = n1714 ^ x3 ;
  assign n2020 = n2019 ^ n1714 ;
  assign n2021 = n1714 ^ n658 ;
  assign n2022 = n2021 ^ n1714 ;
  assign n2023 = ~n2020 & n2022 ;
  assign n2024 = n2023 ^ n1714 ;
  assign n2025 = x6 & n2024 ;
  assign n2026 = n2025 ^ n1714 ;
  assign n2027 = n765 & n2026 ;
  assign n2028 = n108 & n1535 ;
  assign n2029 = n1706 & n2028 ;
  assign n2030 = n173 & n2029 ;
  assign n2031 = ~n2027 & ~n2030 ;
  assign n2032 = x4 & ~n2031 ;
  assign n2033 = ~x4 & ~x11 ;
  assign n2034 = ~n1722 & ~n2033 ;
  assign n2035 = ~x6 & ~x13 ;
  assign n2036 = n2028 & ~n2035 ;
  assign n2037 = n2034 & n2036 ;
  assign n2038 = x12 & n2037 ;
  assign n2039 = x11 & n256 ;
  assign n2040 = x4 & x9 ;
  assign n2041 = n2039 & n2040 ;
  assign n2042 = n1982 & n2001 ;
  assign n2043 = ~x11 & n1535 ;
  assign n2044 = n1899 & n2043 ;
  assign n2045 = ~n2042 & ~n2044 ;
  assign n2046 = ~n2041 & n2045 ;
  assign n2047 = n64 & ~n2046 ;
  assign n2048 = ~n2038 & ~n2047 ;
  assign n2049 = ~n2032 & n2048 ;
  assign n2050 = n2049 ^ n2016 ;
  assign n2051 = ~n2018 & n2050 ;
  assign n2052 = n2051 ^ n2016 ;
  assign n2053 = n1987 & n2052 ;
  assign n2054 = n34 & ~n2053 ;
  assign n2055 = n846 & n1935 ;
  assign n2056 = ~x2 & n540 ;
  assign n2057 = x12 & ~n2056 ;
  assign n2058 = n385 & ~n2057 ;
  assign n2059 = x1 & n1944 ;
  assign n2060 = x7 & ~n2059 ;
  assign n2061 = ~n1959 & n2060 ;
  assign n2062 = ~x12 & n499 ;
  assign n2063 = ~n540 & ~n969 ;
  assign n2064 = ~n134 & ~n2063 ;
  assign n2065 = ~n2062 & n2064 ;
  assign n2066 = n2061 & n2065 ;
  assign n2067 = ~n2058 & n2066 ;
  assign n2068 = ~n2055 & ~n2067 ;
  assign n2069 = x9 & ~n2068 ;
  assign n2070 = n438 & n738 ;
  assign n2071 = ~n824 & n1944 ;
  assign n2072 = ~n2070 & ~n2071 ;
  assign n2073 = ~n606 & ~n2072 ;
  assign n2074 = n543 & n658 ;
  assign n2075 = n362 ^ x12 ;
  assign n2076 = x12 ^ x2 ;
  assign n2077 = n2075 & n2076 ;
  assign n2078 = n2077 ^ x12 ;
  assign n2079 = n2074 & n2078 ;
  assign n2080 = ~n2073 & ~n2079 ;
  assign n2081 = ~n2069 & n2080 ;
  assign n2082 = n17 & ~n2081 ;
  assign n2083 = x0 & ~x4 ;
  assign n2084 = ~x6 & n2083 ;
  assign n2085 = ~x9 & n695 ;
  assign n2086 = n941 & n2085 ;
  assign n2087 = n2084 & n2086 ;
  assign n2088 = n87 & n2087 ;
  assign n2089 = ~n2082 & ~n2088 ;
  assign n2090 = n1293 & ~n2089 ;
  assign n2091 = ~n2054 & ~n2090 ;
  assign n2092 = ~n1977 & n2091 ;
  assign n2093 = ~n1932 & n2092 ;
  assign n2094 = ~n1830 & n2093 ;
  assign n2095 = ~x3 & ~x6 ;
  assign n2096 = ~n1817 & ~n2095 ;
  assign n2097 = ~n824 & n1809 ;
  assign n2098 = n253 & n658 ;
  assign n2099 = x1 & x4 ;
  assign n2100 = n560 & n2099 ;
  assign n2101 = n2098 & n2100 ;
  assign n2102 = ~n2097 & ~n2101 ;
  assign n2103 = x0 & ~n2102 ;
  assign n2104 = ~x4 & n410 ;
  assign n2105 = n499 & n1535 ;
  assign n2106 = n2104 & n2105 ;
  assign n2107 = x12 & n2106 ;
  assign n2108 = ~n2103 & ~n2107 ;
  assign n2109 = ~n2096 & ~n2108 ;
  assign n2110 = n913 & n1715 ;
  assign n2111 = n2110 ^ n2109 ;
  assign n2112 = n437 & n1753 ;
  assign n2113 = x4 & ~x12 ;
  assign n2114 = n629 & n2113 ;
  assign n2115 = n2112 & n2114 ;
  assign n2116 = n286 & n2115 ;
  assign n2117 = n2056 & n2113 ;
  assign n2118 = n1696 & n2117 ;
  assign n2119 = n1731 & n1753 ;
  assign n2120 = x0 & x12 ;
  assign n2121 = n2120 ^ x1 ;
  assign n2122 = n2119 & n2121 ;
  assign n2123 = ~n2118 & ~n2122 ;
  assign n2124 = n287 & ~n2123 ;
  assign n2125 = ~n2116 & ~n2124 ;
  assign n2126 = n2125 ^ x11 ;
  assign n2127 = n2126 ^ n2125 ;
  assign n2128 = ~x5 & ~x6 ;
  assign n2129 = n1535 & n2128 ;
  assign n2130 = ~x0 & n166 ;
  assign n2131 = n2129 & n2130 ;
  assign n2132 = n1960 & n2131 ;
  assign n2133 = n69 & n1535 ;
  assign n2134 = n1722 & n1764 ;
  assign n2135 = ~x12 & n2134 ;
  assign n2136 = ~x0 & ~x4 ;
  assign n2137 = x4 ^ x3 ;
  assign n2138 = n1776 & n2137 ;
  assign n2139 = ~n2136 & ~n2138 ;
  assign n2140 = ~n1706 & ~n1712 ;
  assign n2141 = x5 & ~n2140 ;
  assign n2142 = ~n2139 & n2141 ;
  assign n2143 = ~n2135 & ~n2142 ;
  assign n2144 = n2133 & ~n2143 ;
  assign n2145 = n108 & n719 ;
  assign n2147 = x5 & x6 ;
  assign n2148 = ~n2128 & ~n2147 ;
  assign n2149 = x4 & n2148 ;
  assign n2150 = ~n16 & ~n2149 ;
  assign n2146 = ~x6 & n1808 ;
  assign n2151 = n2150 ^ n2146 ;
  assign n2152 = n2150 ^ x12 ;
  assign n2153 = n2152 ^ n2150 ;
  assign n2154 = n2153 ^ n2145 ;
  assign n2155 = ~n2151 & n2154 ;
  assign n2156 = n2155 ^ n2146 ;
  assign n2157 = n2145 & n2156 ;
  assign n2158 = n2157 ^ x9 ;
  assign n2159 = x6 & n166 ;
  assign n2160 = n1835 & n2159 ;
  assign n2161 = n2160 ^ x5 ;
  assign n2162 = n2161 ^ n2160 ;
  assign n2163 = n1705 & ~n2140 ;
  assign n2164 = n2163 ^ n2160 ;
  assign n2165 = n2162 & n2164 ;
  assign n2166 = n2165 ^ n2160 ;
  assign n2167 = n2166 ^ n2157 ;
  assign n2168 = ~n2158 & ~n2167 ;
  assign n2169 = n2168 ^ n2165 ;
  assign n2170 = n2169 ^ n2160 ;
  assign n2171 = n2170 ^ x9 ;
  assign n2172 = ~n2157 & n2171 ;
  assign n2173 = n2172 ^ n2157 ;
  assign n2174 = n2173 ^ n2157 ;
  assign n2175 = n890 & ~n2174 ;
  assign n2177 = x0 & ~n1718 ;
  assign n2176 = n890 & n1718 ;
  assign n2178 = n2177 ^ n2176 ;
  assign n2179 = n2178 ^ x9 ;
  assign n2186 = n2179 ^ n2178 ;
  assign n2180 = n2179 ^ n2003 ;
  assign n2181 = n2180 ^ n2178 ;
  assign n2182 = n2179 ^ n2176 ;
  assign n2183 = n2182 ^ n2003 ;
  assign n2184 = n2183 ^ n2181 ;
  assign n2185 = ~n2181 & ~n2184 ;
  assign n2187 = n2186 ^ n2185 ;
  assign n2188 = n2187 ^ n2181 ;
  assign n2189 = n2178 ^ n125 ;
  assign n2190 = n2185 ^ n2181 ;
  assign n2191 = ~n2189 & ~n2190 ;
  assign n2192 = n2191 ^ n2178 ;
  assign n2193 = ~n2188 & n2192 ;
  assign n2194 = n2193 ^ n2178 ;
  assign n2195 = n2194 ^ n2177 ;
  assign n2196 = n2195 ^ n2178 ;
  assign n2197 = n1751 & n2196 ;
  assign n2198 = ~x0 & n1865 ;
  assign n2199 = n1706 & n2198 ;
  assign n2200 = n1698 & n2199 ;
  assign n2201 = n606 & n920 ;
  assign n2202 = n1713 & n2201 ;
  assign n2203 = ~n2200 & ~n2202 ;
  assign n2204 = ~n2197 & n2203 ;
  assign n2205 = n2204 ^ n17 ;
  assign n2206 = n2205 ^ n2204 ;
  assign n2207 = n1698 & n1770 ;
  assign n2208 = n2207 ^ n2204 ;
  assign n2209 = n2208 ^ n2204 ;
  assign n2210 = n2206 & n2209 ;
  assign n2211 = n2210 ^ n2204 ;
  assign n2212 = ~x3 & ~n2211 ;
  assign n2213 = n2212 ^ n2204 ;
  assign n2214 = ~n2175 & n2213 ;
  assign n2215 = x1 & ~n2214 ;
  assign n2216 = ~n2144 & ~n2215 ;
  assign n2217 = ~n2132 & n2216 ;
  assign n2218 = n2217 ^ n2125 ;
  assign n2219 = n2127 & n2218 ;
  assign n2220 = n2219 ^ n2125 ;
  assign n2221 = n2220 ^ n2109 ;
  assign n2222 = n2111 & ~n2221 ;
  assign n2223 = n2222 ^ n2219 ;
  assign n2224 = n2223 ^ n2125 ;
  assign n2225 = n2224 ^ n2110 ;
  assign n2226 = ~n2109 & ~n2225 ;
  assign n2227 = n2226 ^ n2109 ;
  assign n2228 = x13 & n2227 ;
  assign n2240 = ~x1 & ~n513 ;
  assign n2241 = n1817 & n2033 ;
  assign n2242 = x4 & x5 ;
  assign n2243 = ~x6 & n2242 ;
  assign n2244 = ~x11 & n2243 ;
  assign n2245 = ~n2241 & ~n2244 ;
  assign n2246 = n2240 & ~n2245 ;
  assign n2247 = x0 & ~x5 ;
  assign n2248 = ~x6 & n1946 ;
  assign n2249 = n2247 & n2248 ;
  assign n2231 = x5 & ~x6 ;
  assign n2232 = n1835 & n2231 ;
  assign n2233 = ~x4 & x6 ;
  assign n2234 = n142 & n2233 ;
  assign n2235 = ~n2232 & ~n2234 ;
  assign n2250 = n437 & ~n2235 ;
  assign n2251 = n540 & ~n1720 ;
  assign n2252 = ~n2250 & ~n2251 ;
  assign n2253 = ~n2249 & n2252 ;
  assign n2254 = n1232 & ~n2253 ;
  assign n2255 = ~n2246 & ~n2254 ;
  assign n2229 = n1946 & n2128 ;
  assign n2230 = n437 & n2229 ;
  assign n2236 = x0 & ~x11 ;
  assign n2237 = n544 & ~n2236 ;
  assign n2238 = ~n2235 & n2237 ;
  assign n2239 = ~n2230 & ~n2238 ;
  assign n2256 = n2255 ^ n2239 ;
  assign n2257 = n2256 ^ n2255 ;
  assign n2258 = n2255 ^ x2 ;
  assign n2259 = n2258 ^ n2255 ;
  assign n2260 = ~n2257 & ~n2259 ;
  assign n2261 = n2260 ^ n2255 ;
  assign n2262 = x12 & ~n2261 ;
  assign n2263 = n2262 ^ n2255 ;
  assign n2264 = n1535 & ~n2263 ;
  assign n2265 = x12 & n1579 ;
  assign n2266 = n108 & n543 ;
  assign n2267 = n2265 & n2266 ;
  assign n2268 = n2146 & n2267 ;
  assign n2269 = ~x1 & ~x11 ;
  assign n2270 = ~x0 & n2269 ;
  assign n2271 = n1707 & n2270 ;
  assign n2272 = n2271 ^ n829 ;
  assign n2273 = n2272 ^ n2271 ;
  assign n2274 = n2271 ^ n2084 ;
  assign n2275 = n2274 ^ n2271 ;
  assign n2276 = ~n2273 & n2275 ;
  assign n2277 = n2276 ^ n2271 ;
  assign n2278 = ~x9 & n2277 ;
  assign n2279 = n2278 ^ n2271 ;
  assign n2280 = n84 & n2279 ;
  assign n2281 = ~n2268 & ~n2280 ;
  assign n2282 = ~n248 & ~n2281 ;
  assign n2283 = n16 & n87 ;
  assign n2284 = ~n1862 & ~n2283 ;
  assign n2285 = x0 & ~n2284 ;
  assign n2286 = ~n1934 & ~n2285 ;
  assign n2287 = n837 & ~n2286 ;
  assign n2288 = ~x0 & n17 ;
  assign n2289 = n1134 & n2288 ;
  assign n2290 = x1 & n2289 ;
  assign n2291 = ~n2287 & ~n2290 ;
  assign n2292 = n249 & ~n2291 ;
  assign n2293 = n410 & n2095 ;
  assign n2294 = n1817 & n2269 ;
  assign n2295 = ~n2293 & ~n2294 ;
  assign n2296 = n2130 & n2242 ;
  assign n2297 = ~n2295 & n2296 ;
  assign n2298 = ~x4 & x12 ;
  assign n2299 = ~x0 & n218 ;
  assign n2300 = n533 & n2299 ;
  assign n2301 = n218 & n543 ;
  assign n2302 = ~n2300 & ~n2301 ;
  assign n2303 = n2231 & ~n2302 ;
  assign n2304 = x11 & n1776 ;
  assign n2305 = ~n92 & ~n189 ;
  assign n2306 = n2304 & ~n2305 ;
  assign n2307 = x6 & x11 ;
  assign n2308 = ~x0 & n142 ;
  assign n2309 = n2307 & n2308 ;
  assign n2310 = n333 & n2309 ;
  assign n2311 = ~n2306 & ~n2310 ;
  assign n2312 = ~n2303 & n2311 ;
  assign n2313 = n2298 & ~n2312 ;
  assign n2314 = ~n2297 & ~n2313 ;
  assign n2315 = ~n2292 & n2314 ;
  assign n2316 = n658 & ~n2315 ;
  assign n2317 = ~n220 & ~n2043 ;
  assign n2318 = ~n1886 & ~n2317 ;
  assign n2319 = n333 & n2318 ;
  assign n2320 = n964 & n1681 ;
  assign n2321 = n533 & ~n1888 ;
  assign n2322 = ~n2320 & ~n2321 ;
  assign n2323 = ~n2319 & n2322 ;
  assign n2324 = n1835 & ~n2323 ;
  assign n2325 = n396 & n2318 ;
  assign n2326 = n969 & n1854 ;
  assign n2327 = ~n2325 & ~n2326 ;
  assign n2328 = n1960 & ~n2327 ;
  assign n2329 = ~n2324 & ~n2328 ;
  assign n2330 = n1759 & ~n2329 ;
  assign n2331 = n1946 & n2247 ;
  assign n2332 = n300 & n1884 ;
  assign n2333 = n87 & n658 ;
  assign n2334 = n388 & n1232 ;
  assign n2335 = ~n2333 & ~n2334 ;
  assign n2336 = ~n623 & ~n1704 ;
  assign n2337 = ~n2335 & ~n2336 ;
  assign n2338 = ~n598 & n2085 ;
  assign n2339 = ~n2337 & ~n2338 ;
  assign n2340 = ~n2332 & n2339 ;
  assign n2341 = n2331 & ~n2340 ;
  assign n2342 = n605 & n827 ;
  assign n2343 = n20 & n112 ;
  assign n2344 = n21 & n48 ;
  assign n2345 = ~n2343 & ~n2344 ;
  assign n2346 = ~n303 & ~n2345 ;
  assign n2347 = ~x1 & x9 ;
  assign n2348 = n99 & ~n410 ;
  assign n2349 = ~n172 & n2348 ;
  assign n2350 = ~n2347 & n2349 ;
  assign n2351 = ~n2346 & ~n2350 ;
  assign n2352 = ~n2342 & n2351 ;
  assign n2353 = x0 & n1788 ;
  assign n2354 = ~n2352 & n2353 ;
  assign n2355 = ~x2 & n1939 ;
  assign n2356 = n850 & n2355 ;
  assign n2357 = n747 & n2356 ;
  assign n2358 = n658 & n2357 ;
  assign n2359 = ~n2354 & ~n2358 ;
  assign n2360 = ~n2341 & n2359 ;
  assign n2361 = ~n2330 & n2360 ;
  assign n2362 = n2035 & ~n2361 ;
  assign n2363 = ~n2316 & ~n2362 ;
  assign n2364 = n134 & n256 ;
  assign n2365 = n20 & n2364 ;
  assign n2366 = ~n2346 & ~n2365 ;
  assign n2367 = x13 & ~n2366 ;
  assign n2368 = ~x2 & n533 ;
  assign n2369 = n1837 & n2368 ;
  assign n2370 = ~x0 & ~n2369 ;
  assign n2371 = n127 & n396 ;
  assign n2372 = x1 & ~n377 ;
  assign n2373 = n255 & n2372 ;
  assign n2374 = ~n2371 & ~n2373 ;
  assign n2375 = n2043 & ~n2374 ;
  assign n2376 = n510 & n1550 ;
  assign n2377 = n1264 & n2376 ;
  assign n2378 = ~n2375 & ~n2377 ;
  assign n2379 = n2370 & n2378 ;
  assign n2380 = ~n2367 & n2379 ;
  assign n2381 = n1946 & n2147 ;
  assign n2382 = n1939 & n2128 ;
  assign n2383 = ~n2381 & ~n2382 ;
  assign n2384 = n377 & n1535 ;
  assign n2385 = n127 & n658 ;
  assign n2386 = ~n2384 & ~n2385 ;
  assign n2387 = n2386 ^ x12 ;
  assign n2388 = n2387 ^ n2386 ;
  assign n2389 = n2386 ^ n659 ;
  assign n2390 = n2389 ^ n2386 ;
  assign n2391 = ~n2388 & n2390 ;
  assign n2392 = n2391 ^ n2386 ;
  assign n2393 = x2 & ~n2392 ;
  assign n2394 = n2393 ^ n2386 ;
  assign n2395 = n1694 & ~n2394 ;
  assign n2396 = n134 & ~n1233 ;
  assign n2397 = ~n822 & ~n2396 ;
  assign n2398 = n658 & ~n2397 ;
  assign n2399 = n385 & n1535 ;
  assign n2400 = n304 & n2399 ;
  assign n2401 = x0 & ~n2400 ;
  assign n2402 = ~n2398 & n2401 ;
  assign n2403 = ~n2395 & n2402 ;
  assign n2404 = ~n2383 & ~n2403 ;
  assign n2405 = ~n2380 & n2404 ;
  assign n2406 = ~n658 & n1134 ;
  assign n2407 = ~n963 & ~n2406 ;
  assign n2408 = ~x0 & n557 ;
  assign n2409 = n1247 & n2408 ;
  assign n2410 = ~n2407 & n2409 ;
  assign n2411 = n606 & n2410 ;
  assign n2412 = x7 & ~x12 ;
  assign n2413 = ~n1704 & ~n2412 ;
  assign n2414 = n397 & n2413 ;
  assign n2415 = n2056 & n2414 ;
  assign n2416 = ~x0 & ~n303 ;
  assign n2417 = ~n1770 & ~n2416 ;
  assign n2418 = n1656 & ~n2417 ;
  assign n2419 = n1535 & n2062 ;
  assign n2420 = n91 & n2419 ;
  assign n2421 = ~n2418 & ~n2420 ;
  assign n2422 = n2269 & ~n2421 ;
  assign n2423 = ~n2415 & ~n2422 ;
  assign n2424 = ~n2411 & n2423 ;
  assign n2425 = n2424 ^ x4 ;
  assign n2426 = n2425 ^ n2424 ;
  assign n2427 = n2308 & ~n2323 ;
  assign n2428 = n2427 ^ n2424 ;
  assign n2429 = ~n2426 & ~n2428 ;
  assign n2430 = n2429 ^ n2424 ;
  assign n2431 = n1847 & ~n2430 ;
  assign n2432 = ~n2405 & ~n2431 ;
  assign n2433 = n2363 & n2432 ;
  assign n2434 = x4 & ~x11 ;
  assign n2435 = x6 & n2434 ;
  assign n2436 = n231 & n2435 ;
  assign n2437 = n471 & n606 ;
  assign n2438 = n2436 & n2437 ;
  assign n2439 = n16 & n442 ;
  assign n2440 = ~x9 & x13 ;
  assign n2441 = n606 & ~n2440 ;
  assign n2442 = ~n886 & n2441 ;
  assign n2443 = ~n2086 & ~n2442 ;
  assign n2444 = n2443 ^ x1 ;
  assign n2445 = n2444 ^ n2443 ;
  assign n2446 = x7 & x12 ;
  assign n2447 = ~x9 & n344 ;
  assign n2448 = ~n2446 & ~n2447 ;
  assign n2449 = ~n604 & ~n2448 ;
  assign n2450 = n2449 ^ n2443 ;
  assign n2451 = ~n2445 & ~n2450 ;
  assign n2452 = n2451 ^ n2443 ;
  assign n2453 = n2439 & ~n2452 ;
  assign n2454 = ~n2438 & ~n2453 ;
  assign n2455 = ~x7 & ~n1891 ;
  assign n2456 = ~n1550 & ~n2455 ;
  assign n2457 = n410 & n2456 ;
  assign n2458 = n1707 & n2457 ;
  assign n2459 = n99 & n1550 ;
  assign n2460 = n533 & n2459 ;
  assign n2468 = n255 & n1535 ;
  assign n2461 = n166 & ~n2043 ;
  assign n2462 = n659 & ~n1264 ;
  assign n2463 = ~n1256 & ~n2462 ;
  assign n2464 = ~n2461 & ~n2463 ;
  assign n2465 = n255 & n1025 ;
  assign n2466 = ~n1704 & n2465 ;
  assign n2467 = ~n2464 & ~n2466 ;
  assign n2469 = n2468 ^ n2467 ;
  assign n2470 = n2469 ^ x1 ;
  assign n2477 = n2470 ^ n2469 ;
  assign n2471 = n2470 ^ n300 ;
  assign n2472 = n2471 ^ n2469 ;
  assign n2473 = n2470 ^ n2467 ;
  assign n2474 = n2473 ^ n300 ;
  assign n2475 = n2474 ^ n2472 ;
  assign n2476 = ~n2472 & ~n2475 ;
  assign n2478 = n2477 ^ n2476 ;
  assign n2479 = n2478 ^ n2472 ;
  assign n2480 = n2469 ^ n377 ;
  assign n2481 = n2476 ^ n2472 ;
  assign n2482 = ~n2480 & ~n2481 ;
  assign n2483 = n2482 ^ n2469 ;
  assign n2484 = ~n2479 & ~n2483 ;
  assign n2485 = n2484 ^ n2469 ;
  assign n2486 = n2485 ^ n2468 ;
  assign n2487 = n2486 ^ n2469 ;
  assign n2488 = ~n2460 & ~n2487 ;
  assign n2489 = n16 & ~n2488 ;
  assign n2490 = ~n2458 & ~n2489 ;
  assign n2491 = n2490 ^ x0 ;
  assign n2492 = n2491 ^ n2490 ;
  assign n2493 = n2492 ^ n2454 ;
  assign n2530 = x11 & ~n1891 ;
  assign n2531 = ~n1550 & ~n2530 ;
  assign n2532 = n166 & ~n2531 ;
  assign n2533 = n24 & n855 ;
  assign n2534 = ~n2532 & ~n2533 ;
  assign n2494 = ~n659 & ~n2043 ;
  assign n2495 = n166 & ~n2494 ;
  assign n2496 = n2495 ^ n24 ;
  assign n2497 = n2496 ^ n385 ;
  assign n2505 = n2497 ^ n2496 ;
  assign n2498 = ~n362 & n658 ;
  assign n2499 = n2498 ^ n2497 ;
  assign n2500 = n2499 ^ n2496 ;
  assign n2501 = n2497 ^ n2495 ;
  assign n2502 = n2501 ^ n2498 ;
  assign n2503 = n2502 ^ n2500 ;
  assign n2504 = n2500 & ~n2503 ;
  assign n2506 = n2505 ^ n2504 ;
  assign n2507 = n2506 ^ n2500 ;
  assign n2508 = n2496 ^ n1535 ;
  assign n2509 = n2504 ^ n2500 ;
  assign n2510 = n2508 & n2509 ;
  assign n2511 = n2510 ^ n2496 ;
  assign n2512 = ~n2507 & n2511 ;
  assign n2513 = n2512 ^ n2496 ;
  assign n2514 = n2513 ^ n24 ;
  assign n2515 = n2514 ^ n2496 ;
  assign n2535 = n2534 ^ n2515 ;
  assign n2516 = ~n127 & ~n385 ;
  assign n2517 = n255 & ~n2516 ;
  assign n2518 = ~n1134 & n2517 ;
  assign n2519 = n377 & n1233 ;
  assign n2520 = ~n2518 & ~n2519 ;
  assign n2521 = n2520 ^ x13 ;
  assign n2522 = n2521 ^ n2520 ;
  assign n2523 = n2520 ^ n1135 ;
  assign n2524 = n2523 ^ n2520 ;
  assign n2525 = ~n2522 & n2524 ;
  assign n2526 = n2525 ^ n2520 ;
  assign n2527 = ~x9 & ~n2526 ;
  assign n2528 = n2527 ^ n2520 ;
  assign n2529 = n2528 ^ n2515 ;
  assign n2536 = n2535 ^ n2529 ;
  assign n2537 = n2529 ^ x7 ;
  assign n2538 = n2537 ^ n2529 ;
  assign n2539 = n2536 & ~n2538 ;
  assign n2540 = n2539 ^ n2529 ;
  assign n2541 = ~x1 & ~n2540 ;
  assign n2542 = n2541 ^ n2515 ;
  assign n2543 = n2542 ^ n17 ;
  assign n2544 = n17 & n2543 ;
  assign n2545 = n2544 ^ n2490 ;
  assign n2546 = n2545 ^ n17 ;
  assign n2547 = ~n2493 & ~n2546 ;
  assign n2548 = n2547 ^ n2544 ;
  assign n2549 = n2548 ^ n17 ;
  assign n2550 = n2454 & n2549 ;
  assign n2551 = n2550 ^ n2454 ;
  assign n2552 = n1293 & ~n2551 ;
  assign n2553 = n2433 & ~n2552 ;
  assign n2554 = ~n2282 & n2553 ;
  assign n2555 = ~n2264 & n2554 ;
  assign n2556 = ~n2228 & n2555 ;
  assign n2557 = x14 & ~n2556 ;
  assign n2558 = n658 & n1835 ;
  assign n2559 = n828 & n2558 ;
  assign n2560 = x2 & n658 ;
  assign n2561 = x4 & x11 ;
  assign n2562 = n941 & n2033 ;
  assign n2563 = ~n2561 & ~n2562 ;
  assign n2564 = n27 & ~n2563 ;
  assign n2567 = n64 & n2033 ;
  assign n2565 = x4 & n1817 ;
  assign n2566 = ~n300 & n2565 ;
  assign n2568 = n2567 ^ n2566 ;
  assign n2569 = x1 & n2568 ;
  assign n2570 = n2569 ^ n2567 ;
  assign n2571 = ~n2564 & ~n2570 ;
  assign n2572 = n2560 & ~n2571 ;
  assign n2573 = ~n2559 & ~n2572 ;
  assign n2574 = n1759 & ~n2573 ;
  assign n2575 = n1938 & n2265 ;
  assign n2576 = n1960 & n2575 ;
  assign n2577 = n920 & n2576 ;
  assign n2578 = ~n2574 & ~n2577 ;
  assign n2579 = ~x6 & n142 ;
  assign n2580 = ~x3 & n1711 ;
  assign n2581 = ~n2579 & ~n2580 ;
  assign n2582 = n1982 & ~n2581 ;
  assign n2583 = n470 & n2582 ;
  assign n2584 = ~n2345 & ~n2383 ;
  assign n2585 = n2584 ^ x0 ;
  assign n2586 = n2585 ^ n2584 ;
  assign n2587 = n2586 ^ n2583 ;
  assign n2588 = ~x3 & n1816 ;
  assign n2589 = ~x9 & n125 ;
  assign n2590 = ~n606 & n2242 ;
  assign n2591 = ~n2589 & ~n2590 ;
  assign n2592 = n1817 & ~n2591 ;
  assign n2593 = ~n2588 & ~n2592 ;
  assign n2594 = n2593 ^ n2269 ;
  assign n2595 = n2269 & ~n2594 ;
  assign n2596 = n2595 ^ n2584 ;
  assign n2597 = n2596 ^ n2269 ;
  assign n2598 = n2587 & n2597 ;
  assign n2599 = n2598 ^ n2595 ;
  assign n2600 = n2599 ^ n2269 ;
  assign n2601 = ~n2583 & n2600 ;
  assign n2602 = n2601 ^ n2583 ;
  assign n2605 = n2602 ^ n1579 ;
  assign n2606 = n2605 ^ n2602 ;
  assign n2603 = n2602 ^ n2408 ;
  assign n2604 = n2603 ^ n2602 ;
  assign n2607 = n2606 ^ n2604 ;
  assign n2608 = n1765 & n1872 ;
  assign n2609 = n2608 ^ n2602 ;
  assign n2610 = n2609 ^ n2602 ;
  assign n2611 = n2610 ^ n2606 ;
  assign n2612 = n2606 & n2611 ;
  assign n2613 = n2612 ^ n2606 ;
  assign n2614 = n2607 & n2613 ;
  assign n2615 = n2614 ^ n2612 ;
  assign n2616 = n2615 ^ n2602 ;
  assign n2617 = n2616 ^ n2606 ;
  assign n2618 = ~x13 & n2617 ;
  assign n2619 = n2618 ^ n2602 ;
  assign n2620 = ~n303 & n2619 ;
  assign n2621 = n2578 & ~n2620 ;
  assign n2622 = x6 & n106 ;
  assign n2623 = n1753 & ~n1835 ;
  assign n2624 = ~n180 & n2623 ;
  assign n2625 = ~n2622 & ~n2624 ;
  assign n2626 = n658 & ~n2625 ;
  assign n2627 = ~x4 & ~n1847 ;
  assign n2628 = n106 & ~n2627 ;
  assign n2629 = n1832 & n2628 ;
  assign n2630 = ~n2626 & ~n2629 ;
  assign n2631 = x0 & ~n2630 ;
  assign n2632 = n1753 & n1873 ;
  assign n2633 = n941 & n1722 ;
  assign n2634 = n2105 & n2633 ;
  assign n2635 = x6 & ~x7 ;
  assign n2636 = ~x9 & n2635 ;
  assign n2637 = n442 & n2636 ;
  assign n2638 = ~n2634 & ~n2637 ;
  assign n2639 = ~n2632 & n2638 ;
  assign n2640 = x3 & ~n2639 ;
  assign n2641 = n499 & n1835 ;
  assign n2642 = x6 & x13 ;
  assign n2643 = n2641 & n2642 ;
  assign n2644 = n2413 & n2643 ;
  assign n2645 = ~n2640 & ~n2644 ;
  assign n2646 = ~n2631 & n2645 ;
  assign n2647 = n2646 ^ x3 ;
  assign n2648 = n2647 ^ n2646 ;
  assign n2649 = x0 & x6 ;
  assign n2650 = ~n1866 & ~n1906 ;
  assign n2651 = n2649 & ~n2650 ;
  assign n2652 = ~x4 & x7 ;
  assign n2653 = ~n1704 & ~n2652 ;
  assign n2654 = ~x0 & n1753 ;
  assign n2655 = n941 & n2654 ;
  assign n2656 = n2653 & n2655 ;
  assign n2657 = ~n2651 & ~n2656 ;
  assign n2658 = n2657 ^ n2646 ;
  assign n2659 = n2658 ^ n2646 ;
  assign n2660 = n2648 & ~n2659 ;
  assign n2661 = n2660 ^ n2646 ;
  assign n2662 = ~x11 & ~n2661 ;
  assign n2663 = n2662 ^ n2646 ;
  assign n2664 = n501 & ~n2663 ;
  assign n2665 = n2621 & ~n2664 ;
  assign n2666 = ~n2557 & n2665 ;
  assign n2667 = n2094 & n2666 ;
  assign n2668 = ~n1693 & ~n2667 ;
  assign n2669 = n1712 & n1865 ;
  assign n2670 = ~n1707 & ~n2669 ;
  assign n2671 = n277 & n1207 ;
  assign n2672 = ~n362 & n2671 ;
  assign n2673 = n385 ^ x9 ;
  assign n2674 = x9 ^ x3 ;
  assign n2675 = ~n2673 & ~n2674 ;
  assign n2676 = n2675 ^ x3 ;
  assign n2677 = n2672 & ~n2676 ;
  assign n2678 = n601 & n1673 ;
  assign n2679 = x10 & n2678 ;
  assign n2680 = ~n2677 & ~n2679 ;
  assign n2681 = n540 & ~n2680 ;
  assign n2682 = ~x0 & n281 ;
  assign n2683 = n142 & n385 ;
  assign n2684 = n2682 & n2683 ;
  assign n2685 = x0 & ~x8 ;
  assign n2686 = ~x10 & n2685 ;
  assign n2687 = n362 & n2686 ;
  assign n2688 = n143 & n2687 ;
  assign n2689 = ~n2684 & ~n2688 ;
  assign n2690 = ~n606 & ~n2689 ;
  assign n2691 = ~x5 & n614 ;
  assign n2692 = x7 & n753 ;
  assign n2693 = n306 & n2692 ;
  assign n2694 = n2691 & n2693 ;
  assign n2695 = ~x5 & ~n597 ;
  assign n2696 = n167 & n190 ;
  assign n2697 = n1000 & ~n2696 ;
  assign n2698 = x11 & ~n2697 ;
  assign n2699 = ~n2695 & ~n2698 ;
  assign n2700 = ~n182 & n1944 ;
  assign n2701 = ~n1000 & n1831 ;
  assign n2702 = ~n2700 & ~n2701 ;
  assign n2703 = ~n2699 & ~n2702 ;
  assign n2704 = ~n82 & ~n1132 ;
  assign n2705 = n366 & ~n2704 ;
  assign n2706 = ~n167 & ~n642 ;
  assign n2707 = n202 & n2706 ;
  assign n2708 = ~n2705 & ~n2707 ;
  assign n2709 = x0 & ~x13 ;
  assign n2710 = n747 & n2709 ;
  assign n2711 = ~n2708 & n2710 ;
  assign n2712 = ~n2703 & ~n2711 ;
  assign n2713 = x3 & ~n2712 ;
  assign n2714 = ~n2694 & ~n2713 ;
  assign n2715 = ~n2690 & n2714 ;
  assign n2716 = n2715 ^ x1 ;
  assign n2717 = n2716 ^ n2715 ;
  assign n2718 = n2717 ^ n2681 ;
  assign n2719 = n277 & n434 ;
  assign n2720 = ~x0 & n385 ;
  assign n2721 = n2719 & n2720 ;
  assign n2722 = n2709 ^ n597 ;
  assign n2723 = n2722 ^ x11 ;
  assign n2724 = n366 & n1132 ;
  assign n2725 = n2724 ^ n1944 ;
  assign n2726 = ~n597 & ~n2725 ;
  assign n2727 = n2726 ^ n2724 ;
  assign n2728 = ~n2723 & n2727 ;
  assign n2729 = n2728 ^ n2726 ;
  assign n2730 = n2729 ^ n2724 ;
  assign n2731 = n2730 ^ n597 ;
  assign n2732 = x11 & ~n2731 ;
  assign n2733 = ~n2721 & ~n2732 ;
  assign n2734 = ~x3 & ~n2733 ;
  assign n2735 = ~x8 & n831 ;
  assign n2736 = n693 & n2735 ;
  assign n2737 = n199 & n753 ;
  assign n2738 = n191 & n2737 ;
  assign n2739 = ~n2736 & ~n2738 ;
  assign n2740 = n1704 & ~n2739 ;
  assign n2741 = ~n2734 & ~n2740 ;
  assign n2742 = n2741 ^ x5 ;
  assign n2743 = x5 & ~n2742 ;
  assign n2744 = n2743 ^ n2715 ;
  assign n2745 = n2744 ^ x5 ;
  assign n2746 = n2718 & ~n2745 ;
  assign n2747 = n2746 ^ n2743 ;
  assign n2748 = n2747 ^ x5 ;
  assign n2749 = ~n2681 & n2748 ;
  assign n2750 = n2749 ^ n2681 ;
  assign n2751 = x14 & n2750 ;
  assign n2752 = n27 & n802 ;
  assign n2762 = ~n483 & ~n2685 ;
  assign n2763 = ~n539 & ~n2762 ;
  assign n2760 = n2752 ^ x7 ;
  assign n2753 = n277 & n624 ;
  assign n2754 = n747 ^ x3 ;
  assign n2755 = x3 ^ x1 ;
  assign n2756 = n2754 & n2755 ;
  assign n2757 = n2756 ^ x1 ;
  assign n2758 = n2753 & ~n2757 ;
  assign n2759 = n2758 ^ n2752 ;
  assign n2761 = n2760 ^ n2759 ;
  assign n2764 = n2763 ^ n2761 ;
  assign n2765 = n2764 ^ n2761 ;
  assign n2766 = n2761 ^ n2759 ;
  assign n2767 = n2766 ^ n2752 ;
  assign n2768 = n2765 & ~n2767 ;
  assign n2769 = n2768 ^ n2759 ;
  assign n2770 = n625 & n747 ;
  assign n2771 = x10 & n2770 ;
  assign n2772 = ~n2759 & n2771 ;
  assign n2773 = n2772 ^ n2752 ;
  assign n2774 = ~n2769 & ~n2773 ;
  assign n2775 = n2774 ^ n2772 ;
  assign n2776 = ~n2752 & n2775 ;
  assign n2777 = n2776 ^ n2768 ;
  assign n2778 = n2777 ^ n2758 ;
  assign n2779 = n2778 ^ n2759 ;
  assign n2780 = n1891 & ~n2779 ;
  assign n2781 = n199 & n709 ;
  assign n2782 = n626 & n743 ;
  assign n2783 = n2781 & n2782 ;
  assign n2784 = ~n2780 & ~n2783 ;
  assign n2785 = ~n2751 & n2784 ;
  assign n2786 = x8 & n2770 ;
  assign n2787 = ~n2752 & ~n2786 ;
  assign n2788 = n627 & ~n1355 ;
  assign n2789 = x10 ^ x0 ;
  assign n2790 = n2788 & n2789 ;
  assign n2791 = ~n2787 & n2790 ;
  assign n2792 = n2785 & ~n2791 ;
  assign n2793 = ~n2670 & ~n2792 ;
  assign n2794 = x10 ^ x5 ;
  assign n2795 = n606 ^ x10 ;
  assign n2796 = n2795 ^ n606 ;
  assign n2797 = ~x13 & n605 ;
  assign n2798 = n2797 ^ n606 ;
  assign n2799 = ~n2796 & ~n2798 ;
  assign n2800 = n2799 ^ n606 ;
  assign n2801 = ~n2794 & ~n2800 ;
  assign n2802 = n2801 ^ x5 ;
  assign n2803 = n2802 ^ n2801 ;
  assign n2804 = n29 & n167 ;
  assign n2805 = n2804 ^ n2801 ;
  assign n2806 = n2805 ^ n2801 ;
  assign n2807 = ~n2803 & n2806 ;
  assign n2808 = n2807 ^ n2801 ;
  assign n2809 = ~x8 & n2808 ;
  assign n2810 = n2809 ^ n2801 ;
  assign n2811 = n410 & n2810 ;
  assign n2812 = n16 & n2811 ;
  assign n2813 = ~n432 & ~n2128 ;
  assign n2814 = n137 & ~n2147 ;
  assign n2815 = ~x9 & n1719 ;
  assign n2816 = ~n2814 & ~n2815 ;
  assign n2817 = ~x4 & x13 ;
  assign n2818 = ~x6 & ~x10 ;
  assign n2819 = ~x4 & n2818 ;
  assign n2820 = ~n2817 & ~n2819 ;
  assign n2821 = n202 & n2820 ;
  assign n2822 = n2816 & n2821 ;
  assign n2823 = ~x4 & ~x13 ;
  assign n2824 = ~x5 & n2823 ;
  assign n2825 = x7 & n1718 ;
  assign n2826 = ~n2824 & ~n2825 ;
  assign n2827 = ~x6 & ~x9 ;
  assign n2828 = n23 & n2827 ;
  assign n2829 = ~n2826 & n2828 ;
  assign n2830 = ~n2822 & ~n2829 ;
  assign n2831 = n2269 & ~n2830 ;
  assign n2832 = ~n2813 & n2831 ;
  assign n2843 = x1 & ~x8 ;
  assign n2844 = ~n135 & ~n2843 ;
  assign n2838 = ~x4 & n2827 ;
  assign n2839 = ~x10 & ~n410 ;
  assign n2840 = n2838 & ~n2839 ;
  assign n2841 = n2840 ^ n1694 ;
  assign n2833 = n16 & n281 ;
  assign n2834 = n17 & n230 ;
  assign n2835 = ~n2833 & ~n2834 ;
  assign n2836 = x9 & ~n2835 ;
  assign n2837 = n2836 ^ n1694 ;
  assign n2842 = n2841 ^ n2837 ;
  assign n2845 = n2844 ^ n2842 ;
  assign n2846 = n2845 ^ n2842 ;
  assign n2847 = n2842 ^ n2837 ;
  assign n2848 = n2847 ^ n1694 ;
  assign n2849 = n2846 & n2848 ;
  assign n2850 = n2849 ^ n2837 ;
  assign n2851 = ~n281 & n2837 ;
  assign n2852 = n2851 ^ n1694 ;
  assign n2853 = n2850 & n2852 ;
  assign n2854 = n2853 ^ n2851 ;
  assign n2855 = n1694 & n2854 ;
  assign n2856 = n2855 ^ n2849 ;
  assign n2857 = n2856 ^ n2836 ;
  assign n2858 = n2857 ^ n2837 ;
  assign n2859 = n286 & n2858 ;
  assign n2860 = x6 & ~n597 ;
  assign n2861 = ~x6 & n281 ;
  assign n2862 = ~n606 & n2861 ;
  assign n2863 = ~n2860 & ~n2862 ;
  assign n2864 = n410 & ~n2863 ;
  assign n2865 = n1132 & n1938 ;
  assign n2866 = n329 & n2865 ;
  assign n2867 = ~n2864 & ~n2866 ;
  assign n2868 = n1808 & ~n2867 ;
  assign n2869 = ~x4 & n197 ;
  assign n2870 = n843 & n2843 ;
  assign n2871 = x8 & n2269 ;
  assign n2872 = ~n281 & ~n2871 ;
  assign n2873 = n410 ^ x10 ;
  assign n2874 = n2873 ^ n410 ;
  assign n2875 = n1694 ^ n410 ;
  assign n2876 = n2875 ^ n410 ;
  assign n2877 = n2874 & n2876 ;
  assign n2878 = n2877 ^ n410 ;
  assign n2879 = x9 & ~n2878 ;
  assign n2880 = n2879 ^ n410 ;
  assign n2881 = ~n2872 & n2880 ;
  assign n2882 = ~n2870 & ~n2881 ;
  assign n2883 = n2869 & ~n2882 ;
  assign n2884 = ~x6 & n2883 ;
  assign n2885 = ~n2868 & ~n2884 ;
  assign n2886 = ~n2859 & n2885 ;
  assign n2887 = x13 & ~n2886 ;
  assign n2888 = ~n2832 & ~n2887 ;
  assign n2889 = ~n2812 & n2888 ;
  assign n2890 = x3 & ~n2889 ;
  assign n2891 = n410 & ~n591 ;
  assign n2892 = x13 & n596 ;
  assign n2893 = ~n2707 & ~n2892 ;
  assign n2894 = n2232 & ~n2893 ;
  assign n2895 = n2891 & n2894 ;
  assign n2896 = x0 & ~n2895 ;
  assign n2897 = ~n47 & ~n1000 ;
  assign n2898 = n144 & ~n597 ;
  assign n2899 = ~n2897 & ~n2898 ;
  assign n2900 = n410 & ~n2899 ;
  assign n2901 = ~n614 & ~n1550 ;
  assign n2902 = n1207 & n2269 ;
  assign n2903 = ~n190 & n2902 ;
  assign n2904 = ~n2901 & n2903 ;
  assign n2905 = ~n2900 & ~n2904 ;
  assign n2906 = n2248 & ~n2905 ;
  assign n2907 = n410 & n2825 ;
  assign n2908 = n1891 & n2907 ;
  assign n2909 = ~n385 & n2003 ;
  assign n2910 = n606 ^ x4 ;
  assign n2911 = n362 & n2910 ;
  assign n2912 = ~n2909 & ~n2911 ;
  assign n2913 = n639 & ~n2912 ;
  assign n2914 = ~x1 & n2242 ;
  assign n2915 = n51 & n1579 ;
  assign n2916 = n2914 & n2915 ;
  assign n2917 = ~n2913 & ~n2916 ;
  assign n2918 = ~n2908 & n2917 ;
  assign n2919 = n230 & n1716 ;
  assign n2920 = ~n2918 & n2919 ;
  assign n2921 = ~n2906 & ~n2920 ;
  assign n2922 = n2896 & n2921 ;
  assign n2923 = ~n2890 & n2922 ;
  assign n2924 = x6 & ~x8 ;
  assign n2925 = n830 & n2924 ;
  assign n2926 = n1983 & n2925 ;
  assign n2927 = ~x7 & n1579 ;
  assign n2928 = ~n883 & ~n2927 ;
  assign n2929 = x13 & n2833 ;
  assign n2930 = ~n2928 & n2929 ;
  assign n2931 = ~n2926 & ~n2930 ;
  assign n2932 = n35 & ~n2931 ;
  assign n2933 = n614 & n680 ;
  assign n2934 = x10 & ~n1535 ;
  assign n2935 = x8 ^ x7 ;
  assign n2936 = n2440 ^ x8 ;
  assign n2937 = n2935 & ~n2936 ;
  assign n2938 = n2937 ^ x8 ;
  assign n2939 = n2934 & n2938 ;
  assign n2940 = ~n2933 & ~n2939 ;
  assign n2941 = n1722 & ~n2940 ;
  assign n2942 = x4 & n2860 ;
  assign n2943 = ~x4 & x10 ;
  assign n2944 = n601 & n2635 ;
  assign n2945 = ~x6 & x8 ;
  assign n2946 = n248 & n2945 ;
  assign n2947 = ~n604 & n2946 ;
  assign n2948 = ~n2944 & ~n2947 ;
  assign n2949 = n2943 & ~n2948 ;
  assign n2950 = ~n2942 & ~n2949 ;
  assign n2951 = ~n2941 & n2950 ;
  assign n2952 = n837 & ~n2951 ;
  assign n2953 = ~x6 & x10 ;
  assign n2954 = ~x4 & x8 ;
  assign n2955 = x11 & n2954 ;
  assign n2956 = n2953 & n2955 ;
  assign n2957 = n629 & n2956 ;
  assign n2958 = n51 & n2957 ;
  assign n2959 = ~n2952 & ~n2958 ;
  assign n2960 = n501 & ~n2959 ;
  assign n2961 = x5 & n2099 ;
  assign n2962 = n230 & n2636 ;
  assign n2963 = ~n2862 & ~n2962 ;
  assign n2964 = x13 & ~n2963 ;
  assign n2965 = x13 ^ x6 ;
  assign n2966 = ~n1000 & ~n2965 ;
  assign n2967 = ~n2964 & ~n2966 ;
  assign n2968 = n814 & ~n2967 ;
  assign n2969 = n202 & n1817 ;
  assign n2970 = n2440 & n2969 ;
  assign n2971 = n329 & n2970 ;
  assign n2972 = ~n2968 & ~n2971 ;
  assign n2973 = n2961 & ~n2972 ;
  assign n2974 = x6 & ~x10 ;
  assign n2975 = n98 & n2974 ;
  assign n2976 = n52 & n2975 ;
  assign n2977 = ~x11 & n604 ;
  assign n2978 = ~x7 & ~n22 ;
  assign n2979 = ~n2977 & ~n2978 ;
  assign n2980 = n1939 & ~n2979 ;
  assign n2981 = n2976 & n2980 ;
  assign n2982 = ~x0 & ~n2981 ;
  assign n2983 = n629 & n2975 ;
  assign n2984 = n248 & n1914 ;
  assign n2985 = n960 & n2984 ;
  assign n2986 = ~n2983 & ~n2985 ;
  assign n2987 = n2104 & ~n2986 ;
  assign n2988 = x5 & n2987 ;
  assign n2989 = n2982 & ~n2988 ;
  assign n2990 = ~n2973 & n2989 ;
  assign n2991 = ~n2960 & n2990 ;
  assign n2992 = ~n2932 & n2991 ;
  assign n2993 = x14 & ~n2992 ;
  assign n2994 = ~n2923 & n2993 ;
  assign n2995 = x7 & n470 ;
  assign n2996 = n614 & n2953 ;
  assign n2997 = n2033 & n2996 ;
  assign n2998 = n141 & n2997 ;
  assign n2999 = n1808 & n2996 ;
  assign n3000 = x4 & ~x8 ;
  assign n3001 = n2147 & n3000 ;
  assign n3002 = n432 & n3001 ;
  assign n3003 = ~n2999 & ~n3002 ;
  assign n3004 = n837 & ~n3003 ;
  assign n3005 = x8 & n843 ;
  assign n3006 = n2229 & n3005 ;
  assign n3007 = ~n3004 & ~n3006 ;
  assign n3008 = ~n2998 & n3007 ;
  assign n3009 = n2995 & ~n3008 ;
  assign n3010 = n2229 & n2719 ;
  assign n3011 = n202 & n432 ;
  assign n3012 = n1939 & n2147 ;
  assign n3013 = n3011 & n3012 ;
  assign n3014 = ~n3010 & ~n3013 ;
  assign n3015 = x11 ^ x0 ;
  assign n3016 = ~n3014 & n3015 ;
  assign n3017 = x4 & n2649 ;
  assign n3018 = n1459 & n2589 ;
  assign n3019 = n3017 & n3018 ;
  assign n3020 = n3019 ^ x3 ;
  assign n3021 = n3020 ^ n3019 ;
  assign n3022 = n3021 ^ n3016 ;
  assign n3023 = ~n1808 & ~n2242 ;
  assign n3024 = n2860 & n3023 ;
  assign n3025 = ~x0 & n3024 ;
  assign n3026 = n534 & n2128 ;
  assign n3027 = n2954 & n3026 ;
  assign n3028 = ~n606 & n3027 ;
  assign n3029 = n230 & n2649 ;
  assign n3030 = n1816 & n3029 ;
  assign n3031 = ~n3028 & ~n3030 ;
  assign n3032 = ~n3025 & n3031 ;
  assign n3033 = n3032 ^ x11 ;
  assign n3034 = ~n3032 & ~n3033 ;
  assign n3035 = n3034 ^ n3019 ;
  assign n3036 = n3035 ^ n3032 ;
  assign n3037 = n3022 & ~n3036 ;
  assign n3038 = n3037 ^ n3034 ;
  assign n3039 = n3038 ^ n3032 ;
  assign n3040 = ~n3016 & ~n3039 ;
  assign n3041 = n3040 ^ n3016 ;
  assign n3042 = x1 & n3041 ;
  assign n3043 = n230 & n739 ;
  assign n3044 = n3012 & n3043 ;
  assign n3045 = ~n22 & n3044 ;
  assign n3046 = ~n3042 & ~n3045 ;
  assign n3047 = ~n3009 & n3046 ;
  assign n3048 = ~n526 & ~n3047 ;
  assign n3049 = x11 & n17 ;
  assign n3050 = n2408 & n3049 ;
  assign n3051 = ~x1 & ~x4 ;
  assign n3052 = n1914 & n3051 ;
  assign n3053 = n2236 & n3052 ;
  assign n3054 = ~n3050 & ~n3053 ;
  assign n3055 = ~n1000 & ~n3054 ;
  assign n3056 = n625 & n794 ;
  assign n3057 = n2836 & n3056 ;
  assign n3058 = n777 & n2953 ;
  assign n3059 = n1667 & n1835 ;
  assign n3060 = ~n22 & n2954 ;
  assign n3061 = x3 & n3060 ;
  assign n3062 = ~n3059 & ~n3061 ;
  assign n3065 = n3062 ^ x4 ;
  assign n3066 = n3065 ^ n3062 ;
  assign n3063 = n3062 ^ n614 ;
  assign n3064 = n3063 ^ n3062 ;
  assign n3067 = n3066 ^ n3064 ;
  assign n3068 = x3 & x11 ;
  assign n3069 = n3068 ^ n3062 ;
  assign n3070 = n3069 ^ n3062 ;
  assign n3071 = n3070 ^ n3066 ;
  assign n3072 = ~n3066 & ~n3071 ;
  assign n3073 = n3072 ^ n3066 ;
  assign n3074 = ~n3067 & ~n3073 ;
  assign n3075 = n3074 ^ n3072 ;
  assign n3076 = n3075 ^ n3062 ;
  assign n3077 = n3076 ^ n3066 ;
  assign n3078 = ~x1 & n3077 ;
  assign n3079 = n3078 ^ n3062 ;
  assign n3080 = n3058 & ~n3079 ;
  assign n3081 = ~n3057 & ~n3080 ;
  assign n3082 = ~n3055 & n3081 ;
  assign n3083 = n3082 ^ x0 ;
  assign n3084 = n3083 ^ x5 ;
  assign n3111 = n3084 ^ n3083 ;
  assign n3085 = x4 & ~x10 ;
  assign n3086 = n1667 & n1896 ;
  assign n3087 = ~n346 & ~n2827 ;
  assign n3088 = x6 & x9 ;
  assign n3089 = ~n105 & ~n3088 ;
  assign n3090 = x1 & ~n3089 ;
  assign n3091 = ~n3087 & n3090 ;
  assign n3092 = ~n3086 & ~n3091 ;
  assign n3093 = ~x3 & ~n3092 ;
  assign n3094 = n1132 & n2294 ;
  assign n3095 = ~n3093 & ~n3094 ;
  assign n3096 = n3085 & ~n3095 ;
  assign n3097 = n286 & n3096 ;
  assign n3098 = x1 & ~x9 ;
  assign n3099 = ~x11 & n3098 ;
  assign n3100 = ~x1 & ~n22 ;
  assign n3101 = ~n3099 & ~n3100 ;
  assign n3102 = n2833 & ~n3101 ;
  assign n3103 = n287 & n3102 ;
  assign n3104 = ~n3097 & ~n3103 ;
  assign n3105 = n3104 ^ n3084 ;
  assign n3106 = n3105 ^ n3083 ;
  assign n3107 = n3084 ^ n3082 ;
  assign n3108 = n3107 ^ n3104 ;
  assign n3109 = n3108 ^ n3106 ;
  assign n3110 = n3106 & ~n3109 ;
  assign n3112 = n3111 ^ n3110 ;
  assign n3113 = n3112 ^ n3106 ;
  assign n3114 = ~x8 & n2974 ;
  assign n3115 = n2343 & n3114 ;
  assign n3116 = ~n2864 & ~n3115 ;
  assign n3117 = n1960 & ~n3116 ;
  assign n3118 = n557 & n2724 ;
  assign n3119 = n3049 & n3118 ;
  assign n3120 = ~n3117 & ~n3119 ;
  assign n3121 = n3120 ^ n3083 ;
  assign n3122 = n3110 ^ n3106 ;
  assign n3123 = ~n3121 & n3122 ;
  assign n3124 = n3123 ^ n3083 ;
  assign n3125 = n3113 & ~n3124 ;
  assign n3126 = n3125 ^ n3083 ;
  assign n3127 = n3126 ^ x0 ;
  assign n3128 = n3127 ^ n3083 ;
  assign n3129 = ~x13 & n3128 ;
  assign n3130 = n624 & n2945 ;
  assign n3131 = ~n3029 & ~n3130 ;
  assign n3132 = n142 & n173 ;
  assign n3133 = n1836 & n3132 ;
  assign n3134 = n180 & n560 ;
  assign n3135 = ~n606 & n3134 ;
  assign n3136 = n2099 & n3135 ;
  assign n3137 = ~n3133 & ~n3136 ;
  assign n3138 = ~n3131 & ~n3137 ;
  assign n3139 = ~x5 & n173 ;
  assign n3140 = ~n167 & ~n190 ;
  assign n3141 = ~n658 & ~n3140 ;
  assign n3142 = n2084 & n3141 ;
  assign n3143 = ~x7 & n1132 ;
  assign n3144 = ~n1567 & ~n3143 ;
  assign n3145 = n2288 & ~n3144 ;
  assign n3146 = ~n3142 & ~n3145 ;
  assign n3147 = n27 & ~n3146 ;
  assign n3148 = n3139 & n3147 ;
  assign n3149 = ~n3138 & ~n3148 ;
  assign n3150 = ~n3129 & n3149 ;
  assign n3151 = ~n3048 & n3150 ;
  assign n3152 = ~n2994 & n3151 ;
  assign n3153 = n255 & ~n3152 ;
  assign n3154 = ~x4 & x14 ;
  assign n3155 = ~x6 & n3154 ;
  assign n3156 = x1 & n915 ;
  assign n3157 = x0 & n405 ;
  assign n3158 = ~n438 & ~n3157 ;
  assign n3159 = ~n253 & ~n3158 ;
  assign n3160 = ~n3156 & ~n3159 ;
  assign n3161 = n3155 & ~n3160 ;
  assign n3162 = ~x0 & ~n526 ;
  assign n3163 = ~n829 & n3162 ;
  assign n3164 = ~n410 & ~n431 ;
  assign n3165 = n442 & ~n3164 ;
  assign n3166 = ~n540 & n1135 ;
  assign n3167 = ~n3165 & ~n3166 ;
  assign n3168 = ~n3163 & n3167 ;
  assign n3169 = n17 & ~n3168 ;
  assign n3170 = ~n3161 & ~n3169 ;
  assign n3171 = ~n597 & ~n3170 ;
  assign n3172 = x6 ^ x4 ;
  assign n3173 = n404 & n540 ;
  assign n3174 = x0 & x7 ;
  assign n3175 = n540 & n794 ;
  assign n3176 = ~n3174 & ~n3175 ;
  assign n3177 = ~n736 & n3176 ;
  assign n3178 = ~n3173 & n3177 ;
  assign n3179 = ~n604 & ~n3178 ;
  assign n3180 = ~n437 & ~n914 ;
  assign n3181 = n1704 & ~n3180 ;
  assign n3182 = ~n3179 & ~n3181 ;
  assign n3183 = n3182 ^ x6 ;
  assign n3184 = n3183 ^ n3182 ;
  assign n3185 = x0 & ~n1959 ;
  assign n3186 = n1681 & n3185 ;
  assign n3187 = n404 & n658 ;
  assign n3188 = x0 & ~x12 ;
  assign n3189 = ~n658 & n3188 ;
  assign n3190 = ~n410 & ~n1608 ;
  assign n3191 = n3189 & n3190 ;
  assign n3192 = ~n1891 & n2412 ;
  assign n3193 = x11 & n1535 ;
  assign n3194 = ~x0 & ~n3193 ;
  assign n3195 = ~n388 & ~n736 ;
  assign n3196 = ~n1550 & n3195 ;
  assign n3197 = n3194 & ~n3196 ;
  assign n3198 = ~n3192 & n3197 ;
  assign n3199 = ~n3191 & ~n3198 ;
  assign n3200 = ~x1 & n890 ;
  assign n3201 = ~n2269 & ~n3200 ;
  assign n3202 = ~n3199 & n3201 ;
  assign n3203 = x14 & n3202 ;
  assign n3204 = ~n3187 & n3203 ;
  assign n3205 = ~n3186 & ~n3204 ;
  assign n3206 = n3205 ^ n3182 ;
  assign n3207 = ~n3184 & n3206 ;
  assign n3208 = n3207 ^ n3182 ;
  assign n3209 = ~n3172 & ~n3208 ;
  assign n3210 = n281 & n3209 ;
  assign n3211 = n16 & n306 ;
  assign n3212 = x6 & n1872 ;
  assign n3213 = ~x10 & n3212 ;
  assign n3214 = ~n3211 & ~n3213 ;
  assign n3215 = n850 & ~n3214 ;
  assign n3216 = x12 & n3085 ;
  assign n3217 = n739 & n3216 ;
  assign n3218 = n2307 & n3217 ;
  assign n3219 = ~n577 & ~n695 ;
  assign n3220 = n17 & n470 ;
  assign n3221 = n237 & n3220 ;
  assign n3222 = ~n3219 & n3221 ;
  assign n3223 = ~n3218 & ~n3222 ;
  assign n3224 = ~n3215 & n3223 ;
  assign n3225 = n518 & ~n3224 ;
  assign n3226 = ~x9 & n3225 ;
  assign n3227 = n1192 & n2823 ;
  assign n3228 = ~x0 & n3227 ;
  assign n3229 = ~x6 & ~x11 ;
  assign n3230 = n112 & n3229 ;
  assign n3231 = n167 & n3230 ;
  assign n3232 = n3228 & n3231 ;
  assign n3233 = ~x10 & n1192 ;
  assign n3234 = ~x0 & x4 ;
  assign n3235 = n3088 & n3234 ;
  assign n3236 = ~n165 & n3235 ;
  assign n3237 = ~n736 & ~n1608 ;
  assign n3238 = n385 & n3237 ;
  assign n3239 = n2084 & n3238 ;
  assign n3240 = ~n3236 & ~n3239 ;
  assign n3241 = n3233 & ~n3240 ;
  assign n3242 = n1013 & n3220 ;
  assign n3243 = x0 & x4 ;
  assign n3244 = n167 & n3243 ;
  assign n3245 = n1938 & n3244 ;
  assign n3246 = ~n3242 & ~n3245 ;
  assign n3247 = ~n3241 & n3246 ;
  assign n3248 = n3247 ^ x8 ;
  assign n3249 = n3248 ^ n3247 ;
  assign n3250 = ~x7 & n17 ;
  assign n3251 = x9 ^ x1 ;
  assign n3252 = n3251 ^ n646 ;
  assign n3253 = x0 & n3252 ;
  assign n3254 = n3253 ^ n646 ;
  assign n3255 = n3250 & n3254 ;
  assign n3256 = n3255 ^ n3247 ;
  assign n3257 = n3249 & ~n3256 ;
  assign n3258 = n3257 ^ n3247 ;
  assign n3259 = ~n3232 & n3258 ;
  assign n3260 = ~x2 & n3259 ;
  assign n3261 = ~n3226 & n3260 ;
  assign n3262 = ~n3210 & n3261 ;
  assign n3263 = n913 & n992 ;
  assign n3264 = ~n470 & ~n3263 ;
  assign n3265 = n281 & ~n3264 ;
  assign n3266 = n1141 ^ x12 ;
  assign n3267 = ~x1 & ~n3266 ;
  assign n3268 = n3267 ^ x12 ;
  assign n3269 = n2686 & n3268 ;
  assign n3270 = x14 & n3269 ;
  assign n3271 = ~n3265 & ~n3270 ;
  assign n3272 = n2838 & ~n3271 ;
  assign n3273 = n2834 & n3173 ;
  assign n3274 = n16 & n431 ;
  assign n3275 = ~n2288 & ~n3274 ;
  assign n3276 = n281 & ~n3275 ;
  assign n3277 = n17 & ~n343 ;
  assign n3278 = n1113 & n2819 ;
  assign n3279 = ~n3277 & ~n3278 ;
  assign n3280 = n2685 & ~n3279 ;
  assign n3281 = ~n3276 & ~n3280 ;
  assign n3282 = n2347 & ~n3281 ;
  assign n3283 = ~n3273 & ~n3282 ;
  assign n3284 = ~n3272 & n3283 ;
  assign n3285 = ~x9 & n17 ;
  assign n3286 = ~x10 & ~n1113 ;
  assign n3287 = ~x1 & ~n3286 ;
  assign n3288 = n431 ^ x0 ;
  assign n3289 = n1507 ^ n431 ;
  assign n3290 = n3289 ^ n431 ;
  assign n3291 = n3288 & ~n3290 ;
  assign n3292 = n3291 ^ n431 ;
  assign n3293 = ~n3287 & ~n3292 ;
  assign n3294 = n3293 ^ x8 ;
  assign n3295 = n3294 ^ n3293 ;
  assign n3296 = ~n236 & ~n343 ;
  assign n3297 = n543 & n3296 ;
  assign n3298 = n3297 ^ n3293 ;
  assign n3299 = n3295 & ~n3298 ;
  assign n3300 = n3299 ^ n3293 ;
  assign n3301 = n3285 & ~n3300 ;
  assign n3302 = n3284 & ~n3301 ;
  assign n3303 = x7 & ~n3302 ;
  assign n3304 = ~n1580 & n3043 ;
  assign n3305 = ~n1141 & n3304 ;
  assign n3306 = n80 & n483 ;
  assign n3307 = x11 & n3306 ;
  assign n3308 = ~x10 & n170 ;
  assign n3309 = n2685 & n3308 ;
  assign n3310 = ~n3307 & ~n3309 ;
  assign n3311 = n48 & ~n3310 ;
  assign n3312 = n1684 & n1886 ;
  assign n3313 = ~x9 & n199 ;
  assign n3314 = n708 & n3313 ;
  assign n3315 = ~n3312 & ~n3314 ;
  assign n3316 = ~n1371 & n3315 ;
  assign n3317 = n540 & ~n3316 ;
  assign n3318 = ~n3311 & ~n3317 ;
  assign n3319 = ~n3305 & n3318 ;
  assign n3320 = n3155 & ~n3319 ;
  assign n3321 = n79 & n148 ;
  assign n3322 = ~n960 & ~n3321 ;
  assign n3323 = ~x7 & ~n3322 ;
  assign n3324 = ~x8 & n59 ;
  assign n3325 = n799 & n3324 ;
  assign n3326 = ~n3323 & ~n3325 ;
  assign n3327 = x1 & n2084 ;
  assign n3328 = ~n3326 & n3327 ;
  assign n3329 = ~n3320 & ~n3328 ;
  assign n3330 = ~n1507 & ~n2762 ;
  assign n3331 = n1058 & n2843 ;
  assign n3332 = ~n3330 & ~n3331 ;
  assign n3333 = n3332 ^ x9 ;
  assign n3334 = n3333 ^ n3332 ;
  assign n3335 = n3334 ^ n3250 ;
  assign n3336 = n19 & n1915 ;
  assign n3337 = n3250 ^ n1459 ;
  assign n3338 = n3336 & ~n3337 ;
  assign n3339 = n3338 ^ n3332 ;
  assign n3340 = ~n3335 & ~n3339 ;
  assign n3341 = n3340 ^ n3338 ;
  assign n3342 = ~n3250 & n3341 ;
  assign n3343 = n3342 ^ n3338 ;
  assign n3344 = n3343 ^ n3340 ;
  assign n3345 = n3329 & ~n3344 ;
  assign n3346 = ~n1190 & n1684 ;
  assign n3347 = ~n1041 & ~n3346 ;
  assign n3348 = n470 & ~n3347 ;
  assign n3349 = n16 & n3348 ;
  assign n3350 = ~x8 & n17 ;
  assign n3351 = ~n830 & ~n988 ;
  assign n3352 = n3350 & ~n3351 ;
  assign n3353 = ~n2833 & ~n3352 ;
  assign n3354 = n404 & ~n3353 ;
  assign n3355 = x4 & x8 ;
  assign n3356 = ~n1684 & ~n3355 ;
  assign n3357 = ~n18 & ~n3356 ;
  assign n3358 = n2943 & n3229 ;
  assign n3359 = n530 & n3358 ;
  assign n3360 = ~n3357 & ~n3359 ;
  assign n3361 = ~n3354 & n3360 ;
  assign n3362 = n543 & ~n3361 ;
  assign n3363 = n230 & n431 ;
  assign n3364 = n3017 & n3363 ;
  assign n3365 = x6 & ~x11 ;
  assign n3366 = n261 & n3085 ;
  assign n3367 = n3365 & n3366 ;
  assign n3368 = ~n2833 & ~n3367 ;
  assign n3369 = n437 & ~n3368 ;
  assign n3370 = n713 & n3350 ;
  assign n3371 = ~n3369 & ~n3370 ;
  assign n3372 = ~n3364 & n3371 ;
  assign n3373 = ~n3362 & n3372 ;
  assign n3374 = ~n3349 & n3373 ;
  assign n3375 = n1535 & ~n3374 ;
  assign n3376 = n3345 & ~n3375 ;
  assign n3377 = x2 & n3376 ;
  assign n3378 = ~n3303 & n3377 ;
  assign n3379 = ~n3262 & ~n3378 ;
  assign n3380 = ~n134 & ~n253 ;
  assign n3381 = x14 & ~n410 ;
  assign n3382 = ~n912 & n3381 ;
  assign n3383 = ~n3380 & n3382 ;
  assign n3384 = x1 & ~n978 ;
  assign n3385 = ~n344 & n3384 ;
  assign n3386 = n3385 ^ n405 ;
  assign n3387 = n3386 ^ n3385 ;
  assign n3388 = n3387 ^ x2 ;
  assign n3389 = x13 ^ x1 ;
  assign n3390 = ~x13 & n3389 ;
  assign n3391 = n3390 ^ n3385 ;
  assign n3392 = n3391 ^ x13 ;
  assign n3393 = n3388 & n3392 ;
  assign n3394 = n3393 ^ n3390 ;
  assign n3395 = n3394 ^ x13 ;
  assign n3396 = x2 & ~n3395 ;
  assign n3397 = ~n3383 & ~n3396 ;
  assign n3398 = x0 & ~n3397 ;
  assign n3399 = x14 & n442 ;
  assign n3400 = n3268 & n3399 ;
  assign n3401 = ~n3398 & ~n3400 ;
  assign n3402 = n16 & ~n3401 ;
  assign n3403 = n438 & n2435 ;
  assign n3404 = ~n3402 & ~n3403 ;
  assign n3405 = ~n1000 & ~n3404 ;
  assign n3406 = x4 & x12 ;
  assign n3407 = n167 & n890 ;
  assign n3408 = x0 & ~x10 ;
  assign n3409 = ~n606 & n3408 ;
  assign n3410 = ~n3407 & ~n3409 ;
  assign n3411 = n129 & n2924 ;
  assign n3412 = ~n3410 & n3411 ;
  assign n3413 = n3406 & n3412 ;
  assign n3414 = ~n3405 & ~n3413 ;
  assign n3415 = ~n3379 & n3414 ;
  assign n3416 = ~n3171 & n3415 ;
  assign n3417 = n1293 & ~n3416 ;
  assign n3418 = ~n3153 & ~n3417 ;
  assign n3419 = n265 & n2943 ;
  assign n3420 = ~n3366 & ~n3419 ;
  assign n3421 = ~n3132 & ~n3134 ;
  assign n3422 = n2112 & ~n3421 ;
  assign n3423 = ~x3 & n2147 ;
  assign n3424 = n570 & n3423 ;
  assign n3425 = ~n513 & n3424 ;
  assign n3426 = ~n3422 & ~n3425 ;
  assign n3427 = n1704 & ~n3426 ;
  assign n3428 = ~x3 & n286 ;
  assign n3429 = ~x0 & ~n2642 ;
  assign n3430 = n3428 & ~n3429 ;
  assign n3431 = n21 & ~n2649 ;
  assign n3432 = n69 & n3431 ;
  assign n3433 = n3430 & n3432 ;
  assign n3434 = n141 & n362 ;
  assign n3435 = ~n2683 & ~n3434 ;
  assign n3436 = n605 & n2001 ;
  assign n3437 = n540 & n3436 ;
  assign n3438 = n1704 & n2112 ;
  assign n3439 = ~n3437 & ~n3438 ;
  assign n3440 = ~n3435 & ~n3439 ;
  assign n3441 = ~n3433 & ~n3440 ;
  assign n3442 = n2498 ^ n2399 ;
  assign n3443 = x2 & n3442 ;
  assign n3444 = n3443 ^ n2399 ;
  assign n3445 = n753 & n3444 ;
  assign n3446 = n2147 & n3445 ;
  assign n3447 = n512 & n3135 ;
  assign n3448 = n2299 & n3139 ;
  assign n3449 = n3448 ^ n1704 ;
  assign n3450 = n3449 ^ n3448 ;
  assign n3451 = n385 & n940 ;
  assign n3452 = n3451 ^ n362 ;
  assign n3453 = n3452 ^ n3451 ;
  assign n3454 = n3451 ^ n944 ;
  assign n3455 = n3454 ^ n3451 ;
  assign n3456 = n3453 & n3455 ;
  assign n3457 = n3456 ^ n3451 ;
  assign n3458 = ~x5 & n3457 ;
  assign n3459 = n3458 ^ n3451 ;
  assign n3460 = n3459 ^ n3448 ;
  assign n3461 = ~n3450 & n3460 ;
  assign n3462 = n3461 ^ n3448 ;
  assign n3463 = ~n3447 & ~n3462 ;
  assign n3464 = n3463 ^ x6 ;
  assign n3465 = n3464 ^ n3463 ;
  assign n3466 = ~x2 & n142 ;
  assign n3467 = x0 & ~n385 ;
  assign n3468 = n1535 & n3467 ;
  assign n3469 = n743 & n1626 ;
  assign n3470 = ~n3468 & ~n3469 ;
  assign n3471 = n3466 & ~n3470 ;
  assign n3472 = n3471 ^ n3463 ;
  assign n3473 = n3465 & ~n3472 ;
  assign n3474 = n3473 ^ n3463 ;
  assign n3475 = ~n3446 & n3474 ;
  assign n3476 = n3475 ^ x1 ;
  assign n3477 = n3476 ^ n3475 ;
  assign n3478 = n3477 ^ n3441 ;
  assign n3479 = n605 & n3423 ;
  assign n3480 = n344 & n3479 ;
  assign n3481 = ~n1891 & ~n3229 ;
  assign n3482 = x3 & n556 ;
  assign n3483 = ~x6 & x9 ;
  assign n3484 = ~n173 & ~n3483 ;
  assign n3485 = n3482 & n3484 ;
  assign n3486 = ~n3481 & n3485 ;
  assign n3487 = ~n3480 & ~n3486 ;
  assign n3488 = ~x11 & n1891 ;
  assign n3489 = ~n2447 & ~n3488 ;
  assign n3490 = x9 ^ x6 ;
  assign n3491 = ~n3489 & n3490 ;
  assign n3492 = n3428 & n3491 ;
  assign n3493 = n3487 & ~n3492 ;
  assign n3494 = n3493 ^ n513 ;
  assign n3495 = ~n3493 & n3494 ;
  assign n3496 = n3495 ^ n3475 ;
  assign n3497 = n3496 ^ n3493 ;
  assign n3498 = ~n3478 & n3497 ;
  assign n3499 = n3498 ^ n3495 ;
  assign n3500 = n3499 ^ n3493 ;
  assign n3501 = n3441 & ~n3500 ;
  assign n3502 = n3501 ^ n3441 ;
  assign n3503 = x14 & ~n3502 ;
  assign n3504 = n540 & n1232 ;
  assign n3505 = n512 & ~n1694 ;
  assign n3506 = ~n3504 & ~n3505 ;
  assign n3507 = n556 & n591 ;
  assign n3508 = n1817 & n3507 ;
  assign n3509 = ~n3506 & n3508 ;
  assign n3510 = n173 & n658 ;
  assign n3511 = n141 & n3510 ;
  assign n3512 = n2240 & n3511 ;
  assign n3513 = n1697 & n2266 ;
  assign n3514 = n362 & n3513 ;
  assign n3515 = ~n3512 & ~n3514 ;
  assign n3516 = ~n3509 & n3515 ;
  assign n3517 = ~n3503 & n3516 ;
  assign n3518 = ~n3427 & n3517 ;
  assign n3519 = ~n3420 & ~n3518 ;
  assign n3520 = n23 & n992 ;
  assign n3521 = ~x0 & n1705 ;
  assign n3522 = n128 & n2083 ;
  assign n3523 = ~n3521 & ~n3522 ;
  assign n3524 = n3520 & ~n3523 ;
  assign n3525 = n79 & ~n526 ;
  assign n3526 = n443 & n3525 ;
  assign n3527 = n920 & n3324 ;
  assign n3528 = ~n3526 & ~n3527 ;
  assign n3529 = n1946 & ~n3528 ;
  assign n3530 = ~n3524 & ~n3529 ;
  assign n3531 = n1632 & ~n3530 ;
  assign n3532 = n944 & n1731 ;
  assign n3533 = n307 ^ x12 ;
  assign n3534 = n3533 ^ n79 ;
  assign n3535 = n3534 ^ n307 ;
  assign n3536 = n3535 ^ n3534 ;
  assign n3537 = ~x8 & n1147 ;
  assign n3538 = n3537 ^ n3534 ;
  assign n3539 = n3538 ^ n3533 ;
  assign n3540 = n3536 & ~n3539 ;
  assign n3541 = n3540 ^ n3537 ;
  assign n3542 = n3351 & ~n3537 ;
  assign n3543 = n3542 ^ n3533 ;
  assign n3544 = ~n3541 & n3543 ;
  assign n3545 = n3544 ^ n3542 ;
  assign n3546 = n3533 & n3545 ;
  assign n3547 = n3546 ^ n3540 ;
  assign n3548 = n3547 ^ x12 ;
  assign n3549 = n3548 ^ n3537 ;
  assign n3550 = n3532 & n3549 ;
  assign n3551 = ~n3531 & ~n3550 ;
  assign n3552 = n3551 ^ x7 ;
  assign n3553 = n3552 ^ n3551 ;
  assign n3554 = ~n54 & n2083 ;
  assign n3555 = ~x13 & n3234 ;
  assign n3556 = ~n1293 & n3555 ;
  assign n3557 = ~n3554 & ~n3556 ;
  assign n3558 = n992 & ~n3557 ;
  assign n3559 = n581 & n3234 ;
  assign n3560 = x3 & ~x12 ;
  assign n3561 = n2242 & n3560 ;
  assign n3562 = n1944 & n3561 ;
  assign n3563 = ~n3559 & ~n3562 ;
  assign n3564 = ~n3558 & n3563 ;
  assign n3565 = n23 & ~n3564 ;
  assign n3566 = n281 & n2136 ;
  assign n3567 = n992 & n3566 ;
  assign n3568 = x3 & n3567 ;
  assign n3569 = x5 & n3000 ;
  assign n3570 = n19 & n80 ;
  assign n3571 = n3569 & n3570 ;
  assign n3572 = n831 & n1808 ;
  assign n3573 = n3324 & n3572 ;
  assign n3574 = ~n3571 & ~n3573 ;
  assign n3575 = ~n3568 & n3574 ;
  assign n3576 = ~n3565 & n3575 ;
  assign n3577 = n181 & ~n3576 ;
  assign n3578 = n812 & n2298 ;
  assign n3579 = n108 & n3578 ;
  assign n3580 = x10 ^ x8 ;
  assign n3581 = n2789 ^ x0 ;
  assign n3582 = n3162 ^ x0 ;
  assign n3583 = n3581 & n3582 ;
  assign n3584 = n3583 ^ x0 ;
  assign n3585 = n3580 & n3584 ;
  assign n3586 = n3579 & n3585 ;
  assign n3587 = n312 & n2943 ;
  assign n3588 = ~x0 & ~n231 ;
  assign n3589 = n3587 & n3588 ;
  assign n3590 = ~x10 & n3000 ;
  assign n3591 = ~x14 & n377 ;
  assign n3592 = n3590 & ~n3591 ;
  assign n3593 = n2247 & n3592 ;
  assign n3594 = ~n3589 & ~n3593 ;
  assign n3595 = n128 & ~n3594 ;
  assign n3596 = n142 & n920 ;
  assign n3597 = ~n1190 & n3590 ;
  assign n3598 = n3596 & n3597 ;
  assign n3599 = ~n3595 & ~n3598 ;
  assign n3600 = x9 & ~n3599 ;
  assign n3601 = ~x5 & n1939 ;
  assign n3602 = n2062 & n3537 ;
  assign n3603 = n3601 & n3602 ;
  assign n3604 = ~n3600 & ~n3603 ;
  assign n3605 = ~n3586 & n3604 ;
  assign n3606 = ~n3577 & n3605 ;
  assign n3607 = n3606 ^ n3551 ;
  assign n3608 = n3553 & n3607 ;
  assign n3609 = n3608 ^ n3551 ;
  assign n3610 = x6 & ~n3609 ;
  assign n3611 = x10 & n2232 ;
  assign n3612 = ~n2943 & ~n3085 ;
  assign n3613 = n142 & ~n3612 ;
  assign n3614 = x6 & n3613 ;
  assign n3615 = ~n3611 & ~n3614 ;
  assign n3616 = ~x12 & n529 ;
  assign n3617 = ~x0 & n452 ;
  assign n3618 = n3616 & n3617 ;
  assign n3619 = ~n3615 & n3618 ;
  assign n3620 = n432 & n1364 ;
  assign n3621 = n60 & n3620 ;
  assign n3622 = ~x0 & n526 ;
  assign n3623 = n3621 & ~n3622 ;
  assign n3624 = x12 & n1132 ;
  assign n3625 = n624 & n3624 ;
  assign n3626 = x0 & ~x9 ;
  assign n3627 = n167 & ~n526 ;
  assign n3628 = x0 & ~n3351 ;
  assign n3629 = ~n3627 & ~n3628 ;
  assign n3630 = n265 & ~n3629 ;
  assign n3631 = ~n3626 & n3630 ;
  assign n3632 = ~n3625 & ~n3631 ;
  assign n3633 = n1805 & ~n3632 ;
  assign n3634 = ~n3623 & ~n3633 ;
  assign n3635 = n2565 & ~n3634 ;
  assign n3636 = n642 & n1835 ;
  assign n3637 = n167 & n1960 ;
  assign n3638 = ~n3636 & ~n3637 ;
  assign n3639 = ~x2 & n312 ;
  assign n3640 = x12 & n3639 ;
  assign n3641 = ~n3638 & n3640 ;
  assign n3642 = n529 & n3000 ;
  assign n3643 = n1960 & n3313 ;
  assign n3644 = ~n3642 & ~n3643 ;
  assign n3645 = n80 & n1805 ;
  assign n3646 = ~n3644 & n3645 ;
  assign n3647 = ~n434 & ~n989 ;
  assign n3648 = n1939 & ~n3647 ;
  assign n3649 = ~x4 & n629 ;
  assign n3650 = n1147 & n3649 ;
  assign n3651 = ~n3648 & ~n3650 ;
  assign n3652 = n60 & n1627 ;
  assign n3653 = ~n3651 & n3652 ;
  assign n3654 = ~n3646 & ~n3653 ;
  assign n3655 = ~n3641 & n3654 ;
  assign n3656 = n1776 & ~n3655 ;
  assign n3657 = ~n3635 & ~n3656 ;
  assign n3658 = n3657 ^ x7 ;
  assign n3659 = n3658 ^ n3657 ;
  assign n3660 = n3659 ^ n3619 ;
  assign n3661 = n992 & n3639 ;
  assign n3662 = n218 & n313 ;
  assign n3663 = n527 & n3662 ;
  assign n3664 = ~n3661 & ~n3663 ;
  assign n3665 = n624 & ~n3664 ;
  assign n3666 = n79 & n3596 ;
  assign n3667 = x8 & n3666 ;
  assign n3668 = ~n3665 & ~n3667 ;
  assign n3669 = n1728 & ~n3668 ;
  assign n3670 = n142 & n499 ;
  assign n3671 = n59 & n614 ;
  assign n3672 = n3670 & n3671 ;
  assign n3673 = ~x3 & n3324 ;
  assign n3674 = ~n3520 & ~n3673 ;
  assign n3675 = n3626 & ~n3674 ;
  assign n3676 = n1805 & n3675 ;
  assign n3677 = ~n3672 & ~n3676 ;
  assign n3678 = n3677 ^ x4 ;
  assign n3679 = n3678 ^ n3677 ;
  assign n3680 = n3679 ^ n3669 ;
  assign n3681 = n614 & ~n1460 ;
  assign n3682 = n303 & n764 ;
  assign n3683 = n3681 & n3682 ;
  assign n3684 = x2 & x5 ;
  assign n3685 = ~x0 & n3684 ;
  assign n3686 = n1550 & n1577 ;
  assign n3687 = n1192 & n3686 ;
  assign n3688 = n3685 & n3687 ;
  assign n3689 = ~n3683 & ~n3688 ;
  assign n3690 = n3689 ^ x10 ;
  assign n3691 = ~n3689 & ~n3690 ;
  assign n3692 = n3691 ^ n3677 ;
  assign n3693 = n3692 ^ n3689 ;
  assign n3694 = n3680 & n3693 ;
  assign n3695 = n3694 ^ n3691 ;
  assign n3696 = n3695 ^ n3689 ;
  assign n3697 = ~n3669 & ~n3696 ;
  assign n3698 = n3697 ^ n3669 ;
  assign n3699 = n3698 ^ x6 ;
  assign n3700 = n3698 & ~n3699 ;
  assign n3701 = n3700 ^ n3657 ;
  assign n3702 = n3701 ^ n3698 ;
  assign n3703 = ~n3660 & ~n3702 ;
  assign n3704 = n3703 ^ n3700 ;
  assign n3705 = n3704 ^ n3698 ;
  assign n3706 = ~n3619 & n3705 ;
  assign n3707 = n3706 ^ n3619 ;
  assign n3708 = ~n3610 & ~n3707 ;
  assign n3709 = ~n1694 & ~n3708 ;
  assign n3710 = ~n3519 & ~n3709 ;
  assign n3711 = n3418 & n3710 ;
  assign n3712 = ~n2793 & n3711 ;
  assign n3713 = ~n2668 & n3712 ;
  assign n3714 = ~n1692 & n3713 ;
  assign n3715 = n1718 & n1776 ;
  assign n3716 = n254 & n3715 ;
  assign n3717 = n596 & n3716 ;
  assign n3718 = ~x6 & n920 ;
  assign n3719 = n1853 & n3718 ;
  assign n3720 = n82 & ~n513 ;
  assign n3721 = x2 & ~n1944 ;
  assign n3722 = ~n19 & ~n3721 ;
  assign n3723 = n1132 & ~n3722 ;
  assign n3724 = ~n3720 & ~n3723 ;
  assign n3727 = n3724 ^ n1891 ;
  assign n3728 = n3727 ^ n3724 ;
  assign n3725 = n3724 ^ n518 ;
  assign n3726 = n3725 ^ n3724 ;
  assign n3729 = n3728 ^ n3726 ;
  assign n3730 = n3724 ^ n499 ;
  assign n3731 = n3730 ^ n3724 ;
  assign n3732 = n3731 ^ n3728 ;
  assign n3733 = n3728 & n3732 ;
  assign n3734 = n3733 ^ n3728 ;
  assign n3735 = n3729 & n3734 ;
  assign n3736 = n3735 ^ n3733 ;
  assign n3737 = n3736 ^ n3724 ;
  assign n3738 = n3737 ^ n3728 ;
  assign n3739 = ~x12 & ~n3738 ;
  assign n3740 = n3739 ^ n3724 ;
  assign n3741 = x6 & ~n3740 ;
  assign n3742 = ~n3719 & ~n3741 ;
  assign n3743 = n539 & ~n3742 ;
  assign n3744 = n171 & n1104 ;
  assign n3745 = ~x8 & n3744 ;
  assign n3746 = x12 & n614 ;
  assign n3747 = ~n3745 & ~n3746 ;
  assign n3748 = n1776 & ~n3747 ;
  assign n3749 = n65 & n3748 ;
  assign n3750 = ~x0 & n3745 ;
  assign n3751 = n2001 & n3750 ;
  assign n3752 = n2654 & n3746 ;
  assign n3753 = ~n3751 & ~n3752 ;
  assign n3754 = x10 & ~n3753 ;
  assign n3755 = n3624 & n3718 ;
  assign n3756 = x4 & ~n3755 ;
  assign n3757 = ~x8 & ~x12 ;
  assign n3758 = x0 & n3757 ;
  assign n3759 = n3088 ^ x6 ;
  assign n3760 = n3759 ^ n3088 ;
  assign n3761 = n3088 ^ n1550 ;
  assign n3762 = n3761 ^ n3088 ;
  assign n3763 = ~n3760 & n3762 ;
  assign n3764 = n3763 ^ n3088 ;
  assign n3765 = x2 & n3764 ;
  assign n3766 = n3765 ^ n3088 ;
  assign n3767 = n3758 & n3766 ;
  assign n3768 = ~x0 & x12 ;
  assign n3769 = n1753 & n3768 ;
  assign n3770 = n82 & n3769 ;
  assign n3771 = ~n3767 & ~n3770 ;
  assign n3772 = n988 & ~n3771 ;
  assign n3773 = n3756 & ~n3772 ;
  assign n3774 = ~n3754 & n3773 ;
  assign n3775 = ~n3749 & n3774 ;
  assign n3776 = ~n2242 & ~n3775 ;
  assign n3777 = ~n3743 & ~n3776 ;
  assign n3778 = ~x6 & x14 ;
  assign n3779 = ~x0 & n1805 ;
  assign n3780 = n3671 & n3779 ;
  assign n3781 = ~x9 & n205 ;
  assign n3782 = n1944 ^ n1770 ;
  assign n3783 = n3782 ^ n1770 ;
  assign n3784 = n1770 ^ n254 ;
  assign n3785 = n3784 ^ n1770 ;
  assign n3786 = n3783 & n3785 ;
  assign n3787 = n3786 ^ n1770 ;
  assign n3788 = ~x8 & n3787 ;
  assign n3789 = n3788 ^ n1770 ;
  assign n3790 = n3781 & n3789 ;
  assign n3791 = n80 & n452 ;
  assign n3792 = ~n262 & ~n3791 ;
  assign n3793 = n2247 & ~n3792 ;
  assign n3794 = n205 & n483 ;
  assign n3795 = ~n255 & n3794 ;
  assign n3796 = ~n3793 & ~n3795 ;
  assign n3797 = n1891 & ~n3796 ;
  assign n3798 = ~n3790 & ~n3797 ;
  assign n3799 = ~n3780 & n3798 ;
  assign n3800 = n3778 & ~n3799 ;
  assign n3801 = x12 & n3684 ;
  assign n3802 = n23 & n3626 ;
  assign n3803 = n2704 & n2953 ;
  assign n3804 = ~n1944 & n3803 ;
  assign n3805 = ~n3802 & ~n3804 ;
  assign n3806 = n3801 & ~n3805 ;
  assign n3807 = ~n513 & n2706 ;
  assign n3808 = ~x8 & n642 ;
  assign n3809 = n3721 & n3808 ;
  assign n3810 = ~n3807 & ~n3809 ;
  assign n3813 = n3810 ^ n920 ;
  assign n3814 = n3813 ^ n3810 ;
  assign n3811 = n3810 ^ n591 ;
  assign n3812 = n3811 ^ n3810 ;
  assign n3815 = n3814 ^ n3812 ;
  assign n3816 = n3810 ^ n230 ;
  assign n3817 = n3816 ^ n3810 ;
  assign n3818 = n3817 ^ n3814 ;
  assign n3819 = n3814 & n3818 ;
  assign n3820 = n3819 ^ n3814 ;
  assign n3821 = n3815 & n3820 ;
  assign n3822 = n3821 ^ n3819 ;
  assign n3823 = n3822 ^ n3810 ;
  assign n3824 = n3823 ^ n3814 ;
  assign n3825 = ~x6 & ~n3824 ;
  assign n3826 = n3825 ^ n3810 ;
  assign n3827 = n1627 & ~n3826 ;
  assign n3828 = x6 & x10 ;
  assign n3829 = ~x5 & n3828 ;
  assign n3830 = n525 & n3829 ;
  assign n3831 = ~n513 & n3830 ;
  assign n3832 = ~x4 & ~n3831 ;
  assign n3833 = ~n3827 & n3832 ;
  assign n3834 = ~n3806 & n3833 ;
  assign n3835 = ~n81 & ~n1207 ;
  assign n3836 = n2827 & n3835 ;
  assign n3837 = n917 & n1765 ;
  assign n3838 = ~n3836 & ~n3837 ;
  assign n3839 = ~n513 & ~n3838 ;
  assign n3840 = ~x10 & n1753 ;
  assign n3841 = n2120 & n3840 ;
  assign n3842 = n1632 & n3841 ;
  assign n3843 = ~n3839 & ~n3842 ;
  assign n3844 = n601 & ~n3843 ;
  assign n3845 = n942 & n1132 ;
  assign n3846 = n442 & n1765 ;
  assign n3847 = n3845 & n3846 ;
  assign n3848 = x6 & x8 ;
  assign n3849 = n1247 & n3848 ;
  assign n3850 = n1550 & n3849 ;
  assign n3851 = ~n534 & ~n920 ;
  assign n3852 = ~n65 & ~n203 ;
  assign n3853 = ~x0 & n3852 ;
  assign n3854 = n3851 & ~n3853 ;
  assign n3855 = n3850 & n3854 ;
  assign n3856 = ~n3847 & ~n3855 ;
  assign n3857 = ~n3844 & n3856 ;
  assign n3858 = x14 & ~n3857 ;
  assign n3859 = n3834 & ~n3858 ;
  assign n3860 = ~n3800 & n3859 ;
  assign n3861 = ~n3777 & ~n3860 ;
  assign n3862 = n499 & n1765 ;
  assign n3863 = ~n1106 & n3862 ;
  assign n3864 = x6 & n1355 ;
  assign n3865 = ~n2128 & ~n3864 ;
  assign n3866 = x10 & ~n513 ;
  assign n3867 = ~n3865 & n3866 ;
  assign n3868 = ~n3863 & ~n3867 ;
  assign n3869 = n1853 & ~n3868 ;
  assign n3870 = n1754 & n3408 ;
  assign n3871 = n3746 & n3870 ;
  assign n3872 = x7 & ~n3871 ;
  assign n3873 = ~n3869 & n3872 ;
  assign n3874 = ~n3861 & n3873 ;
  assign n3875 = ~x8 & n254 ;
  assign n3876 = n253 & n1104 ;
  assign n3877 = ~x4 & n3876 ;
  assign n3878 = x8 & n3877 ;
  assign n3879 = ~n3875 & ~n3878 ;
  assign n3880 = n1776 & ~n3879 ;
  assign n3881 = n1104 & n3757 ;
  assign n3882 = n2083 & n3881 ;
  assign n3883 = n2001 & n3882 ;
  assign n3884 = n1105 & n2439 ;
  assign n3885 = x12 & n3884 ;
  assign n3886 = ~n3883 & ~n3885 ;
  assign n3887 = ~n3880 & n3886 ;
  assign n3888 = n1207 & ~n3887 ;
  assign n3889 = ~x4 & n1364 ;
  assign n3890 = ~n17 & ~n3889 ;
  assign n3891 = x8 & ~n3890 ;
  assign n3892 = ~n1031 & ~n1765 ;
  assign n3893 = ~n1711 & n3892 ;
  assign n3894 = ~n1808 & ~n3406 ;
  assign n3895 = ~n1104 & n3894 ;
  assign n3896 = ~n3893 & ~n3895 ;
  assign n3897 = ~x12 & ~n2040 ;
  assign n3898 = ~n614 & n3897 ;
  assign n3899 = ~n1351 & ~n2147 ;
  assign n3900 = ~x10 & n3899 ;
  assign n3901 = ~n3898 & n3900 ;
  assign n3902 = n3896 & n3901 ;
  assign n3903 = ~n3891 & n3902 ;
  assign n3904 = x8 ^ x6 ;
  assign n3905 = n1207 & n3904 ;
  assign n3906 = x12 & n3905 ;
  assign n3907 = ~n3903 & ~n3906 ;
  assign n3908 = ~n513 & ~n3907 ;
  assign n3909 = ~x7 & ~n3908 ;
  assign n3923 = x10 & n2954 ;
  assign n3924 = n1105 & n3216 ;
  assign n3925 = ~n3923 & ~n3924 ;
  assign n3926 = n1753 & ~n3925 ;
  assign n3927 = ~x6 & n1104 ;
  assign n3928 = n3216 & n3927 ;
  assign n3929 = ~n59 & ~n3227 ;
  assign n3930 = ~n3928 & n3929 ;
  assign n3931 = n452 & ~n3930 ;
  assign n3932 = ~n3926 & ~n3931 ;
  assign n3933 = x5 & ~n3932 ;
  assign n3910 = n65 & n2954 ;
  assign n3911 = n2231 & n3910 ;
  assign n3912 = x4 & x14 ;
  assign n3913 = ~x13 & ~n3912 ;
  assign n3914 = n3791 & ~n3913 ;
  assign n3915 = n60 & n3525 ;
  assign n3916 = ~n3914 & ~n3915 ;
  assign n3917 = n3916 ^ n2128 ;
  assign n3918 = n3917 ^ n3916 ;
  assign n3919 = n3916 ^ n262 ;
  assign n3920 = ~n3918 & ~n3919 ;
  assign n3921 = n3920 ^ n3916 ;
  assign n3922 = ~n3911 & n3921 ;
  assign n3934 = n3933 ^ n3922 ;
  assign n3935 = n3934 ^ n3922 ;
  assign n3936 = n79 & n1865 ;
  assign n3937 = n1104 & n2924 ;
  assign n3938 = n3936 & n3937 ;
  assign n3939 = ~n144 & ~n3912 ;
  assign n3940 = x6 & ~n3939 ;
  assign n3941 = ~n3792 & n3940 ;
  assign n3942 = ~n3938 & ~n3941 ;
  assign n3943 = n3942 ^ n3922 ;
  assign n3944 = n3943 ^ n3922 ;
  assign n3945 = ~n3935 & n3944 ;
  assign n3946 = n3945 ^ n3922 ;
  assign n3947 = ~x0 & n3946 ;
  assign n3948 = n3947 ^ n3922 ;
  assign n3949 = ~x9 & ~n3948 ;
  assign n3950 = n1693 ^ x0 ;
  assign n3956 = n3950 ^ n1693 ;
  assign n3951 = n3950 ^ x6 ;
  assign n3952 = n3951 ^ n1693 ;
  assign n3953 = n3904 ^ x6 ;
  assign n3954 = n3953 ^ n3952 ;
  assign n3955 = ~n3952 & ~n3954 ;
  assign n3957 = n3956 ^ n3955 ;
  assign n3958 = n3957 ^ n3952 ;
  assign n3959 = n3351 ^ n1693 ;
  assign n3960 = n3955 ^ n3952 ;
  assign n3961 = n3959 & ~n3960 ;
  assign n3962 = n3961 ^ n1693 ;
  assign n3963 = ~n3958 & ~n3962 ;
  assign n3964 = n3963 ^ n1693 ;
  assign n3965 = n3964 ^ n1693 ;
  assign n3966 = n3684 & n3965 ;
  assign n3967 = x6 ^ x5 ;
  assign n3968 = n3967 ^ x5 ;
  assign n3969 = ~x10 & n1104 ;
  assign n3970 = n3969 ^ x5 ;
  assign n3971 = ~n3968 & ~n3970 ;
  assign n3972 = n3971 ^ x5 ;
  assign n3973 = n3617 & ~n3972 ;
  assign n3974 = ~n3966 & ~n3973 ;
  assign n3975 = n170 & ~n3974 ;
  assign n3976 = n3975 ^ x9 ;
  assign n3977 = n3976 ^ n3975 ;
  assign n3978 = ~x2 & ~x5 ;
  assign n3979 = n124 & n2649 ;
  assign n3980 = n992 & n3979 ;
  assign n3981 = n3978 & n3980 ;
  assign n3982 = ~n1753 & ~n2001 ;
  assign n3983 = n1831 & ~n3982 ;
  assign n3984 = ~n2974 & n3983 ;
  assign n3985 = ~n137 & n3399 ;
  assign n3986 = n2128 & n3985 ;
  assign n3987 = ~n3984 & ~n3986 ;
  assign n3988 = n261 & ~n3987 ;
  assign n3989 = n1104 & n2062 ;
  assign n3990 = n23 & n1765 ;
  assign n3991 = n3989 & n3990 ;
  assign n3992 = ~n3988 & ~n3991 ;
  assign n3993 = ~n3981 & n3992 ;
  assign n3994 = n3993 ^ n3975 ;
  assign n3995 = n3994 ^ n3975 ;
  assign n3996 = n3977 & ~n3995 ;
  assign n3997 = n3996 ^ n3975 ;
  assign n3998 = x4 & n3997 ;
  assign n3999 = n3998 ^ n3975 ;
  assign n4000 = ~n3949 & ~n3999 ;
  assign n4001 = n3909 & n4000 ;
  assign n4002 = ~n3888 & n4001 ;
  assign n4003 = ~n3874 & ~n4002 ;
  assign n4004 = n1754 & n3802 ;
  assign n4005 = ~x5 & ~n2704 ;
  assign n4006 = n2974 & n4005 ;
  assign n4007 = n1356 & n2827 ;
  assign n4008 = ~n4006 & ~n4007 ;
  assign n4009 = n1305 & ~n4008 ;
  assign n4010 = ~x0 & n4009 ;
  assign n4011 = ~n4004 & ~n4010 ;
  assign n4012 = n2298 & ~n4011 ;
  assign n4013 = n1355 & n2953 ;
  assign n4014 = ~n3990 & ~n4013 ;
  assign n4015 = x4 & n1853 ;
  assign n4016 = ~n4014 & n4015 ;
  assign n4017 = n1711 & n2945 ;
  assign n4018 = n434 & n4017 ;
  assign n4019 = n992 & n4018 ;
  assign n4020 = ~n4016 & ~n4019 ;
  assign n4021 = ~n513 & ~n4020 ;
  assign n4022 = ~n4012 & ~n4021 ;
  assign n4023 = ~n4003 & n4022 ;
  assign n4024 = x3 & n4023 ;
  assign n4025 = ~x6 & n205 ;
  assign n4026 = ~n170 & ~n525 ;
  assign n4027 = n4025 & ~n4026 ;
  assign n4028 = ~x6 & n1853 ;
  assign n4029 = ~n1031 & n2035 ;
  assign n4030 = ~n1314 & n4029 ;
  assign n4031 = ~n2704 & n4030 ;
  assign n4032 = ~n4028 & ~n4031 ;
  assign n4033 = x5 & ~n4032 ;
  assign n4034 = n1031 & n1696 ;
  assign n4035 = x8 & ~n3744 ;
  assign n4036 = ~n525 & n1765 ;
  assign n4037 = ~n4035 & n4036 ;
  assign n4038 = ~n4034 & ~n4037 ;
  assign n4039 = ~n4033 & n4038 ;
  assign n4040 = ~x10 & ~n4039 ;
  assign n4041 = ~n4027 & ~n4040 ;
  assign n4042 = n1872 & ~n4041 ;
  assign n4043 = ~x5 & n17 ;
  assign n4044 = ~x10 & n525 ;
  assign n4045 = ~n3143 & ~n4044 ;
  assign n4046 = n4043 & ~n4045 ;
  assign n4047 = n658 & n2833 ;
  assign n4048 = ~n4046 & ~n4047 ;
  assign n4049 = n1315 & ~n4048 ;
  assign n4050 = n1336 & ~n2706 ;
  assign n4051 = ~n59 & ~n4050 ;
  assign n4052 = n2954 & ~n4051 ;
  assign n4053 = n2147 & n4052 ;
  assign n4054 = n432 & ~n1104 ;
  assign n4055 = n1355 & n3406 ;
  assign n4056 = ~n4054 & n4055 ;
  assign n4057 = ~n1632 & ~n3744 ;
  assign n4058 = n3085 & ~n4057 ;
  assign n4059 = ~x5 & ~x10 ;
  assign n4060 = n3227 & n4059 ;
  assign n4061 = x14 & n1042 ;
  assign n4062 = ~n1364 & ~n4061 ;
  assign n4063 = n1731 & ~n4062 ;
  assign n4064 = ~n4060 & ~n4063 ;
  assign n4065 = ~n4058 & n4064 ;
  assign n4066 = n2945 & ~n4065 ;
  assign n4067 = ~n4056 & ~n4066 ;
  assign n4068 = ~n4053 & n4067 ;
  assign n4069 = n4068 ^ x7 ;
  assign n4070 = n4069 ^ n4068 ;
  assign n4071 = n4070 ^ n4049 ;
  assign n4072 = n335 & n992 ;
  assign n4073 = n812 & n2924 ;
  assign n4074 = n4072 & n4073 ;
  assign n4075 = n812 & ~n1106 ;
  assign n4076 = n2147 ^ n281 ;
  assign n4077 = n4076 ^ n2147 ;
  assign n4078 = n1104 & n2128 ;
  assign n4079 = n4078 ^ n2147 ;
  assign n4080 = ~n4077 & n4079 ;
  assign n4081 = n4080 ^ n2147 ;
  assign n4082 = x9 & n4081 ;
  assign n4083 = ~n4075 & ~n4082 ;
  assign n4084 = x12 & ~n4083 ;
  assign n4085 = ~n4074 & ~n4084 ;
  assign n4086 = n4085 ^ x4 ;
  assign n4087 = ~n4085 & n4086 ;
  assign n4088 = n4087 ^ n4068 ;
  assign n4089 = n4088 ^ n4085 ;
  assign n4090 = ~n4071 & n4089 ;
  assign n4091 = n4090 ^ n4087 ;
  assign n4092 = n4091 ^ n4085 ;
  assign n4093 = ~n4049 & ~n4092 ;
  assign n4094 = n4093 ^ n4049 ;
  assign n4095 = ~n4042 & ~n4094 ;
  assign n4096 = ~n513 & ~n4095 ;
  assign n4097 = n4096 ^ x3 ;
  assign n4098 = n170 & n4017 ;
  assign n4099 = n3406 & n4013 ;
  assign n4100 = ~n4098 & ~n4099 ;
  assign n4101 = n1104 & ~n4100 ;
  assign n4102 = ~n167 & ~n1632 ;
  assign n4103 = n2945 & ~n4102 ;
  assign n4104 = ~n144 & n518 ;
  assign n4105 = ~n137 & n4104 ;
  assign n4106 = ~n2691 & ~n4105 ;
  assign n4107 = ~n1765 & ~n3088 ;
  assign n4108 = ~n4106 & ~n4107 ;
  assign n4109 = ~n167 & n4108 ;
  assign n4110 = ~n4103 & ~n4109 ;
  assign n4111 = n3406 & ~n4110 ;
  assign n4112 = n529 & n1718 ;
  assign n4113 = n3848 & n4112 ;
  assign n4114 = n231 & n4113 ;
  assign n4115 = ~n4111 & ~n4114 ;
  assign n4116 = ~n4101 & n4115 ;
  assign n4117 = n499 & ~n4116 ;
  assign n4118 = ~n432 & n1355 ;
  assign n4119 = ~x6 & n2691 ;
  assign n4120 = ~n4118 & ~n4119 ;
  assign n4121 = n254 & ~n4120 ;
  assign n4122 = n174 & n2035 ;
  assign n4123 = n4102 & n4122 ;
  assign n4124 = n3490 ^ x9 ;
  assign n4125 = n601 ^ x9 ;
  assign n4126 = ~n4124 & n4125 ;
  assign n4127 = n4126 ^ x9 ;
  assign n4128 = n205 & n4127 ;
  assign n4129 = ~n572 & n4128 ;
  assign n4130 = ~n4123 & ~n4129 ;
  assign n4131 = n992 & ~n4130 ;
  assign n4132 = ~x5 & x14 ;
  assign n4133 = n1753 & n4132 ;
  assign n4134 = ~n167 & n4133 ;
  assign n4135 = n1597 & n4134 ;
  assign n4136 = ~n4131 & ~n4135 ;
  assign n4137 = ~n4121 & n4136 ;
  assign n4138 = n2083 & ~n4137 ;
  assign n4139 = n3243 & n3621 ;
  assign n4140 = ~n4138 & ~n4139 ;
  assign n4141 = ~n4117 & n4140 ;
  assign n4142 = n4141 ^ x7 ;
  assign n4143 = n4142 ^ n4141 ;
  assign n4144 = ~x4 & n265 ;
  assign n4145 = n812 & n988 ;
  assign n4146 = ~n1699 & n4145 ;
  assign n4147 = n4144 & n4146 ;
  assign n4148 = n79 & n1132 ;
  assign n4149 = n2243 & n4148 ;
  assign n4150 = n539 & ~n3483 ;
  assign n4151 = ~n3848 & n4150 ;
  assign n4152 = ~n281 & ~n1132 ;
  assign n4153 = n2128 & ~n4152 ;
  assign n4154 = ~n3848 & ~n4078 ;
  assign n4155 = n432 & ~n4154 ;
  assign n4156 = ~n4153 & ~n4155 ;
  assign n4157 = ~n4151 & n4156 ;
  assign n4158 = n2298 & ~n4157 ;
  assign n4159 = ~n4149 & ~n4158 ;
  assign n4160 = ~n4147 & n4159 ;
  assign n4161 = n920 & ~n4160 ;
  assign n4162 = n1197 & n1711 ;
  assign n4163 = n2996 & n4162 ;
  assign n4164 = n3848 & n4145 ;
  assign n4165 = ~n4075 & ~n4164 ;
  assign n4166 = x4 & ~n4165 ;
  assign n4167 = n432 & n1104 ;
  assign n4168 = n4152 & ~n4167 ;
  assign n4169 = n4043 & ~n4168 ;
  assign n4170 = ~n4166 & ~n4169 ;
  assign n4171 = ~n4163 & n4170 ;
  assign n4172 = n2130 & ~n4171 ;
  assign n4173 = n2823 & n3778 ;
  assign n4174 = n3626 & n4173 ;
  assign n4175 = n3791 & n4174 ;
  assign n4176 = x5 & n4175 ;
  assign n4177 = ~n4172 & ~n4176 ;
  assign n4178 = ~n4161 & n4177 ;
  assign n4179 = n4178 ^ n4141 ;
  assign n4180 = n4143 & n4179 ;
  assign n4181 = n4180 ^ n4141 ;
  assign n4182 = n4181 ^ n4096 ;
  assign n4183 = n4097 & ~n4182 ;
  assign n4184 = n4183 ^ n4180 ;
  assign n4185 = n4184 ^ n4141 ;
  assign n4186 = n4185 ^ x3 ;
  assign n4187 = ~n4096 & ~n4186 ;
  assign n4188 = n4187 ^ n4096 ;
  assign n4189 = ~n4024 & n4188 ;
  assign n4190 = n2869 & n3746 ;
  assign n4191 = n190 & n1853 ;
  assign n4192 = n1101 & n3616 ;
  assign n4193 = ~n4191 & ~n4192 ;
  assign n4194 = n2242 & ~n4193 ;
  assign n4195 = ~x9 & n1104 ;
  assign n4196 = n125 & n4144 ;
  assign n4197 = n4195 & n4196 ;
  assign n4198 = ~n4194 & ~n4197 ;
  assign n4199 = ~n4190 & n4198 ;
  assign n4200 = n2974 & ~n4199 ;
  assign n4201 = ~n513 & n4200 ;
  assign n4202 = n60 & n1207 ;
  assign n4203 = n3639 & n3969 ;
  assign n4204 = ~n4202 & ~n4203 ;
  assign n4205 = n2083 & ~n4204 ;
  assign n4206 = n2242 & n3969 ;
  assign n4207 = n3617 & n4206 ;
  assign n4208 = ~n4205 & ~n4207 ;
  assign n4209 = n2827 & ~n4208 ;
  assign n4210 = n499 & n1718 ;
  assign n4211 = n124 & n1696 ;
  assign n4212 = n4210 & n4211 ;
  assign n4213 = n1132 & n1759 ;
  assign n4214 = n1104 & n2818 ;
  assign n4215 = n1705 & n4214 ;
  assign n4216 = n4213 & n4215 ;
  assign n4217 = ~n4212 & ~n4216 ;
  assign n4218 = ~n4209 & n4217 ;
  assign n4219 = n1527 & ~n4218 ;
  assign n4220 = ~x4 & n3862 ;
  assign n4221 = n1315 & n4220 ;
  assign n4222 = n2696 & n4221 ;
  assign n4223 = ~n4219 & ~n4222 ;
  assign n4224 = ~n4201 & n4223 ;
  assign n4225 = ~n4189 & n4224 ;
  assign n4226 = ~n3717 & n4225 ;
  assign n4227 = n2269 & ~n4226 ;
  assign n4228 = ~n2113 & ~n2298 ;
  assign n4229 = ~x1 & x8 ;
  assign n4230 = n141 & n3365 ;
  assign n4231 = n362 & n2579 ;
  assign n4232 = ~n4230 & ~n4231 ;
  assign n4233 = n100 & n432 ;
  assign n4234 = n65 & ~n606 ;
  assign n4235 = ~n4233 & ~n4234 ;
  assign n4236 = n4235 ^ x2 ;
  assign n4237 = n4236 ^ n4235 ;
  assign n4238 = n4235 ^ n1567 ;
  assign n4239 = n4238 ^ n4235 ;
  assign n4240 = ~n4237 & n4239 ;
  assign n4241 = n4240 ^ n4235 ;
  assign n4242 = x0 & ~n4241 ;
  assign n4243 = n4242 ^ n4235 ;
  assign n4244 = ~n4232 & ~n4243 ;
  assign n4245 = ~n2706 & n2720 ;
  assign n4246 = ~n1765 & ~n3483 ;
  assign n4247 = ~x3 & n4246 ;
  assign n4248 = n4245 & n4247 ;
  assign n4249 = n537 & n2128 ;
  assign n4250 = n1995 & n4249 ;
  assign n4251 = ~n4248 & ~n4250 ;
  assign n4252 = n99 & ~n4251 ;
  assign n4253 = ~n4244 & ~n4252 ;
  assign n4254 = x14 & ~n4253 ;
  assign n4255 = n141 & n658 ;
  assign n4256 = n499 & n755 ;
  assign n4257 = n4255 & n4256 ;
  assign n4258 = ~n4254 & ~n4257 ;
  assign n4259 = n4229 & ~n4258 ;
  assign n4260 = ~x2 & ~n1198 ;
  assign n4261 = n152 & n2309 ;
  assign n4262 = x9 & n4261 ;
  assign n4263 = n604 & n1766 ;
  assign n4264 = n191 & n4263 ;
  assign n4265 = n1831 & n3229 ;
  assign n4266 = ~n616 & n629 ;
  assign n4267 = n4265 & n4266 ;
  assign n4268 = ~n4264 & ~n4267 ;
  assign n4269 = ~n4262 & n4268 ;
  assign n4270 = n4260 & ~n4269 ;
  assign n4271 = ~x10 & n1579 ;
  assign n4272 = n743 & n4271 ;
  assign n4273 = n218 & n1765 ;
  assign n4274 = ~n1198 & n4273 ;
  assign n4275 = n4272 & n4274 ;
  assign n4276 = n792 & n3428 ;
  assign n4277 = ~x13 & n1579 ;
  assign n4278 = ~x5 & n25 ;
  assign n4279 = n4277 & n4278 ;
  assign n4280 = ~n4276 & ~n4279 ;
  assign n4281 = n19 & n2974 ;
  assign n4282 = ~n4280 & n4281 ;
  assign n4283 = ~x2 & n4282 ;
  assign n4284 = ~n4275 & ~n4283 ;
  assign n4285 = ~n4270 & n4284 ;
  assign n4286 = x1 & ~n4285 ;
  assign n4290 = n182 & n1914 ;
  assign n4287 = ~n606 & n624 ;
  assign n4288 = x0 & n1567 ;
  assign n4289 = ~n4287 & ~n4288 ;
  assign n4291 = n4290 ^ n4289 ;
  assign n4292 = n130 & n2147 ;
  assign n4293 = n4292 ^ n4291 ;
  assign n4294 = n4293 ^ n4289 ;
  assign n4295 = n4294 ^ n4293 ;
  assign n4296 = ~n2133 & ~n2333 ;
  assign n4297 = n624 & ~n4296 ;
  assign n4298 = n471 & n1704 ;
  assign n4299 = n4298 ^ x10 ;
  assign n4300 = n4299 ^ n4298 ;
  assign n4301 = n4300 ^ n4297 ;
  assign n4302 = n846 ^ n604 ;
  assign n4303 = n604 & n4302 ;
  assign n4304 = n4303 ^ n4298 ;
  assign n4305 = n4304 ^ n604 ;
  assign n4306 = n4301 & n4305 ;
  assign n4307 = n4306 ^ n4303 ;
  assign n4308 = n4307 ^ n604 ;
  assign n4309 = ~n4297 & n4308 ;
  assign n4310 = n4309 ^ n4297 ;
  assign n4311 = n4310 ^ n4293 ;
  assign n4312 = n4311 ^ n4291 ;
  assign n4313 = ~n4295 & ~n4312 ;
  assign n4314 = n4313 ^ n4310 ;
  assign n4315 = ~n396 & ~n4310 ;
  assign n4316 = n4315 ^ n4291 ;
  assign n4317 = ~n4314 & n4316 ;
  assign n4318 = n4317 ^ n4315 ;
  assign n4319 = n4291 & n4318 ;
  assign n4320 = n4319 ^ n4313 ;
  assign n4321 = n4320 ^ n4290 ;
  assign n4322 = n4321 ^ n4310 ;
  assign n4323 = ~n526 & ~n4322 ;
  assign n4324 = ~n4286 & ~n4323 ;
  assign n4325 = n4324 ^ x8 ;
  assign n4326 = n4325 ^ n4324 ;
  assign n4327 = n128 & n4265 ;
  assign n4328 = n142 & n2307 ;
  assign n4329 = x2 & n4328 ;
  assign n4330 = ~n534 & n4329 ;
  assign n4331 = ~n4327 & ~n4330 ;
  assign n4332 = ~n167 & ~n920 ;
  assign n4333 = ~n606 & ~n1198 ;
  assign n4334 = ~n4332 & n4333 ;
  assign n4335 = ~n4331 & n4334 ;
  assign n4336 = ~n1054 & ~n3851 ;
  assign n4337 = n4230 & n4336 ;
  assign n4338 = n2128 & n2299 ;
  assign n4339 = n191 & n4338 ;
  assign n4340 = ~n4337 & ~n4339 ;
  assign n4341 = n605 & ~n4340 ;
  assign n4342 = ~x3 & n801 ;
  assign n4343 = n2649 & n4342 ;
  assign n4344 = n4233 & n4343 ;
  assign n4345 = ~n4341 & ~n4344 ;
  assign n4346 = n4345 ^ x14 ;
  assign n4347 = n4345 ^ x13 ;
  assign n4348 = n4347 ^ x13 ;
  assign n4349 = ~x3 & n197 ;
  assign n4350 = n3488 & n4349 ;
  assign n4351 = n2447 & n3482 ;
  assign n4352 = ~n4350 & ~n4351 ;
  assign n4353 = n624 & ~n4352 ;
  assign n4354 = ~x5 & n3068 ;
  assign n4355 = ~n2456 & n4354 ;
  assign n4356 = n562 & n855 ;
  assign n4357 = ~n4355 & ~n4356 ;
  assign n4358 = n3408 & ~n4357 ;
  assign n4359 = ~n4353 & ~n4358 ;
  assign n4360 = n2001 & ~n4359 ;
  assign n4361 = n1586 & n2308 ;
  assign n4362 = x0 & ~n1704 ;
  assign n4363 = n142 ^ n141 ;
  assign n4364 = n4363 ^ n4362 ;
  assign n4365 = n141 ^ x13 ;
  assign n4366 = n141 ^ x11 ;
  assign n4367 = n4366 ^ n4365 ;
  assign n4368 = n4365 & n4367 ;
  assign n4369 = n4368 ^ n141 ;
  assign n4370 = n4369 ^ n4365 ;
  assign n4371 = n4364 & n4370 ;
  assign n4372 = n4371 ^ n4368 ;
  assign n4373 = n4372 ^ n4365 ;
  assign n4374 = n4362 & n4373 ;
  assign n4375 = ~n4361 & ~n4374 ;
  assign n4376 = n3840 & ~n4375 ;
  assign n4378 = n142 & n3193 ;
  assign n4377 = n1944 ^ x0 ;
  assign n4379 = n4378 ^ n4377 ;
  assign n4380 = n4379 ^ n1944 ;
  assign n4386 = n4380 ^ n4377 ;
  assign n4387 = n4386 ^ n1944 ;
  assign n4388 = n4387 ^ n1944 ;
  assign n4389 = ~n606 & n4342 ;
  assign n4390 = n4389 ^ n4377 ;
  assign n4391 = n4390 ^ n4377 ;
  assign n4392 = n4391 ^ n1944 ;
  assign n4393 = n4388 & n4392 ;
  assign n4381 = n799 & n4349 ;
  assign n4382 = n4381 ^ n4377 ;
  assign n4383 = n4382 ^ n4380 ;
  assign n4384 = n4383 ^ n1944 ;
  assign n4385 = n4380 & n4384 ;
  assign n4394 = n4393 ^ n4385 ;
  assign n4395 = n4394 ^ n4380 ;
  assign n4396 = n4385 ^ n1944 ;
  assign n4397 = n4396 ^ n4387 ;
  assign n4398 = ~n1944 & n4397 ;
  assign n4399 = n4398 ^ n4385 ;
  assign n4400 = n4395 & n4399 ;
  assign n4401 = n4400 ^ n4393 ;
  assign n4402 = n4401 ^ n4398 ;
  assign n4403 = n4402 ^ n4380 ;
  assign n4404 = n4403 ^ n1944 ;
  assign n4405 = n4404 ^ n4387 ;
  assign n4406 = n4405 ^ x0 ;
  assign n4407 = n2974 & n4406 ;
  assign n4408 = x2 & n4407 ;
  assign n4409 = ~n4376 & ~n4408 ;
  assign n4410 = ~n4360 & n4409 ;
  assign n4411 = n4410 ^ x13 ;
  assign n4412 = n4348 & n4411 ;
  assign n4413 = n4412 ^ x13 ;
  assign n4414 = ~n4346 & n4413 ;
  assign n4415 = n4414 ^ x14 ;
  assign n4416 = ~n4335 & ~n4415 ;
  assign n4417 = x1 & ~n4416 ;
  assign n4418 = x14 & n540 ;
  assign n4419 = ~x3 & n2231 ;
  assign n4420 = n306 & n4419 ;
  assign n4421 = ~x7 & n4420 ;
  assign n4422 = n754 & n1732 ;
  assign n4423 = n830 & n1729 ;
  assign n4424 = ~n4422 & ~n4423 ;
  assign n4425 = n4354 & ~n4424 ;
  assign n4426 = n3365 & n4349 ;
  assign n4427 = ~n137 & n4426 ;
  assign n4428 = ~n4425 & ~n4427 ;
  assign n4429 = x9 & ~n4428 ;
  assign n4430 = ~n4421 & ~n4429 ;
  assign n4433 = n4430 ^ x3 ;
  assign n4434 = n4433 ^ n4430 ;
  assign n4431 = n4430 ^ n1847 ;
  assign n4432 = n4431 ^ n4430 ;
  assign n4435 = n4434 ^ n4432 ;
  assign n4436 = ~x9 & n305 ;
  assign n4437 = n286 & n4436 ;
  assign n4438 = n4437 ^ n4430 ;
  assign n4439 = n4438 ^ n4430 ;
  assign n4440 = n4439 ^ n4434 ;
  assign n4441 = ~n4434 & ~n4440 ;
  assign n4442 = n4441 ^ n4434 ;
  assign n4443 = ~n4435 & ~n4442 ;
  assign n4444 = n4443 ^ n4441 ;
  assign n4445 = n4444 ^ n4430 ;
  assign n4446 = n4445 ^ n4434 ;
  assign n4447 = ~x2 & n4446 ;
  assign n4448 = n4447 ^ n4430 ;
  assign n4449 = n4418 & ~n4448 ;
  assign n4450 = n4449 ^ n470 ;
  assign n4452 = x10 ^ x6 ;
  assign n4451 = n4354 ^ n4230 ;
  assign n4453 = n4452 ^ n4451 ;
  assign n4458 = n4453 ^ n4451 ;
  assign n4454 = n4453 ^ n4354 ;
  assign n4455 = n4454 ^ x13 ;
  assign n4456 = n4455 ^ x10 ;
  assign n4457 = n4456 ^ n4451 ;
  assign n4459 = n4458 ^ n4457 ;
  assign n4461 = n4456 ^ x10 ;
  assign n4460 = n4457 ^ n221 ;
  assign n4462 = n4461 ^ n4460 ;
  assign n4463 = n4459 & n4462 ;
  assign n4464 = n4463 ^ n4456 ;
  assign n4465 = n4464 ^ n221 ;
  assign n4466 = n4465 ^ n4461 ;
  assign n4467 = n4460 ^ n4458 ;
  assign n4468 = ~n4464 & ~n4467 ;
  assign n4469 = n4468 ^ n4456 ;
  assign n4470 = n4469 ^ n4457 ;
  assign n4471 = n4470 ^ n4458 ;
  assign n4472 = n4466 & ~n4471 ;
  assign n4473 = n4472 ^ n4230 ;
  assign n4474 = x9 & n4473 ;
  assign n4475 = ~n4420 & ~n4474 ;
  assign n4476 = n1255 & ~n4475 ;
  assign n4477 = n432 & n4342 ;
  assign n4478 = n843 & n2579 ;
  assign n4479 = ~n4477 & ~n4478 ;
  assign n4480 = x2 & ~n4479 ;
  assign n4481 = ~n526 & n4480 ;
  assign n4482 = ~n4476 & ~n4481 ;
  assign n4483 = n4482 ^ x7 ;
  assign n4484 = n4483 ^ n4482 ;
  assign n4485 = n1696 & n3466 ;
  assign n4486 = n1439 & n4485 ;
  assign n4487 = n859 & n2128 ;
  assign n4488 = n65 & n978 ;
  assign n4489 = n4487 & n4488 ;
  assign n4490 = ~x11 & ~n1198 ;
  assign n4491 = n4419 & n4490 ;
  assign n4492 = n4491 ^ n1104 ;
  assign n4493 = n4492 ^ n4491 ;
  assign n4494 = n4491 ^ n4328 ;
  assign n4495 = n4494 ^ n4491 ;
  assign n4496 = n4493 & n4495 ;
  assign n4497 = n4496 ^ n4491 ;
  assign n4498 = ~x2 & n4497 ;
  assign n4499 = n4498 ^ n4491 ;
  assign n4500 = n642 & n4499 ;
  assign n4501 = ~n4489 & ~n4500 ;
  assign n4502 = ~n4486 & n4501 ;
  assign n4503 = n4502 ^ n4482 ;
  assign n4504 = n4484 & n4503 ;
  assign n4505 = n4504 ^ n4482 ;
  assign n4506 = n4505 ^ n4449 ;
  assign n4507 = ~n4450 & n4506 ;
  assign n4508 = n4507 ^ n4504 ;
  assign n4509 = n4508 ^ n4482 ;
  assign n4510 = n4509 ^ n470 ;
  assign n4511 = ~n4449 & ~n4510 ;
  assign n4512 = n4511 ^ n4449 ;
  assign n4513 = n4512 ^ n4449 ;
  assign n4514 = ~n4417 & n4513 ;
  assign n4515 = n4514 ^ n4324 ;
  assign n4516 = ~n4326 & n4515 ;
  assign n4517 = n4516 ^ n4324 ;
  assign n4518 = ~n4259 & n4517 ;
  assign n4519 = ~n4228 & ~n4518 ;
  assign n4520 = x4 & n1766 ;
  assign n4521 = n262 & n4520 ;
  assign n4522 = n106 & n1718 ;
  assign n4523 = n124 & n1712 ;
  assign n4524 = n4522 & n4523 ;
  assign n4525 = n141 & n1865 ;
  assign n4526 = n236 & n3848 ;
  assign n4527 = n4525 & n4526 ;
  assign n4528 = ~n4524 & ~n4527 ;
  assign n4529 = x0 & ~n4528 ;
  assign n4530 = ~n4521 & ~n4529 ;
  assign n4531 = x13 & ~n4530 ;
  assign n4532 = n1042 & n1788 ;
  assign n4533 = n442 & n2945 ;
  assign n4534 = n4532 & n4533 ;
  assign n4535 = n236 & n2147 ;
  assign n4536 = n1165 & n2035 ;
  assign n4537 = ~n4535 & ~n4536 ;
  assign n4538 = n1705 & ~n4537 ;
  assign n4539 = ~x6 & n1865 ;
  assign n4540 = x12 ^ x5 ;
  assign n4541 = n830 ^ n754 ;
  assign n4542 = n830 ^ x12 ;
  assign n4543 = n4542 ^ n830 ;
  assign n4544 = n4541 & ~n4543 ;
  assign n4545 = n4544 ^ n830 ;
  assign n4546 = ~n4540 & n4545 ;
  assign n4547 = n4546 ^ x3 ;
  assign n4548 = n4547 ^ n4546 ;
  assign n4549 = n249 & n754 ;
  assign n4550 = n4549 ^ n4546 ;
  assign n4551 = ~n4548 & n4550 ;
  assign n4552 = n4551 ^ n4546 ;
  assign n4553 = n4539 & n4552 ;
  assign n4554 = ~n4538 & ~n4553 ;
  assign n4555 = n2685 & ~n4554 ;
  assign n4556 = ~x13 & n142 ;
  assign n4557 = n2834 & n4556 ;
  assign n4558 = n1150 & n2833 ;
  assign n4559 = n2095 & n2954 ;
  assign n4560 = n1207 & n4559 ;
  assign n4561 = ~n4558 & ~n4560 ;
  assign n4562 = ~n4557 & n4561 ;
  assign n4563 = x12 & ~n4562 ;
  assign n4564 = n137 & n265 ;
  assign n4565 = n2381 & n4564 ;
  assign n4566 = ~n4563 & ~n4565 ;
  assign n4567 = n442 & ~n4566 ;
  assign n4568 = x13 ^ x0 ;
  assign n4569 = n4524 ^ x13 ;
  assign n4570 = n4569 ^ n4524 ;
  assign n4571 = n4570 ^ n4568 ;
  assign n4572 = ~x6 & n207 ;
  assign n4573 = n108 & ~n2148 ;
  assign n4574 = ~x10 & n4573 ;
  assign n4575 = ~n4572 & ~n4574 ;
  assign n4576 = n4575 ^ n4144 ;
  assign n4577 = n4144 & ~n4576 ;
  assign n4578 = n4577 ^ n4524 ;
  assign n4579 = n4578 ^ n4144 ;
  assign n4580 = ~n4571 & n4579 ;
  assign n4581 = n4580 ^ n4577 ;
  assign n4582 = n4581 ^ n4144 ;
  assign n4583 = n4568 & n4582 ;
  assign n4584 = ~n4567 & ~n4583 ;
  assign n4585 = ~n4555 & n4584 ;
  assign n4586 = x14 & ~n4585 ;
  assign n4587 = ~n4534 & ~n4586 ;
  assign n4588 = ~n4531 & n4587 ;
  assign n4589 = x11 ^ x9 ;
  assign n4590 = n112 ^ n48 ;
  assign n4591 = n112 ^ x11 ;
  assign n4592 = n4591 ^ n112 ;
  assign n4593 = n4590 & ~n4592 ;
  assign n4594 = n4593 ^ n112 ;
  assign n4595 = n4589 & n4594 ;
  assign n4596 = ~n4588 & n4595 ;
  assign n4597 = ~x7 & n1718 ;
  assign n4598 = n3296 & n4597 ;
  assign n4599 = n191 & n286 ;
  assign n4600 = n2298 & n4599 ;
  assign n4601 = ~n4598 & ~n4600 ;
  assign n4602 = n3626 & ~n4601 ;
  assign n4603 = ~x4 & n1831 ;
  assign n4604 = n329 & n4603 ;
  assign n4605 = n604 & n4604 ;
  assign n4606 = n125 & n3234 ;
  assign n4607 = n4271 & n4606 ;
  assign n4608 = x10 & n2652 ;
  assign n4609 = n1759 & n4608 ;
  assign n4610 = ~n799 & ~n1586 ;
  assign n4611 = n4609 & ~n4610 ;
  assign n4612 = ~n4607 & ~n4611 ;
  assign n4613 = ~n4605 & n4612 ;
  assign n4614 = n992 & ~n4613 ;
  assign n4615 = ~n4602 & ~n4614 ;
  assign n4616 = n2945 & ~n4615 ;
  assign n4617 = n556 & n3085 ;
  assign n4618 = n152 & n1711 ;
  assign n4619 = ~n4617 & ~n4618 ;
  assign n4620 = x0 & n20 ;
  assign n4621 = ~n4619 & n4620 ;
  assign n4622 = n709 & n1718 ;
  assign n4623 = n890 & n4622 ;
  assign n4624 = ~n4621 & ~n4623 ;
  assign n4625 = n3757 & n3778 ;
  assign n4626 = ~n4624 & n4625 ;
  assign n4627 = ~x11 & n992 ;
  assign n4628 = n890 & n3808 ;
  assign n4629 = n4627 & n4628 ;
  assign n4630 = ~x7 & n167 ;
  assign n4631 = ~x8 & ~n4630 ;
  assign n4632 = n4631 ^ x0 ;
  assign n4633 = n4632 ^ n4631 ;
  assign n4634 = n4633 ^ n4629 ;
  assign n4635 = n979 & n3808 ;
  assign n4636 = ~n960 & ~n4635 ;
  assign n4637 = n4636 ^ x7 ;
  assign n4638 = ~n4636 & n4637 ;
  assign n4639 = n4638 ^ n4631 ;
  assign n4640 = n4639 ^ n4636 ;
  assign n4641 = n4634 & n4640 ;
  assign n4642 = n4641 ^ n4638 ;
  assign n4643 = n4642 ^ n4636 ;
  assign n4644 = ~n4629 & ~n4643 ;
  assign n4645 = n4644 ^ n4629 ;
  assign n4646 = n4043 & n4645 ;
  assign n4647 = ~x10 & ~n1376 ;
  assign n4648 = n3212 & n4213 ;
  assign n4649 = ~n4647 & n4648 ;
  assign n4650 = ~n4646 & ~n4649 ;
  assign n4651 = ~n4626 & n4650 ;
  assign n4652 = ~n4616 & n4651 ;
  assign n4653 = n218 & ~n4652 ;
  assign n4676 = n2368 & n3423 ;
  assign n4677 = n1197 & n3143 ;
  assign n4678 = n4676 & n4677 ;
  assign n4679 = x14 & n108 ;
  assign n4680 = n2945 & n4679 ;
  assign n4681 = ~x8 & n1817 ;
  assign n4682 = n4260 & n4681 ;
  assign n4683 = ~n4680 & ~n4682 ;
  assign n4684 = n34 & n2977 ;
  assign n4685 = ~n4683 & n4684 ;
  assign n4686 = ~n4678 & ~n4685 ;
  assign n4687 = ~x4 & ~n4686 ;
  assign n4688 = ~n518 & ~n601 ;
  assign n4689 = n3012 & ~n4688 ;
  assign n4690 = n2977 & n4689 ;
  assign n4691 = n333 & n4690 ;
  assign n4692 = ~n4687 & ~n4691 ;
  assign n4654 = x1 & ~n2128 ;
  assign n4655 = ~n4539 & n4654 ;
  assign n4656 = ~n34 & ~n48 ;
  assign n4657 = ~n2635 & n4656 ;
  assign n4658 = ~n4655 & ~n4657 ;
  assign n4659 = ~n52 & ~n1197 ;
  assign n4660 = ~n98 & ~n518 ;
  assign n4661 = ~n4659 & ~n4660 ;
  assign n4662 = ~n639 & ~n2355 ;
  assign n4663 = n4661 & ~n4662 ;
  assign n4664 = n4658 & n4663 ;
  assign n4665 = n1117 & n3927 ;
  assign n4666 = n1865 & n4665 ;
  assign n4667 = ~x1 & n4666 ;
  assign n4668 = ~n4664 & ~n4667 ;
  assign n4669 = n1579 & ~n4668 ;
  assign n4670 = x13 & n801 ;
  assign n4671 = n498 & n604 ;
  assign n4672 = n3155 & n4671 ;
  assign n4673 = n87 & n4672 ;
  assign n4674 = n4670 & n4673 ;
  assign n4675 = ~n4669 & ~n4674 ;
  assign n4693 = n4692 ^ n4675 ;
  assign n4694 = n4693 ^ n4675 ;
  assign n4695 = ~x6 & x7 ;
  assign n4696 = n2580 & n4695 ;
  assign n4697 = n83 & n87 ;
  assign n4698 = n4696 & n4697 ;
  assign n4699 = n1862 & n4278 ;
  assign n4700 = n1667 & n4699 ;
  assign n4701 = ~n4698 & ~n4700 ;
  assign n4702 = ~n526 & ~n4701 ;
  assign n4703 = n4702 ^ n4675 ;
  assign n4704 = n4703 ^ n4675 ;
  assign n4705 = n4694 & ~n4704 ;
  assign n4706 = n4705 ^ n4675 ;
  assign n4707 = x0 & n4706 ;
  assign n4708 = n4707 ^ n4675 ;
  assign n4709 = ~n81 & ~n4708 ;
  assign n4710 = ~n4653 & ~n4709 ;
  assign n4711 = x0 & ~n526 ;
  assign n4712 = ~n1197 & ~n4711 ;
  assign n4713 = ~x7 & n170 ;
  assign n4714 = n2580 & n4713 ;
  assign n4715 = n1351 & n3560 ;
  assign n4716 = n1872 & n4715 ;
  assign n4717 = ~n4714 & ~n4716 ;
  assign n4718 = n60 & n2953 ;
  assign n4719 = n129 & n4718 ;
  assign n4720 = n452 & n1896 ;
  assign n4721 = n343 & n4720 ;
  assign n4722 = ~n4719 & ~n4721 ;
  assign n4723 = ~n4717 & ~n4722 ;
  assign n4724 = ~n4712 & n4723 ;
  assign n4725 = n59 & n190 ;
  assign n4726 = n230 & n1197 ;
  assign n4727 = n2412 & n4726 ;
  assign n4728 = ~n4725 & ~n4727 ;
  assign n4729 = n3285 & ~n4728 ;
  assign n4730 = n1031 & n2818 ;
  assign n4731 = n3154 & n4730 ;
  assign n4732 = n627 & n4731 ;
  assign n4733 = n941 & n3778 ;
  assign n4734 = ~x4 & n4733 ;
  assign n4735 = n595 & n4734 ;
  assign n4736 = ~n4732 & ~n4735 ;
  assign n4737 = ~n4729 & n4736 ;
  assign n4738 = n560 & ~n4737 ;
  assign n4739 = n1376 & n2146 ;
  assign n4740 = n2719 & n4739 ;
  assign n4741 = ~n4738 & ~n4740 ;
  assign n4742 = ~x0 & ~n4741 ;
  assign n4743 = n2040 & n2147 ;
  assign n4744 = x0 & n190 ;
  assign n4745 = n708 & n4744 ;
  assign n4746 = n4743 & ~n4745 ;
  assign n4747 = ~n2753 & n4746 ;
  assign n4748 = n4747 ^ n4743 ;
  assign n4749 = ~n4742 & ~n4748 ;
  assign n4750 = n106 & ~n4749 ;
  assign n4751 = ~n4724 & ~n4750 ;
  assign n4752 = n4710 & n4751 ;
  assign n4753 = ~n4596 & n4752 ;
  assign n4754 = ~n205 & ~n1939 ;
  assign n4755 = ~n1946 & ~n4059 ;
  assign n4756 = ~n4754 & ~n4755 ;
  assign n4757 = n1696 & n2412 ;
  assign n4759 = n4757 ^ n135 ;
  assign n4768 = n4759 ^ n4757 ;
  assign n4758 = n4757 ^ n1867 ;
  assign n4760 = n4759 ^ n4758 ;
  assign n4761 = n4760 ^ n4759 ;
  assign n4762 = n4761 ^ n4757 ;
  assign n4763 = x9 & n48 ;
  assign n4764 = n4763 ^ n4760 ;
  assign n4765 = n4764 ^ n4760 ;
  assign n4766 = n4765 ^ n4762 ;
  assign n4767 = n4762 & n4766 ;
  assign n4769 = n4768 ^ n4767 ;
  assign n4770 = n4769 ^ n4762 ;
  assign n4771 = n4757 ^ n148 ;
  assign n4772 = n4767 ^ n4762 ;
  assign n4773 = ~n4771 & n4772 ;
  assign n4774 = n4773 ^ n4757 ;
  assign n4775 = n4770 & ~n4774 ;
  assign n4776 = n4775 ^ n4757 ;
  assign n4777 = n4776 ^ n135 ;
  assign n4778 = n4777 ^ n4757 ;
  assign n4779 = n442 & n4778 ;
  assign n4780 = ~n1944 & ~n2709 ;
  assign n4781 = ~x9 & n1101 ;
  assign n4782 = n822 & n4781 ;
  assign n4785 = n4782 ^ n823 ;
  assign n4786 = n4785 ^ n4782 ;
  assign n4783 = n4782 ^ n614 ;
  assign n4784 = n4783 ^ n4782 ;
  assign n4787 = n4786 ^ n4784 ;
  assign n4788 = n4782 ^ x7 ;
  assign n4789 = n4788 ^ n4782 ;
  assign n4790 = n4789 ^ n4786 ;
  assign n4791 = n4786 & ~n4790 ;
  assign n4792 = n4791 ^ n4786 ;
  assign n4793 = n4787 & n4792 ;
  assign n4794 = n4793 ^ n4791 ;
  assign n4795 = n4794 ^ n4782 ;
  assign n4796 = n4795 ^ n4786 ;
  assign n4797 = ~x6 & n4796 ;
  assign n4798 = n4797 ^ n4782 ;
  assign n4799 = ~n4780 & n4798 ;
  assign n4800 = n98 & n1732 ;
  assign n4801 = n471 & n2265 ;
  assign n4802 = n4800 & n4801 ;
  assign n4803 = ~n4799 & ~n4802 ;
  assign n4804 = n470 & n1732 ;
  assign n4805 = n199 & n1886 ;
  assign n4806 = n4804 & n4805 ;
  assign n4807 = x8 ^ x1 ;
  assign n4808 = n2412 & n4807 ;
  assign n4809 = n4808 ^ x1 ;
  assign n4810 = n4809 ^ n4808 ;
  assign n4811 = n4808 ^ n268 ;
  assign n4812 = n4811 ^ n4808 ;
  assign n4813 = n4810 & n4812 ;
  assign n4814 = n4813 ^ n4808 ;
  assign n4815 = ~x0 & n4814 ;
  assign n4816 = n4815 ^ n4808 ;
  assign n4817 = n1696 & n4816 ;
  assign n4818 = ~n4806 & ~n4817 ;
  assign n4819 = n969 & ~n4818 ;
  assign n4820 = n4803 & ~n4819 ;
  assign n4821 = ~n4779 & n4820 ;
  assign n4822 = x14 & ~n4821 ;
  assign n4823 = n1853 & n2924 ;
  assign n4824 = n1886 & n2945 ;
  assign n4825 = n173 & n4824 ;
  assign n4826 = ~n4823 & ~n4825 ;
  assign n4827 = n777 & ~n4826 ;
  assign n4828 = n87 & n4827 ;
  assign n4829 = n69 & n3174 ;
  assign n4830 = n362 & n4829 ;
  assign n4831 = n4823 & n4830 ;
  assign n4832 = ~n416 & n1699 ;
  assign n4833 = n4713 & n4832 ;
  assign n4834 = n846 & n4833 ;
  assign n4835 = ~n4831 & ~n4834 ;
  assign n4836 = ~n4828 & n4835 ;
  assign n4837 = ~n4822 & n4836 ;
  assign n4838 = n4756 & ~n4837 ;
  assign n4839 = ~x3 & n17 ;
  assign n4840 = n4202 & n4839 ;
  assign n4841 = n300 & n1197 ;
  assign n4842 = n379 & n2242 ;
  assign n4843 = n4841 & n4842 ;
  assign n4844 = ~x4 & n4059 ;
  assign n4845 = x10 & n2242 ;
  assign n4846 = ~n4844 & ~n4845 ;
  assign n4847 = x2 & ~n3286 ;
  assign n4848 = ~n4846 & n4847 ;
  assign n4849 = ~n4843 & ~n4848 ;
  assign n4850 = n4681 & ~n4849 ;
  assign n4851 = n47 & n3155 ;
  assign n4852 = ~n814 & ~n837 ;
  assign n4853 = n3791 & ~n4852 ;
  assign n4854 = n108 & n3363 ;
  assign n4855 = ~n4853 & ~n4854 ;
  assign n4856 = n4851 & ~n4855 ;
  assign n4857 = n281 & n2242 ;
  assign n4858 = n2622 & n4857 ;
  assign n4859 = ~n4856 & ~n4858 ;
  assign n4860 = ~n4850 & n4859 ;
  assign n4861 = ~n4840 & n4860 ;
  assign n4862 = n437 & ~n4861 ;
  assign n4863 = n708 & n1899 ;
  assign n4864 = n2147 & n3877 ;
  assign n4865 = n191 & n4864 ;
  assign n4866 = ~n4863 & ~n4865 ;
  assign n4867 = n27 & ~n4866 ;
  assign n4868 = n87 & n3828 ;
  assign n4869 = n1835 & n4868 ;
  assign n4870 = ~n128 & ~n3051 ;
  assign n4871 = ~x2 & ~x4 ;
  assign n4872 = n404 & ~n4871 ;
  assign n4873 = n2974 & n4872 ;
  assign n4874 = ~n4870 & n4873 ;
  assign n4875 = n129 & n4072 ;
  assign n4876 = ~n1705 & ~n1865 ;
  assign n4877 = n1914 & ~n4876 ;
  assign n4878 = n4875 & n4877 ;
  assign n4879 = ~n4874 & ~n4878 ;
  assign n4880 = ~n4869 & n4879 ;
  assign n4881 = ~x5 & ~n4880 ;
  assign n4882 = ~n4867 & ~n4881 ;
  assign n4883 = n483 & ~n4882 ;
  assign n4884 = n27 & n2083 ;
  assign n4885 = n1753 & n4884 ;
  assign n4886 = n3321 & n4885 ;
  assign n4887 = ~x5 & n2233 ;
  assign n4888 = ~n1760 & ~n4887 ;
  assign n4889 = n3321 & ~n4888 ;
  assign n4890 = n84 & ~n2835 ;
  assign n4891 = n1376 & n4890 ;
  assign n4892 = ~n4889 & ~n4891 ;
  assign n4893 = n471 & ~n4892 ;
  assign n4894 = ~x11 & n230 ;
  assign n4895 = n1764 & n4894 ;
  assign n4896 = n34 & n1955 ;
  assign n4897 = n4895 & n4896 ;
  assign n4898 = n3227 & n4897 ;
  assign n4899 = ~n4893 & ~n4898 ;
  assign n4900 = ~n4886 & n4899 ;
  assign n4901 = ~n4883 & n4900 ;
  assign n4902 = ~n4862 & n4901 ;
  assign n4903 = n606 & ~n4902 ;
  assign n4904 = ~x2 & n3243 ;
  assign n4905 = ~x5 & n190 ;
  assign n4906 = n4904 & n4905 ;
  assign n4907 = x4 & x10 ;
  assign n4908 = n3978 & n4907 ;
  assign n4909 = n2446 & n4908 ;
  assign n4910 = n571 & n992 ;
  assign n4911 = ~x4 & n3684 ;
  assign n4912 = n4910 & n4911 ;
  assign n4913 = ~n4909 & ~n4912 ;
  assign n4914 = ~x0 & n105 ;
  assign n4915 = ~n4913 & n4914 ;
  assign n4916 = ~x4 & n286 ;
  assign n4917 = n4627 & n4916 ;
  assign n4918 = n920 & n4917 ;
  assign n4919 = n230 & n4918 ;
  assign n4920 = ~n4915 & ~n4919 ;
  assign n4923 = n4920 ^ x8 ;
  assign n4924 = n4923 ^ n4920 ;
  assign n4921 = n4920 ^ x7 ;
  assign n4922 = n4921 ^ n4920 ;
  assign n4925 = n4924 ^ n4922 ;
  assign n4926 = ~n3286 & n4210 ;
  assign n4927 = x0 & n3296 ;
  assign n4928 = n4911 & n4927 ;
  assign n4929 = ~n4926 & ~n4928 ;
  assign n4930 = n4929 ^ n4920 ;
  assign n4931 = n4930 ^ n4920 ;
  assign n4932 = n4931 ^ n4924 ;
  assign n4933 = n4924 & ~n4932 ;
  assign n4934 = n4933 ^ n4924 ;
  assign n4935 = ~n4925 & n4934 ;
  assign n4936 = n4935 ^ n4933 ;
  assign n4937 = n4936 ^ n4920 ;
  assign n4938 = n4937 ^ n4924 ;
  assign n4939 = ~x9 & ~n4938 ;
  assign n4940 = n4939 ^ n4920 ;
  assign n4941 = ~n4906 & n4940 ;
  assign n4942 = n1716 & ~n4941 ;
  assign n4943 = ~n4903 & ~n4942 ;
  assign n4944 = ~n4838 & n4943 ;
  assign n4945 = ~n2927 & ~n3099 ;
  assign n4946 = ~n48 & ~n4945 ;
  assign n4947 = n4522 & n4730 ;
  assign n4948 = n1944 & n4947 ;
  assign n4949 = n3864 ^ x13 ;
  assign n4950 = n4949 ^ n3864 ;
  assign n4951 = n307 & n1914 ;
  assign n4952 = n4951 ^ n3864 ;
  assign n4953 = n4952 ^ n3864 ;
  assign n4954 = ~n4950 & n4953 ;
  assign n4955 = n4954 ^ n3864 ;
  assign n4956 = x12 & n4955 ;
  assign n4957 = n4956 ^ n3864 ;
  assign n4958 = n1705 & n4957 ;
  assign n4959 = n1454 ^ n530 ;
  assign n4960 = n4959 ^ n4539 ;
  assign n4961 = n1597 ^ n141 ;
  assign n4962 = n1454 & ~n4961 ;
  assign n4963 = n4962 ^ n141 ;
  assign n4964 = n4960 & n4963 ;
  assign n4965 = n4964 ^ n4962 ;
  assign n4966 = n4965 ^ n141 ;
  assign n4967 = n4966 ^ n1454 ;
  assign n4968 = n4539 & n4967 ;
  assign n4969 = ~n4958 & ~n4968 ;
  assign n4970 = n3408 & ~n4969 ;
  assign n4971 = n754 & n2381 ;
  assign n4972 = n3757 & n4971 ;
  assign n4973 = ~n4563 & ~n4972 ;
  assign n4974 = n442 & ~n4973 ;
  assign n4975 = n1914 & n3639 ;
  assign n4976 = ~x3 & ~n3865 ;
  assign n4977 = ~n572 & n4976 ;
  assign n4978 = ~n4975 & ~n4977 ;
  assign n4979 = n811 & n2083 ;
  assign n4980 = ~n4978 & n4979 ;
  assign n4981 = ~n4974 & ~n4980 ;
  assign n4982 = ~n4970 & n4981 ;
  assign n4983 = ~n4948 & n4982 ;
  assign n4984 = x14 & ~n4983 ;
  assign n4985 = n124 & n1706 ;
  assign n4986 = n4525 & n4985 ;
  assign n4987 = ~n4947 & ~n4986 ;
  assign n4988 = x0 & ~n4987 ;
  assign n4989 = ~n4521 & ~n4988 ;
  assign n4990 = x13 & ~n4989 ;
  assign n4991 = ~n4534 & ~n4990 ;
  assign n4992 = ~n4984 & n4991 ;
  assign n4993 = n4946 & ~n4992 ;
  assign n4994 = n4944 & ~n4993 ;
  assign n4995 = n4753 & n4994 ;
  assign n4996 = n396 & n3363 ;
  assign n4997 = n129 & n265 ;
  assign n4998 = n65 & n4997 ;
  assign n4999 = ~n4996 & ~n4998 ;
  assign n5000 = ~n2383 & ~n4999 ;
  assign n5001 = ~x6 & x11 ;
  assign n5002 = n4229 & n5001 ;
  assign n5003 = n1329 & n2580 ;
  assign n5004 = n5002 & n5003 ;
  assign n5005 = n3114 & n3601 ;
  assign n5006 = n823 & n5005 ;
  assign n5007 = ~n5004 & ~n5006 ;
  assign n5008 = ~n5000 & n5007 ;
  assign n5009 = n4711 & ~n5008 ;
  assign n5010 = ~n802 & n3791 ;
  assign n5011 = n3801 & n4894 ;
  assign n5012 = ~n5010 & ~n5011 ;
  assign n5013 = ~x1 & n2565 ;
  assign n5014 = ~n5012 & n5013 ;
  assign n5015 = n334 & n1955 ;
  assign n5016 = n1058 & n5015 ;
  assign n5017 = n404 & n2861 ;
  assign n5018 = n3466 & n5017 ;
  assign n5019 = n230 & n2147 ;
  assign n5020 = n963 & n5019 ;
  assign n5021 = x12 ^ x3 ;
  assign n5022 = n5020 & n5021 ;
  assign n5023 = ~n5018 & ~n5022 ;
  assign n5024 = ~n5016 & n5023 ;
  assign n5025 = n2099 & ~n5024 ;
  assign n5026 = ~x5 & n2861 ;
  assign n5027 = ~n5019 & ~n5026 ;
  assign n5028 = n431 & n1865 ;
  assign n5029 = n557 & n5028 ;
  assign n5030 = ~n5027 & n5029 ;
  assign n5031 = ~n5025 & ~n5030 ;
  assign n5032 = ~n5014 & n5031 ;
  assign n5033 = n3162 & ~n5032 ;
  assign n5034 = ~n5009 & ~n5033 ;
  assign n5035 = n281 & n431 ;
  assign n5036 = n2134 & n5035 ;
  assign n5037 = n91 & n2834 ;
  assign n5038 = n19 & ~n1141 ;
  assign n5039 = ~n3185 & ~n5038 ;
  assign n5040 = n5037 & ~n5039 ;
  assign n5041 = ~n5036 & ~n5040 ;
  assign n5042 = ~x3 & n281 ;
  assign n5043 = ~n1776 & ~n3768 ;
  assign n5044 = n5042 & ~n5043 ;
  assign n5045 = n763 & n1867 ;
  assign n5046 = ~n231 & ~n941 ;
  assign n5047 = n2095 & ~n5046 ;
  assign n5048 = n5047 ^ n231 ;
  assign n5049 = n5048 ^ n5047 ;
  assign n5050 = n5047 ^ n1817 ;
  assign n5051 = n5050 ^ n5047 ;
  assign n5052 = ~n5049 & n5051 ;
  assign n5053 = n5052 ^ n5047 ;
  assign n5054 = ~x0 & n5053 ;
  assign n5055 = n5054 ^ n5047 ;
  assign n5056 = x14 & n5055 ;
  assign n5057 = ~n5045 & ~n5056 ;
  assign n5058 = n230 & ~n5057 ;
  assign n5059 = ~n5044 & ~n5058 ;
  assign n5060 = n2434 & ~n5059 ;
  assign n5061 = n1717 & n2686 ;
  assign n5062 = n1192 & n5061 ;
  assign n5063 = ~x3 & ~x8 ;
  assign n5064 = n236 & n2649 ;
  assign n5065 = n5063 & n5064 ;
  assign n5066 = n1104 & n5065 ;
  assign n5067 = ~x3 & n3306 ;
  assign n5068 = ~x14 & ~n1847 ;
  assign n5069 = ~n1699 & ~n5068 ;
  assign n5070 = n5067 & n5069 ;
  assign n5071 = n2120 & n2861 ;
  assign n5072 = ~n5070 & ~n5071 ;
  assign n5073 = ~n5066 & n5072 ;
  assign n5074 = n2561 & ~n5073 ;
  assign n5075 = ~x0 & n1197 ;
  assign n5076 = n300 & n1716 ;
  assign n5077 = n5075 & n5076 ;
  assign n5078 = n837 & n3927 ;
  assign n5079 = ~n2307 & ~n5078 ;
  assign n5080 = n3768 & ~n5079 ;
  assign n5081 = n2120 & ~n2307 ;
  assign n5082 = ~n1914 & n5081 ;
  assign n5083 = ~n1328 & n5082 ;
  assign n5084 = ~n5080 & ~n5083 ;
  assign n5085 = ~n5077 & n5084 ;
  assign n5086 = n3923 & ~n5085 ;
  assign n5087 = ~n5074 & ~n5086 ;
  assign n5088 = ~n5062 & n5087 ;
  assign n5089 = ~n5060 & n5088 ;
  assign n5090 = n5089 ^ x5 ;
  assign n5091 = n5090 ^ n5089 ;
  assign n5092 = n5091 ^ n5041 ;
  assign n5093 = n2307 & n2682 ;
  assign n5094 = ~n281 & ~n3365 ;
  assign n5095 = ~n2304 & ~n2686 ;
  assign n5096 = ~n5094 & ~n5095 ;
  assign n5097 = ~n5093 & ~n5096 ;
  assign n5098 = n2823 & ~n5097 ;
  assign n5099 = n992 & n5098 ;
  assign n5100 = n992 & n2434 ;
  assign n5101 = n1699 & n2682 ;
  assign n5102 = n5100 & n5101 ;
  assign n5103 = ~x8 & n988 ;
  assign n5104 = x13 & n431 ;
  assign n5105 = ~n1712 & ~n5104 ;
  assign n5106 = n5103 & ~n5105 ;
  assign n5107 = n3243 & n5106 ;
  assign n5108 = ~n5102 & ~n5107 ;
  assign n5109 = n344 & n3366 ;
  assign n5110 = x6 & n5109 ;
  assign n5111 = n3365 & n3923 ;
  assign n5112 = ~n5017 & ~n5111 ;
  assign n5113 = ~n5110 & n5112 ;
  assign n5114 = n5113 ^ x0 ;
  assign n5115 = n5114 ^ n5113 ;
  assign n5116 = n5115 ^ n5108 ;
  assign n5117 = n3848 ^ n1041 ;
  assign n5118 = n1041 & n5117 ;
  assign n5119 = n5118 ^ n5113 ;
  assign n5120 = n5119 ^ n1041 ;
  assign n5121 = ~n5116 & ~n5120 ;
  assign n5122 = n5121 ^ n5118 ;
  assign n5123 = n5122 ^ n1041 ;
  assign n5124 = n5108 & n5123 ;
  assign n5125 = n5124 ^ n5108 ;
  assign n5126 = ~n5099 & n5125 ;
  assign n5127 = n5126 ^ x3 ;
  assign n5128 = ~n5126 & ~n5127 ;
  assign n5129 = n5128 ^ n5089 ;
  assign n5130 = n5129 ^ n5126 ;
  assign n5131 = ~n5092 & n5130 ;
  assign n5132 = n5131 ^ n5128 ;
  assign n5133 = n5132 ^ n5126 ;
  assign n5134 = n5041 & ~n5133 ;
  assign n5135 = n5134 ^ n5041 ;
  assign n5136 = n333 & ~n5135 ;
  assign n5137 = n5136 ^ n5034 ;
  assign n5138 = x1 & n4603 ;
  assign n5139 = n5017 & n5138 ;
  assign n5140 = x4 ^ x0 ;
  assign n5141 = n322 & n2099 ;
  assign n5142 = n405 & n5141 ;
  assign n5143 = n129 & ~n4228 ;
  assign n5144 = n5143 ^ n2824 ;
  assign n5145 = n5144 ^ n533 ;
  assign n5146 = n5145 ^ n5143 ;
  assign n5147 = n5146 ^ n5145 ;
  assign n5148 = n5145 ^ n2242 ;
  assign n5149 = n5148 ^ n5144 ;
  assign n5150 = ~n5147 & ~n5149 ;
  assign n5151 = n5150 ^ n2242 ;
  assign n5152 = n377 & n2242 ;
  assign n5153 = n5152 ^ n5144 ;
  assign n5154 = n5151 & ~n5153 ;
  assign n5155 = n5154 ^ n5152 ;
  assign n5156 = ~n5144 & n5155 ;
  assign n5157 = n5156 ^ n5150 ;
  assign n5158 = n5157 ^ n2824 ;
  assign n5159 = n5158 ^ n2242 ;
  assign n5160 = ~n5142 & ~n5159 ;
  assign n5161 = n1776 & ~n5160 ;
  assign n5162 = n5161 ^ n5140 ;
  assign n5163 = n2231 & n3268 ;
  assign n5164 = n1168 & n1706 ;
  assign n5165 = x1 & n5164 ;
  assign n5166 = ~n5163 & ~n5165 ;
  assign n5167 = n5166 ^ x0 ;
  assign n5168 = n5167 ^ n5166 ;
  assign n5169 = n231 & n3365 ;
  assign n5170 = n52 & n5169 ;
  assign n5171 = n5170 ^ n5166 ;
  assign n5172 = n5168 & ~n5171 ;
  assign n5173 = n5172 ^ n5166 ;
  assign n5174 = n5173 ^ n5140 ;
  assign n5175 = ~n5162 & ~n5174 ;
  assign n5176 = n5175 ^ n5172 ;
  assign n5177 = n5176 ^ n5166 ;
  assign n5178 = n5177 ^ n5161 ;
  assign n5179 = n5140 & n5178 ;
  assign n5180 = n5179 ^ n5140 ;
  assign n5181 = n5180 ^ n5161 ;
  assign n5182 = n5103 & n5181 ;
  assign n5183 = n34 & n3017 ;
  assign n5184 = n470 & n2242 ;
  assign n5185 = n2818 & n5184 ;
  assign n5186 = ~n1959 & n5185 ;
  assign n5187 = ~n5183 & ~n5186 ;
  assign n5188 = ~x8 & ~n5187 ;
  assign n5189 = n801 & n1336 ;
  assign n5190 = ~n2242 & ~n5189 ;
  assign n5191 = ~x6 & n540 ;
  assign n5192 = ~n5190 & n5191 ;
  assign n5193 = n437 & n3274 ;
  assign n5194 = ~n5192 & ~n5193 ;
  assign n5195 = n5194 ^ n281 ;
  assign n5196 = n388 & ~n1808 ;
  assign n5197 = ~x5 & n3051 ;
  assign n5198 = n1336 & n5197 ;
  assign n5199 = ~n5196 & ~n5198 ;
  assign n5200 = n5001 & ~n5199 ;
  assign n5201 = ~x1 & n1711 ;
  assign n5202 = n992 & n3365 ;
  assign n5203 = n5201 & n5202 ;
  assign n5204 = ~n5200 & ~n5203 ;
  assign n5205 = ~x0 & ~n5204 ;
  assign n5206 = n5205 ^ n5042 ;
  assign n5207 = n5195 & n5206 ;
  assign n5208 = n5207 ^ n5205 ;
  assign n5209 = n5042 & n5208 ;
  assign n5210 = n5209 ^ x3 ;
  assign n5211 = ~n5188 & ~n5210 ;
  assign n5212 = ~n5182 & n5211 ;
  assign n5213 = ~x0 & ~x8 ;
  assign n5214 = n2242 & n3296 ;
  assign n5215 = n1192 & n4844 ;
  assign n5216 = n236 & n1197 ;
  assign n5217 = ~x5 & n2434 ;
  assign n5218 = n5216 & n5217 ;
  assign n5219 = ~n5215 & ~n5218 ;
  assign n5220 = ~n5214 & n5219 ;
  assign n5221 = n5213 & ~n5220 ;
  assign n5222 = x1 & n5221 ;
  assign n5223 = n230 & n1104 ;
  assign n5224 = n34 & n2083 ;
  assign n5225 = n5223 & n5224 ;
  assign n5226 = n230 & n470 ;
  assign n5227 = n5226 ^ n1808 ;
  assign n5228 = n5226 ^ n2242 ;
  assign n5229 = n5228 ^ n2242 ;
  assign n5230 = n281 & n543 ;
  assign n5231 = n5230 ^ n2242 ;
  assign n5232 = ~n5229 & ~n5231 ;
  assign n5233 = n5232 ^ n2242 ;
  assign n5234 = n5227 & n5233 ;
  assign n5235 = n5234 ^ n1808 ;
  assign n5236 = ~n1198 & n5235 ;
  assign n5237 = ~n5225 & ~n5236 ;
  assign n5238 = n405 & ~n5237 ;
  assign n5239 = n237 & n313 ;
  assign n5240 = n3154 & n5239 ;
  assign n5241 = ~n4857 & ~n5240 ;
  assign n5242 = n540 & ~n5241 ;
  assign n5243 = ~n5238 & ~n5242 ;
  assign n5244 = n1192 & n5197 ;
  assign n5245 = ~n2961 & ~n5244 ;
  assign n5246 = ~x0 & ~n5245 ;
  assign n5247 = n1576 & ~n2136 ;
  assign n5248 = ~n3023 & n5247 ;
  assign n5249 = ~n5246 & ~n5248 ;
  assign n5250 = n1459 & ~n5249 ;
  assign n5251 = ~n2269 & ~n4627 ;
  assign n5252 = n4844 & ~n5251 ;
  assign n5253 = n2685 & ~n5252 ;
  assign n5254 = n79 & n801 ;
  assign n5255 = ~n4845 & ~n5254 ;
  assign n5256 = n5255 ^ n2242 ;
  assign n5257 = n5255 ^ x1 ;
  assign n5258 = n5257 ^ n5255 ;
  assign n5259 = n5258 ^ n5253 ;
  assign n5260 = n5259 ^ n5252 ;
  assign n5261 = ~n5256 & ~n5260 ;
  assign n5262 = n5261 ^ n5255 ;
  assign n5263 = n5253 & ~n5262 ;
  assign n5264 = n5263 ^ n5253 ;
  assign n5265 = n5264 ^ n2685 ;
  assign n5266 = ~n5250 & ~n5265 ;
  assign n5267 = n5243 & n5266 ;
  assign n5268 = ~n5222 & n5267 ;
  assign n5269 = x6 & ~n5268 ;
  assign n5270 = ~x12 & n5223 ;
  assign n5271 = ~n281 & ~n5270 ;
  assign n5272 = n3229 & n5201 ;
  assign n5273 = ~n5271 & n5272 ;
  assign n5274 = x0 & n5273 ;
  assign n5275 = ~x11 & n2914 ;
  assign n5276 = ~n2104 & ~n5275 ;
  assign n5277 = n2682 & ~n5276 ;
  assign n5278 = ~n47 & n470 ;
  assign n5279 = n4894 & n5278 ;
  assign n5280 = ~n2242 & n5279 ;
  assign n5281 = ~x4 & n34 ;
  assign n5282 = n281 & n5281 ;
  assign n5283 = n2236 & n5282 ;
  assign n5284 = ~n5280 & ~n5283 ;
  assign n5285 = ~n5277 & n5284 ;
  assign n5286 = n1712 & ~n5285 ;
  assign n5287 = n3173 & n3587 ;
  assign n5288 = ~n5286 & ~n5287 ;
  assign n5289 = x3 & n5288 ;
  assign n5290 = ~n5274 & n5289 ;
  assign n5291 = ~n5269 & n5290 ;
  assign n5292 = ~n5212 & ~n5291 ;
  assign n5293 = n2682 & ~n3164 ;
  assign n5294 = ~n2269 & n3467 ;
  assign n5295 = n5294 ^ x0 ;
  assign n5296 = n5295 ^ n5294 ;
  assign n5297 = n5294 ^ n570 ;
  assign n5298 = n5297 ^ n5294 ;
  assign n5299 = ~n5296 & n5298 ;
  assign n5300 = n5299 ^ n5294 ;
  assign n5301 = x12 & n5300 ;
  assign n5302 = n5301 ^ n5294 ;
  assign n5303 = n5103 & n5302 ;
  assign n5304 = ~n5293 & ~n5303 ;
  assign n5305 = ~n2383 & ~n5304 ;
  assign n5306 = x6 & n913 ;
  assign n5307 = n236 & n518 ;
  assign n5308 = n2914 & n5307 ;
  assign n5309 = n388 & n2954 ;
  assign n5310 = n1207 & n5309 ;
  assign n5311 = ~n5308 & ~n5310 ;
  assign n5312 = n5306 & ~n5311 ;
  assign n5313 = ~n5305 & ~n5312 ;
  assign n5314 = ~n5292 & n5313 ;
  assign n5315 = ~n5139 & n5314 ;
  assign n5316 = n5315 ^ x2 ;
  assign n5317 = n5316 ^ n5315 ;
  assign n5318 = x4 & n837 ;
  assign n5319 = n5071 & n5318 ;
  assign n5320 = x5 & n5319 ;
  assign n5321 = n5320 ^ x1 ;
  assign n5322 = ~n2096 & n2242 ;
  assign n5323 = n431 & n1939 ;
  assign n5324 = n5323 ^ x5 ;
  assign n5325 = n5324 ^ x6 ;
  assign n5331 = n5325 ^ n5324 ;
  assign n5326 = n5325 ^ n5323 ;
  assign n5327 = n5326 ^ n2567 ;
  assign n5328 = n5325 ^ n2567 ;
  assign n5329 = n5328 ^ n5324 ;
  assign n5330 = ~n5327 & n5329 ;
  assign n5332 = n5331 ^ n5330 ;
  assign n5333 = x11 & n2298 ;
  assign n5334 = n5333 ^ n5325 ;
  assign n5335 = ~n5331 & ~n5334 ;
  assign n5336 = n5335 ^ n5333 ;
  assign n5337 = ~n5332 & n5336 ;
  assign n5338 = n5337 ^ n5330 ;
  assign n5339 = n5338 ^ n5325 ;
  assign n5340 = n5339 ^ x5 ;
  assign n5341 = n5340 ^ n5324 ;
  assign n5342 = ~n5322 & n5341 ;
  assign n5343 = n281 & ~n5342 ;
  assign n5344 = ~x3 & n2242 ;
  assign n5345 = n232 & n5344 ;
  assign n5346 = n3778 & n5345 ;
  assign n5347 = n2925 ^ x11 ;
  assign n5348 = n5347 ^ n2925 ;
  assign n5349 = n2925 ^ n2861 ;
  assign n5350 = n5349 ^ n2925 ;
  assign n5351 = ~n5348 & n5350 ;
  assign n5352 = n5351 ^ n2925 ;
  assign n5353 = x4 & n5352 ;
  assign n5354 = n5353 ^ n2925 ;
  assign n5355 = n3560 & n5354 ;
  assign n5356 = n2248 & n5035 ;
  assign n5357 = ~n5355 & ~n5356 ;
  assign n5358 = n4132 & ~n5357 ;
  assign n5359 = ~n5346 & ~n5358 ;
  assign n5360 = ~n5343 & n5359 ;
  assign n5361 = n5360 ^ x0 ;
  assign n5362 = n5361 ^ n5360 ;
  assign n5363 = n182 & n4839 ;
  assign n5364 = n5223 & n5363 ;
  assign n5365 = x5 & x14 ;
  assign n5366 = ~n664 & ~n5104 ;
  assign n5367 = ~x4 & x11 ;
  assign n5368 = ~n2434 & ~n5367 ;
  assign n5369 = n2095 & ~n5368 ;
  assign n5370 = ~n5366 & n5369 ;
  assign n5371 = n5365 & n5370 ;
  assign n5372 = n64 & n3155 ;
  assign n5373 = ~n2566 & ~n5372 ;
  assign n5374 = n5373 ^ n1939 ;
  assign n5375 = n5374 ^ n5373 ;
  assign n5376 = n5373 ^ n5202 ;
  assign n5377 = n5376 ^ n5373 ;
  assign n5378 = n5375 & n5377 ;
  assign n5379 = n5378 ^ n5373 ;
  assign n5380 = ~x5 & ~n5379 ;
  assign n5381 = n5380 ^ n5373 ;
  assign n5382 = ~n5371 & n5381 ;
  assign n5383 = n281 & ~n5382 ;
  assign n5384 = ~n5364 & ~n5383 ;
  assign n5385 = n5384 ^ n5360 ;
  assign n5386 = ~n5362 & n5385 ;
  assign n5387 = n5386 ^ n5360 ;
  assign n5388 = n5387 ^ n5320 ;
  assign n5389 = n5321 & n5388 ;
  assign n5390 = n5389 ^ n5386 ;
  assign n5391 = n5390 ^ n5360 ;
  assign n5392 = n5391 ^ x1 ;
  assign n5393 = ~n5320 & n5392 ;
  assign n5394 = n5393 ^ n5320 ;
  assign n5395 = n5394 ^ n5320 ;
  assign n5396 = n5395 ^ n5315 ;
  assign n5397 = ~n5317 & n5396 ;
  assign n5398 = n5397 ^ n5315 ;
  assign n5399 = n5398 ^ n5034 ;
  assign n5400 = ~n5137 & n5399 ;
  assign n5401 = n5400 ^ n5397 ;
  assign n5402 = n5401 ^ n5315 ;
  assign n5403 = n5402 ^ n5136 ;
  assign n5404 = n5034 & ~n5403 ;
  assign n5405 = n5404 ^ n5034 ;
  assign n5406 = n1704 & ~n5405 ;
  assign n5407 = n4995 & ~n5406 ;
  assign n5408 = ~n4519 & n5407 ;
  assign n5409 = n5408 ^ n4227 ;
  assign n5410 = x3 & n2696 ;
  assign n5411 = ~x4 & n2231 ;
  assign n5412 = n5410 & n5411 ;
  assign n5413 = n1535 & n5037 ;
  assign n5414 = ~n1000 & ~n2235 ;
  assign n5415 = ~n5413 & ~n5414 ;
  assign n5416 = ~n5412 & n5415 ;
  assign n5417 = n3989 & ~n5416 ;
  assign n5418 = x3 & x14 ;
  assign n5419 = n24 & n2233 ;
  assign n5420 = ~n597 & n5419 ;
  assign n5421 = n256 & n1722 ;
  assign n5422 = n3845 & n5421 ;
  assign n5423 = ~n5420 & ~n5422 ;
  assign n5424 = n5418 & ~n5423 ;
  assign n5425 = ~x3 & x14 ;
  assign n5426 = ~n180 & ~n5425 ;
  assign n5427 = n277 & ~n5426 ;
  assign n5428 = ~n519 & ~n5427 ;
  assign n5429 = ~x6 & ~x12 ;
  assign n5430 = ~n5428 & n5429 ;
  assign n5431 = ~n2969 & ~n5430 ;
  assign n5432 = x2 & n4907 ;
  assign n5433 = ~n5431 & n5432 ;
  assign n5434 = n5046 ^ n127 ;
  assign n5435 = x6 & ~n5434 ;
  assign n5436 = n5435 ^ n127 ;
  assign n5437 = n1101 & n5436 ;
  assign n5438 = n530 & n1732 ;
  assign n5439 = ~n5437 & ~n5438 ;
  assign n5440 = n4679 & ~n5439 ;
  assign n5441 = ~n1448 & ~n2096 ;
  assign n5442 = ~x2 & ~n64 ;
  assign n5443 = ~x7 & ~n5442 ;
  assign n5444 = n5441 & n5443 ;
  assign n5445 = n174 & n5418 ;
  assign n5446 = n377 & n2635 ;
  assign n5447 = n5445 & n5446 ;
  assign n5448 = x12 & n1716 ;
  assign n5449 = n1994 & n5448 ;
  assign n5450 = n1101 & n5449 ;
  assign n5451 = ~n5447 & ~n5450 ;
  assign n5452 = ~n5444 & n5451 ;
  assign n5453 = ~x7 & n2095 ;
  assign n5454 = n1031 & n5453 ;
  assign n5455 = n377 & n4681 ;
  assign n5456 = ~n5454 & ~n5455 ;
  assign n5457 = n1255 & ~n5456 ;
  assign n5458 = n5452 & ~n5457 ;
  assign n5459 = ~n5440 & n5458 ;
  assign n5460 = n3085 & ~n5459 ;
  assign n5461 = ~x2 & ~n231 ;
  assign n5462 = n1462 & n5461 ;
  assign n5463 = ~n64 & ~n5462 ;
  assign n5464 = n2861 & ~n5463 ;
  assign n5465 = n1955 & n5042 ;
  assign n5466 = n2159 & n4726 ;
  assign n5467 = ~n5465 & ~n5466 ;
  assign n5468 = ~n5464 & n5467 ;
  assign n5469 = n2652 & ~n5468 ;
  assign n5470 = n71 & n3355 ;
  assign n5471 = n2095 & n5470 ;
  assign n5472 = ~n5469 & ~n5471 ;
  assign n5473 = ~n5460 & n5472 ;
  assign n5474 = ~n5433 & n5473 ;
  assign n5475 = n1632 & ~n5474 ;
  assign n5476 = ~n5424 & ~n5475 ;
  assign n5477 = n1732 & n2355 ;
  assign n5478 = ~x9 & n1147 ;
  assign n5479 = ~n1448 & n5478 ;
  assign n5480 = n5477 & n5479 ;
  assign n5481 = n1729 & n3671 ;
  assign n5482 = n1960 & n5481 ;
  assign n5483 = n1817 & n5223 ;
  assign n5484 = ~n526 & n2095 ;
  assign n5485 = n281 & n5484 ;
  assign n5486 = ~n5483 & ~n5485 ;
  assign n5487 = n1724 & ~n5486 ;
  assign n5488 = ~n526 & n658 ;
  assign n5489 = n1535 & ~n3591 ;
  assign n5490 = ~n5488 & ~n5489 ;
  assign n5491 = n230 & ~n5490 ;
  assign n5492 = n3144 & ~n5491 ;
  assign n5493 = n4839 & ~n5492 ;
  assign n5494 = x3 & n2945 ;
  assign n5497 = n2653 ^ x4 ;
  assign n5498 = n5497 ^ n2653 ;
  assign n5495 = n2653 ^ n526 ;
  assign n5496 = n5495 ^ n2653 ;
  assign n5499 = n5498 ^ n5496 ;
  assign n5500 = n4713 ^ n2653 ;
  assign n5501 = n5500 ^ n2653 ;
  assign n5502 = n5501 ^ n5498 ;
  assign n5503 = n5498 & n5502 ;
  assign n5504 = n5503 ^ n5498 ;
  assign n5505 = ~n5499 & n5504 ;
  assign n5506 = n5505 ^ n5503 ;
  assign n5507 = n5506 ^ n2653 ;
  assign n5508 = n5507 ^ n5498 ;
  assign n5509 = ~x10 & n5508 ;
  assign n5510 = n5509 ^ n2653 ;
  assign n5511 = n5494 & n5510 ;
  assign n5512 = n1817 & ~n3591 ;
  assign n5513 = ~x3 & n3927 ;
  assign n5514 = ~n5512 & ~n5513 ;
  assign n5515 = ~n1000 & ~n5514 ;
  assign n5516 = ~x4 & n5515 ;
  assign n5517 = ~n5511 & ~n5516 ;
  assign n5518 = ~n5493 & n5517 ;
  assign n5519 = ~n5487 & n5518 ;
  assign n5520 = n5519 ^ x2 ;
  assign n5521 = n5520 ^ n5519 ;
  assign n5522 = n5521 ^ n5482 ;
  assign n5523 = ~n595 & ~n2705 ;
  assign n5524 = n1835 & ~n5523 ;
  assign n5525 = ~n1000 & n1960 ;
  assign n5526 = ~n5524 & ~n5525 ;
  assign n5527 = n1192 & ~n5526 ;
  assign n5528 = n2113 & n5425 ;
  assign n5529 = n595 & n5528 ;
  assign n5530 = ~x13 & n5529 ;
  assign n5531 = n1835 & n3141 ;
  assign n5532 = ~n5410 & ~n5531 ;
  assign n5533 = ~n5530 & n5532 ;
  assign n5534 = ~n5527 & n5533 ;
  assign n5535 = n5534 ^ x6 ;
  assign n5536 = ~n5534 & ~n5535 ;
  assign n5537 = n5536 ^ n5519 ;
  assign n5538 = n5537 ^ n5534 ;
  assign n5539 = n5522 & n5538 ;
  assign n5540 = n5539 ^ n5536 ;
  assign n5541 = n5540 ^ n5534 ;
  assign n5542 = ~n5482 & ~n5541 ;
  assign n5543 = n5542 ^ n5482 ;
  assign n5544 = ~n5480 & ~n5543 ;
  assign n5545 = n5544 ^ x5 ;
  assign n5546 = n5545 ^ n5544 ;
  assign n5547 = n5546 ^ n5476 ;
  assign n5548 = x12 & n2096 ;
  assign n5549 = n5548 ^ n1753 ;
  assign n5550 = n5548 ^ n1255 ;
  assign n5551 = n5550 ^ n1255 ;
  assign n5552 = n1255 ^ n1190 ;
  assign n5553 = ~n5551 & n5552 ;
  assign n5554 = n5553 ^ n1255 ;
  assign n5555 = n5549 & n5554 ;
  assign n5556 = n5555 ^ n1753 ;
  assign n5557 = ~n108 & ~n5556 ;
  assign n5558 = ~x7 & ~n5557 ;
  assign n5559 = n1336 & n1914 ;
  assign n5560 = n100 & n5559 ;
  assign n5561 = ~n5558 & ~n5560 ;
  assign n5562 = n3923 & ~n5561 ;
  assign n5563 = ~x2 & ~x8 ;
  assign n5564 = x6 ^ x3 ;
  assign n5565 = n1147 ^ x6 ;
  assign n5566 = n5565 ^ n1147 ;
  assign n5567 = ~x10 & ~n526 ;
  assign n5568 = n5567 ^ n1147 ;
  assign n5569 = n5566 & n5568 ;
  assign n5570 = n5569 ^ n1147 ;
  assign n5571 = ~n5564 & n5570 ;
  assign n5572 = n2446 & n5571 ;
  assign n5573 = n5563 & n5572 ;
  assign n5574 = n1105 & n5453 ;
  assign n5575 = ~x12 & n3778 ;
  assign n5576 = ~n1817 & ~n5575 ;
  assign n5577 = x8 & ~n5576 ;
  assign n5578 = ~n220 & n5577 ;
  assign n5579 = ~n5574 & ~n5578 ;
  assign n5580 = n203 & ~n5579 ;
  assign n5581 = n1190 & ~n1712 ;
  assign n5582 = n60 & n70 ;
  assign n5583 = ~n2096 & n5582 ;
  assign n5584 = ~n5581 & n5583 ;
  assign n5585 = ~x2 & n281 ;
  assign n5586 = n562 & n5585 ;
  assign n5587 = n71 & n4681 ;
  assign n5588 = ~n5586 & ~n5587 ;
  assign n5589 = ~n5584 & n5588 ;
  assign n5590 = ~n5580 & n5589 ;
  assign n5591 = ~n5573 & n5590 ;
  assign n5592 = x4 & ~n5591 ;
  assign n5593 = ~n5562 & ~n5592 ;
  assign n5594 = n5593 ^ x9 ;
  assign n5595 = ~x9 & n5594 ;
  assign n5596 = n5595 ^ n5544 ;
  assign n5597 = n5596 ^ x9 ;
  assign n5598 = n5547 & n5597 ;
  assign n5599 = n5598 ^ n5595 ;
  assign n5600 = n5599 ^ x9 ;
  assign n5601 = n5476 & ~n5600 ;
  assign n5602 = n5601 ^ n5476 ;
  assign n5603 = ~x0 & ~n5602 ;
  assign n5604 = n1101 & n3012 ;
  assign n5605 = n3308 & n5604 ;
  assign n5606 = n999 & ~n3023 ;
  assign n5607 = n1817 & n5606 ;
  assign n5608 = ~n1000 & n2232 ;
  assign n5609 = n2095 & n2719 ;
  assign n5610 = n2242 & n5609 ;
  assign n5611 = ~n5608 & ~n5610 ;
  assign n5612 = ~n5607 & n5611 ;
  assign n5613 = ~n1198 & ~n5612 ;
  assign n5614 = ~n199 & ~n3864 ;
  assign n5615 = n4976 & ~n5614 ;
  assign n5616 = ~n4951 & ~n5615 ;
  assign n5617 = n2652 & n5478 ;
  assign n5618 = ~n5616 & n5617 ;
  assign n5619 = ~n5613 & ~n5618 ;
  assign n5620 = ~x12 & ~n5619 ;
  assign n5621 = n137 & n842 ;
  assign n5622 = x12 & n287 ;
  assign n5623 = ~n5621 & ~n5622 ;
  assign n5624 = n3350 & ~n5623 ;
  assign n5625 = n1716 & n4617 ;
  assign n5626 = n2943 & n4349 ;
  assign n5627 = ~n220 & n2565 ;
  assign n5628 = n1197 & n2446 ;
  assign n5629 = n2248 & n5628 ;
  assign n5630 = ~n5627 & ~n5629 ;
  assign n5631 = n539 & ~n5630 ;
  assign n5632 = ~x14 & n180 ;
  assign n5633 = n152 & n2128 ;
  assign n5634 = ~n1835 & n5633 ;
  assign n5635 = ~n5632 & n5634 ;
  assign n5636 = ~n5631 & ~n5635 ;
  assign n5637 = ~n5626 & n5636 ;
  assign n5638 = n5637 ^ x8 ;
  assign n5639 = n5638 ^ n5637 ;
  assign n5640 = n5639 ^ n5625 ;
  assign n5641 = ~x3 & n2149 ;
  assign n5642 = ~n2234 & ~n5641 ;
  assign n5643 = n680 & ~n5642 ;
  assign n5644 = ~n1808 & ~n2817 ;
  assign n5645 = n1981 & n5644 ;
  assign n5646 = ~n144 & ~n2818 ;
  assign n5647 = ~x3 & n5646 ;
  assign n5648 = ~n5645 & ~n5647 ;
  assign n5649 = ~n2242 & ~n4907 ;
  assign n5650 = x7 & n5649 ;
  assign n5651 = ~n249 & n5650 ;
  assign n5652 = ~n5648 & n5651 ;
  assign n5653 = ~n3828 & n5652 ;
  assign n5654 = ~n830 & n5653 ;
  assign n5655 = ~n5643 & ~n5654 ;
  assign n5656 = n5655 ^ x14 ;
  assign n5657 = x14 & ~n5656 ;
  assign n5658 = n5657 ^ n5637 ;
  assign n5659 = n5658 ^ x14 ;
  assign n5660 = n5640 & ~n5659 ;
  assign n5661 = n5660 ^ n5657 ;
  assign n5662 = n5661 ^ x14 ;
  assign n5663 = ~n5625 & n5662 ;
  assign n5664 = n5663 ^ n5625 ;
  assign n5665 = ~n5624 & ~n5664 ;
  assign n5666 = n5665 ^ x9 ;
  assign n5667 = n5666 ^ n5665 ;
  assign n5668 = ~n236 & n347 ;
  assign n5669 = ~n334 & ~n5668 ;
  assign n5670 = n3250 & ~n5669 ;
  assign n5671 = ~x7 & n1946 ;
  assign n5672 = n3969 & n5671 ;
  assign n5673 = n70 & n1939 ;
  assign n5674 = ~n5672 & ~n5673 ;
  assign n5675 = n307 & ~n5674 ;
  assign n5676 = n141 & n3366 ;
  assign n5677 = n507 & n5676 ;
  assign n5678 = ~x10 & n3154 ;
  assign n5679 = n197 & n5678 ;
  assign n5680 = ~n1966 & n5679 ;
  assign n5681 = n70 & ~n5680 ;
  assign n5682 = n5680 ^ n2137 ;
  assign n5683 = n5681 ^ n1711 ;
  assign n5684 = n5682 & n5683 ;
  assign n5685 = n5684 ^ n1711 ;
  assign n5686 = n5681 & n5685 ;
  assign n5687 = n5686 ^ n5680 ;
  assign n5688 = n1031 & n5687 ;
  assign n5689 = ~n5677 & ~n5688 ;
  assign n5690 = ~n5675 & n5689 ;
  assign n5691 = ~x6 & ~n5690 ;
  assign n5692 = ~n84 & n1729 ;
  assign n5693 = ~n1247 & n5692 ;
  assign n5694 = n3923 & n5693 ;
  assign n5695 = ~n5691 & ~n5694 ;
  assign n5696 = ~n5670 & n5695 ;
  assign n5697 = n5696 ^ n5665 ;
  assign n5698 = n5667 & n5697 ;
  assign n5699 = n5698 ^ n5665 ;
  assign n5700 = ~n5620 & n5699 ;
  assign n5701 = n512 & ~n5700 ;
  assign n5702 = ~x9 & n277 ;
  assign n5703 = n2095 & n5215 ;
  assign n5704 = n5702 & n5703 ;
  assign n5705 = n1840 & n2381 ;
  assign n5706 = ~x9 & n197 ;
  assign n5707 = ~n3507 & ~n5706 ;
  assign n5708 = ~x4 & n1981 ;
  assign n5709 = ~n5707 & n5708 ;
  assign n5710 = x12 & n2129 ;
  assign n5711 = n1946 & n5710 ;
  assign n5712 = ~n5709 & ~n5711 ;
  assign n5713 = ~n5705 & n5712 ;
  assign n5714 = n5103 & ~n5713 ;
  assign n5715 = n1535 & n2147 ;
  assign n5716 = n659 & n2128 ;
  assign n5717 = ~n5715 & ~n5716 ;
  assign n5718 = x4 & n3560 ;
  assign n5719 = x14 & n5718 ;
  assign n5720 = ~n5717 & n5719 ;
  assign n5721 = n142 & n2636 ;
  assign n5722 = ~n2588 & ~n5721 ;
  assign n5723 = ~n5720 & n5722 ;
  assign n5724 = n230 & ~n5723 ;
  assign n5725 = ~x9 & n136 ;
  assign n5726 = ~n220 & ~n1314 ;
  assign n5727 = n206 & n5726 ;
  assign n5728 = ~n842 & ~n5727 ;
  assign n5729 = n614 & ~n5728 ;
  assign n5730 = ~n5725 & ~n5729 ;
  assign n5731 = n16 & ~n5730 ;
  assign n5732 = ~n5724 & ~n5731 ;
  assign n5733 = ~n5714 & n5732 ;
  assign n5734 = ~n5704 & n5733 ;
  assign n5735 = n920 & ~n5734 ;
  assign n5736 = ~n5701 & ~n5735 ;
  assign n5737 = ~n5605 & n5736 ;
  assign n5738 = ~n5603 & n5737 ;
  assign n5739 = x11 & ~n5738 ;
  assign n5740 = n434 & n5604 ;
  assign n5749 = n3233 & n5411 ;
  assign n5750 = ~n3829 & ~n5749 ;
  assign n5751 = n82 & ~n5750 ;
  assign n5752 = n313 & n3233 ;
  assign n5753 = ~n3848 & ~n5752 ;
  assign n5754 = ~n1765 & n2040 ;
  assign n5755 = ~n5753 & n5754 ;
  assign n5756 = ~n5751 & ~n5755 ;
  assign n5741 = n16 & n529 ;
  assign n5742 = n1365 & n5741 ;
  assign n5743 = n314 & n3285 ;
  assign n5744 = ~n3757 & n5743 ;
  assign n5745 = ~x5 & n3848 ;
  assign n5746 = n1731 & n5745 ;
  assign n5747 = ~n5744 & ~n5746 ;
  assign n5748 = ~n5742 & n5747 ;
  assign n5757 = n5756 ^ n5748 ;
  assign n5758 = n5757 ^ n5756 ;
  assign n5759 = n5756 ^ x10 ;
  assign n5760 = n5759 ^ n5756 ;
  assign n5761 = ~n5758 & n5760 ;
  assign n5762 = n5761 ^ n5756 ;
  assign n5763 = ~x7 & ~n5762 ;
  assign n5764 = n5763 ^ n5756 ;
  assign n5765 = x3 & ~n5764 ;
  assign n5766 = x14 & n4148 ;
  assign n5767 = n3428 & n5766 ;
  assign n5768 = n2233 & n5767 ;
  assign n5769 = ~x2 & ~n5768 ;
  assign n5770 = n312 & n4630 ;
  assign n5771 = n91 & n168 ;
  assign n5772 = ~n5770 & ~n5771 ;
  assign n5773 = n17 & ~n5772 ;
  assign n5774 = n1760 & n2696 ;
  assign n5775 = ~n5773 & ~n5774 ;
  assign n5776 = n2696 & n4887 ;
  assign n5777 = x7 & ~n230 ;
  assign n5778 = ~n663 & ~n960 ;
  assign n5779 = n4839 & ~n5778 ;
  assign n5780 = n5777 & n5779 ;
  assign n5781 = ~n5776 & ~n5780 ;
  assign n5782 = n5775 & n5781 ;
  assign n5783 = n5769 & n5782 ;
  assign n5784 = ~n5765 & n5783 ;
  assign n5785 = ~x7 & n16 ;
  assign n5786 = n281 & n1293 ;
  assign n5787 = n539 & n859 ;
  assign n5788 = n3881 & n5787 ;
  assign n5789 = ~n960 & ~n5788 ;
  assign n5790 = ~n5786 & n5789 ;
  assign n5791 = n5785 & ~n5790 ;
  assign n5792 = n1355 & ~n4630 ;
  assign n5793 = n17 & ~n142 ;
  assign n5794 = ~n5792 & n5793 ;
  assign n5795 = n1336 & n2248 ;
  assign n5796 = n556 & n3808 ;
  assign n5797 = n5795 & n5796 ;
  assign n5798 = ~n5794 & ~n5797 ;
  assign n5799 = n920 & n5798 ;
  assign n5800 = ~n5791 & n5799 ;
  assign n5801 = n5800 ^ n3172 ;
  assign n5802 = ~n1011 & ~n5702 ;
  assign n5803 = n142 & ~n5802 ;
  assign n5804 = ~n606 & ~n4102 ;
  assign n5805 = n498 & n5804 ;
  assign n5806 = ~n4905 & ~n5805 ;
  assign n5807 = ~n5803 & n5806 ;
  assign n5808 = n5807 ^ x4 ;
  assign n5809 = n5808 ^ n5807 ;
  assign n5810 = n317 & n605 ;
  assign n5811 = n5702 ^ n141 ;
  assign n5812 = n5811 ^ n1520 ;
  assign n5813 = n1207 ^ n1011 ;
  assign n5814 = ~n141 & ~n5813 ;
  assign n5815 = n5814 ^ n1011 ;
  assign n5816 = ~n5812 & ~n5815 ;
  assign n5817 = n5816 ^ n5814 ;
  assign n5818 = n5817 ^ n1011 ;
  assign n5819 = n5818 ^ n141 ;
  assign n5820 = ~n1520 & n5819 ;
  assign n5821 = ~n5810 & n5820 ;
  assign n5822 = n5821 ^ n5807 ;
  assign n5823 = n5809 & n5822 ;
  assign n5824 = n5823 ^ n5807 ;
  assign n5825 = n5824 ^ n3172 ;
  assign n5826 = n5801 & ~n5825 ;
  assign n5827 = n5826 ^ n5823 ;
  assign n5828 = n5827 ^ n5807 ;
  assign n5829 = n5828 ^ n5800 ;
  assign n5830 = n3172 & ~n5829 ;
  assign n5831 = n5830 ^ n3172 ;
  assign n5832 = n5831 ^ n5800 ;
  assign n5833 = ~n5784 & ~n5832 ;
  assign n5834 = ~n5740 & ~n5833 ;
  assign n5835 = n3233 ^ n3088 ;
  assign n5836 = n5835 ^ n3088 ;
  assign n5837 = n3088 ^ n2827 ;
  assign n5838 = n5837 ^ n3088 ;
  assign n5839 = n5836 & n5838 ;
  assign n5840 = n5839 ^ n3088 ;
  assign n5841 = ~x4 & n5840 ;
  assign n5842 = n5841 ^ n3088 ;
  assign n5843 = n316 & n5842 ;
  assign n5844 = n1717 & n5766 ;
  assign n5845 = ~n5843 & ~n5844 ;
  assign n5846 = n286 & ~n5845 ;
  assign n5847 = x4 & n91 ;
  assign n5848 = n4211 & n5847 ;
  assign n5849 = ~n5846 & ~n5848 ;
  assign n5850 = n167 & n3848 ;
  assign n5851 = n3483 & n3590 ;
  assign n5852 = n1192 & n5851 ;
  assign n5853 = ~n5850 & ~n5852 ;
  assign n5854 = n142 & ~n5853 ;
  assign n5855 = n5854 ^ x7 ;
  assign n5856 = n5855 ^ n5854 ;
  assign n5857 = ~n167 & ~n1765 ;
  assign n5858 = ~n142 & ~n1914 ;
  assign n5859 = n3355 & n5858 ;
  assign n5860 = n281 & ~n629 ;
  assign n5861 = n4887 & n5860 ;
  assign n5862 = ~n5859 & ~n5861 ;
  assign n5863 = ~n5857 & ~n5862 ;
  assign n5864 = ~n3285 & ~n5741 ;
  assign n5865 = n581 & ~n5864 ;
  assign n5866 = n124 & n5865 ;
  assign n5867 = ~n5863 & ~n5866 ;
  assign n5868 = n5867 ^ n5854 ;
  assign n5869 = ~n5856 & ~n5868 ;
  assign n5870 = n5869 ^ n5854 ;
  assign n5871 = ~n5780 & ~n5870 ;
  assign n5872 = n5849 & n5871 ;
  assign n5873 = x2 & ~n5872 ;
  assign n5874 = ~x0 & ~n5873 ;
  assign n5875 = ~n5834 & ~n5874 ;
  assign n5876 = ~n5739 & ~n5875 ;
  assign n5877 = ~n5417 & n5876 ;
  assign n5878 = n5877 ^ x1 ;
  assign n5879 = n5878 ^ n5877 ;
  assign n5880 = x5 & n1705 ;
  assign n5881 = n2236 & n5880 ;
  assign n5882 = n1527 & n5881 ;
  assign n5883 = ~n182 & n3421 ;
  assign n5884 = n3188 & ~n5883 ;
  assign n5885 = ~n141 & ~n344 ;
  assign n5886 = ~n143 & n3768 ;
  assign n5887 = ~n5885 & n5886 ;
  assign n5888 = ~n5884 & ~n5887 ;
  assign n5889 = n1255 & ~n5888 ;
  assign n5890 = n3670 & n5104 ;
  assign n5891 = ~x12 & ~n831 ;
  assign n5892 = n1232 & ~n5891 ;
  assign n5893 = n1293 & n5892 ;
  assign n5894 = ~n5890 & ~n5893 ;
  assign n5895 = ~n5889 & n5894 ;
  assign n5896 = n1722 & ~n5895 ;
  assign n5897 = n16 & n218 ;
  assign n5898 = x12 ^ x11 ;
  assign n5899 = n5898 ^ x12 ;
  assign n5900 = n5899 ^ x5 ;
  assign n5901 = n231 ^ n19 ;
  assign n5902 = ~n231 & ~n5901 ;
  assign n5903 = n5902 ^ x12 ;
  assign n5904 = n5903 ^ n231 ;
  assign n5905 = ~n5900 & ~n5904 ;
  assign n5906 = n5905 ^ n5902 ;
  assign n5907 = n5906 ^ n231 ;
  assign n5908 = x5 & ~n5907 ;
  assign n5909 = n5897 & n5908 ;
  assign n5910 = ~n5896 & ~n5909 ;
  assign n5911 = ~n5882 & n5910 ;
  assign n5912 = ~n597 & ~n5911 ;
  assign n5913 = n218 & n4607 ;
  assign n5914 = ~x10 & ~n1305 ;
  assign n5915 = ~x0 & n197 ;
  assign n5916 = n799 & n5915 ;
  assign n5917 = ~n5914 & n5916 ;
  assign n5918 = n256 & n843 ;
  assign n5919 = n2247 & n5918 ;
  assign n5920 = ~n5917 & ~n5919 ;
  assign n5921 = n1946 & ~n5920 ;
  assign n5922 = ~n5913 & ~n5921 ;
  assign n5923 = n1031 & ~n5922 ;
  assign n5924 = x14 & n1891 ;
  assign n5925 = n2652 & n5924 ;
  assign n5926 = x3 & n5925 ;
  assign n5927 = ~n2558 & ~n5926 ;
  assign n5928 = n969 & n1759 ;
  assign n5929 = ~n5927 & n5928 ;
  assign n5930 = n4195 & n5671 ;
  assign n5931 = n1872 & n1995 ;
  assign n5932 = ~n5930 & ~n5931 ;
  assign n5933 = n3978 & ~n5932 ;
  assign n5934 = n913 & n5933 ;
  assign n5935 = n106 & n2003 ;
  assign n5936 = n21 & n5671 ;
  assign n5937 = ~n5935 & ~n5936 ;
  assign n5938 = n2247 & ~n5937 ;
  assign n5939 = ~n5934 & ~n5938 ;
  assign n5940 = ~n5929 & n5939 ;
  assign n5941 = n2861 & ~n5940 ;
  assign n5942 = ~n5923 & ~n5941 ;
  assign n5943 = n1898 & n5213 ;
  assign n5944 = n794 & n1627 ;
  assign n5945 = x3 & n5944 ;
  assign n5946 = n5943 & n5945 ;
  assign n5947 = ~n2706 & n5946 ;
  assign n5948 = n5942 & ~n5947 ;
  assign n5949 = n431 & n605 ;
  assign n5950 = n1711 & n5949 ;
  assign n5951 = n4336 & n5950 ;
  assign n5952 = ~x2 & n1718 ;
  assign n5953 = ~n642 & n5952 ;
  assign n5954 = n990 & n4871 ;
  assign n5955 = ~n5953 & ~n5954 ;
  assign n5956 = x7 & ~n5955 ;
  assign n5957 = n197 & n1112 ;
  assign n5958 = n1058 & n5957 ;
  assign n5959 = x0 & ~n5958 ;
  assign n5960 = n646 & n2869 ;
  assign n5961 = ~n1898 & ~n5960 ;
  assign n5962 = n5959 & n5961 ;
  assign n5963 = x5 & ~n1112 ;
  assign n5964 = ~n561 & ~n5963 ;
  assign n5965 = ~x9 & n431 ;
  assign n5966 = ~n434 & ~n5965 ;
  assign n5967 = ~x2 & n5966 ;
  assign n5968 = n2652 & ~n5967 ;
  assign n5969 = ~n5964 & n5968 ;
  assign n5970 = n5962 & ~n5969 ;
  assign n5971 = ~n5956 & n5970 ;
  assign n5972 = n560 & n4713 ;
  assign n5973 = n203 & n5972 ;
  assign n5974 = ~x2 & n21 ;
  assign n5975 = n992 & n5974 ;
  assign n5976 = n4608 & n5975 ;
  assign n5977 = ~n5973 & ~n5976 ;
  assign n5978 = ~x0 & n5977 ;
  assign n5979 = ~x9 & n70 ;
  assign n5980 = n708 & n1112 ;
  assign n5981 = ~n5979 & ~n5980 ;
  assign n5982 = ~x5 & ~n5981 ;
  assign n5983 = n366 & n5975 ;
  assign n5984 = ~n5982 & ~n5983 ;
  assign n5985 = n912 & n1314 ;
  assign n5986 = n343 & n5985 ;
  assign n5987 = n663 & ~n5986 ;
  assign n5988 = n978 & n1805 ;
  assign n5989 = n592 & n5988 ;
  assign n5990 = ~n3781 & ~n5989 ;
  assign n5991 = ~n5987 & n5990 ;
  assign n5992 = n5991 ^ x7 ;
  assign n5993 = n5992 ^ n5991 ;
  assign n5994 = n5993 ^ n5984 ;
  assign n5995 = n1112 & ~n1402 ;
  assign n5996 = ~n1190 & n1346 ;
  assign n5997 = ~n5995 & ~n5996 ;
  assign n5998 = n5997 ^ x5 ;
  assign n5999 = ~n5997 & n5998 ;
  assign n6000 = n5999 ^ n5991 ;
  assign n6001 = n6000 ^ n5997 ;
  assign n6002 = n5994 & n6001 ;
  assign n6003 = n6002 ^ n5999 ;
  assign n6004 = n6003 ^ n5997 ;
  assign n6005 = n5984 & ~n6004 ;
  assign n6006 = n6005 ^ n5984 ;
  assign n6007 = n6006 ^ x4 ;
  assign n6008 = n6007 ^ n6006 ;
  assign n6009 = n6008 ^ n5978 ;
  assign n6010 = ~x2 & n152 ;
  assign n6011 = ~n377 & ~n526 ;
  assign n6012 = ~x9 & n6011 ;
  assign n6013 = ~n623 & n6012 ;
  assign n6014 = ~n979 & ~n6013 ;
  assign n6015 = n6010 & ~n6014 ;
  assign n6016 = ~n433 & ~n434 ;
  assign n6017 = n100 & ~n6016 ;
  assign n6018 = n2039 & n5216 ;
  assign n6019 = ~n6017 & ~n6018 ;
  assign n6020 = n642 & n1192 ;
  assign n6021 = n99 & n6020 ;
  assign n6022 = ~n5918 & ~n6021 ;
  assign n6023 = n6019 & n6022 ;
  assign n6024 = ~n6015 & n6023 ;
  assign n6025 = n6024 ^ x5 ;
  assign n6026 = x5 & ~n6025 ;
  assign n6027 = n6026 ^ n6006 ;
  assign n6028 = n6027 ^ x5 ;
  assign n6029 = ~n6009 & ~n6028 ;
  assign n6030 = n6029 ^ n6026 ;
  assign n6031 = n6030 ^ x5 ;
  assign n6032 = n5978 & n6031 ;
  assign n6033 = n6032 ^ n5978 ;
  assign n6034 = ~n5971 & ~n6033 ;
  assign n6035 = x8 & ~n6034 ;
  assign n6036 = n434 & n5367 ;
  assign n6037 = n3779 & n6036 ;
  assign n6038 = n377 & n6037 ;
  assign n6039 = x14 & n6038 ;
  assign n6040 = n5217 ^ n21 ;
  assign n6041 = n6040 ^ n5217 ;
  assign n6042 = n5217 ^ n4162 ;
  assign n6043 = n6042 ^ n5217 ;
  assign n6044 = n6041 & n6043 ;
  assign n6045 = n6044 ^ n5217 ;
  assign n6046 = ~x2 & n6045 ;
  assign n6047 = n6046 ^ n5217 ;
  assign n6048 = n79 & n6047 ;
  assign n6049 = n431 & ~n1318 ;
  assign n6050 = ~n1808 & n6049 ;
  assign n6051 = n1141 & n5368 ;
  assign n6052 = n5365 & n6051 ;
  assign n6053 = ~n5100 & ~n6052 ;
  assign n6054 = ~n6050 & n6053 ;
  assign n6055 = n6054 ^ n1333 ;
  assign n6056 = n6055 ^ n6054 ;
  assign n6057 = n6054 ^ n1718 ;
  assign n6058 = n6057 ^ n6054 ;
  assign n6059 = n6056 & n6058 ;
  assign n6060 = n6059 ^ n6054 ;
  assign n6061 = ~x2 & ~n6060 ;
  assign n6062 = n6061 ^ n6054 ;
  assign n6063 = n642 & ~n6062 ;
  assign n6064 = ~n6048 & ~n6063 ;
  assign n6065 = ~x2 & n1959 ;
  assign n6066 = n1718 & ~n6065 ;
  assign n6067 = ~n323 & n405 ;
  assign n6068 = n6067 ^ n1364 ;
  assign n6069 = x4 & n6068 ;
  assign n6070 = n6069 ^ n1364 ;
  assign n6071 = n1255 & n6070 ;
  assign n6072 = n431 & n3684 ;
  assign n6073 = ~n6071 & ~n6072 ;
  assign n6074 = ~n6066 & n6073 ;
  assign n6075 = n167 & ~n6074 ;
  assign n6076 = n6064 & ~n6075 ;
  assign n6077 = n890 & ~n6076 ;
  assign n6078 = n560 & n1695 ;
  assign n6079 = n642 & ~n6078 ;
  assign n6080 = n1306 ^ x5 ;
  assign n6081 = n6080 ^ n1306 ;
  assign n6082 = n6081 ^ x4 ;
  assign n6083 = n1337 ^ n1306 ;
  assign n6084 = n6083 ^ n1306 ;
  assign n6085 = x2 & ~n405 ;
  assign n6086 = n6085 ^ x4 ;
  assign n6087 = ~n6084 & n6086 ;
  assign n6088 = n6087 ^ n6083 ;
  assign n6089 = n6088 ^ n6084 ;
  assign n6090 = ~n6082 & ~n6089 ;
  assign n6091 = n6090 ^ n6087 ;
  assign n6092 = x4 & n6091 ;
  assign n6093 = n6092 ^ x4 ;
  assign n6094 = n6079 & ~n6093 ;
  assign n6095 = n434 & ~n4911 ;
  assign n6096 = ~n305 & ~n1232 ;
  assign n6097 = n3889 & ~n6096 ;
  assign n6098 = ~x9 & ~n4908 ;
  assign n6099 = ~n6097 & n6098 ;
  assign n6100 = ~n6095 & ~n6099 ;
  assign n6101 = n3174 & n6100 ;
  assign n6102 = ~n6094 & n6101 ;
  assign n6103 = ~x8 & ~n6102 ;
  assign n6104 = ~x10 & n3626 ;
  assign n6105 = ~x12 & ~n1248 ;
  assign n6106 = n6104 & ~n6105 ;
  assign n6107 = n377 & ~n1054 ;
  assign n6108 = ~n1314 & ~n3684 ;
  assign n6109 = ~x13 & n432 ;
  assign n6110 = ~x5 & ~n6109 ;
  assign n6111 = ~n4167 & ~n6110 ;
  assign n6112 = n24 & ~n663 ;
  assign n6113 = ~x0 & ~n236 ;
  assign n6114 = ~n6112 & n6113 ;
  assign n6115 = ~n6111 & n6114 ;
  assign n6116 = n6108 & n6115 ;
  assign n6117 = ~n6107 & n6116 ;
  assign n6118 = ~n6106 & ~n6117 ;
  assign n6119 = n2434 & ~n6118 ;
  assign n6120 = x2 & ~x5 ;
  assign n6121 = ~n992 & ~n6120 ;
  assign n6122 = ~n24 & ~n6121 ;
  assign n6123 = n624 & n6122 ;
  assign n6124 = x9 & n6123 ;
  assign n6125 = ~n912 & n4132 ;
  assign n6126 = ~n377 & n6125 ;
  assign n6127 = n6126 ^ x0 ;
  assign n6128 = n6127 ^ n6126 ;
  assign n6129 = n6128 ^ n432 ;
  assign n6130 = n254 ^ x5 ;
  assign n6131 = ~n254 & ~n6130 ;
  assign n6132 = n6131 ^ n6126 ;
  assign n6133 = n6132 ^ n254 ;
  assign n6134 = n6129 & n6133 ;
  assign n6135 = n6134 ^ n6131 ;
  assign n6136 = n6135 ^ n254 ;
  assign n6137 = n432 & ~n6136 ;
  assign n6138 = n6137 ^ n432 ;
  assign n6139 = ~n6124 & ~n6138 ;
  assign n6140 = n2561 & ~n6139 ;
  assign n6141 = n3243 & ~n6120 ;
  assign n6142 = x10 & ~n1632 ;
  assign n6143 = n6141 & n6142 ;
  assign n6144 = ~n6140 & ~n6143 ;
  assign n6145 = n512 & n992 ;
  assign n6146 = n6145 ^ n6036 ;
  assign n6147 = x2 & n1831 ;
  assign n6148 = ~n3801 & ~n6147 ;
  assign n6149 = n6148 ^ n6145 ;
  assign n6150 = n6149 ^ n6148 ;
  assign n6151 = ~x4 & n434 ;
  assign n6152 = n4670 & n6151 ;
  assign n6153 = n6152 ^ n6148 ;
  assign n6154 = n6150 & n6153 ;
  assign n6155 = n6154 ^ n6148 ;
  assign n6156 = n6146 & n6155 ;
  assign n6157 = n6156 ^ n6036 ;
  assign n6158 = n6144 & ~n6157 ;
  assign n6159 = ~n6119 & n6158 ;
  assign n6160 = ~x7 & ~n6159 ;
  assign n6161 = n6103 & ~n6160 ;
  assign n6162 = ~n6077 & n6161 ;
  assign n6163 = ~n6039 & n6162 ;
  assign n6164 = ~n6035 & ~n6163 ;
  assign n6165 = n70 & n3521 ;
  assign n6166 = n1638 & n6165 ;
  assign n6167 = n604 & n708 ;
  assign n6168 = n4210 & n6167 ;
  assign n6169 = ~n6166 & ~n6168 ;
  assign n6170 = ~n6164 & n6169 ;
  assign n6171 = ~n5951 & n6170 ;
  assign n6172 = n1716 & ~n6171 ;
  assign n6173 = n6172 ^ n5948 ;
  assign n6174 = x5 ^ x2 ;
  assign n6175 = n344 & n1946 ;
  assign n6176 = ~n5318 & ~n6175 ;
  assign n6177 = n6176 ^ x5 ;
  assign n6178 = n6177 ^ n6176 ;
  assign n6179 = n362 & n1835 ;
  assign n6180 = n385 & n1960 ;
  assign n6181 = ~n6179 & ~n6180 ;
  assign n6182 = n6181 ^ n6176 ;
  assign n6183 = n6178 & n6182 ;
  assign n6184 = n6183 ^ n6176 ;
  assign n6185 = n6174 & ~n6184 ;
  assign n6186 = n658 & n6185 ;
  assign n6187 = ~n2530 & n4911 ;
  assign n6188 = n182 & n1705 ;
  assign n6189 = ~n6187 & ~n6188 ;
  assign n6190 = n25 & ~n6189 ;
  assign n6191 = n629 & n2817 ;
  assign n6192 = x4 & ~n591 ;
  assign n6193 = n813 & n6192 ;
  assign n6194 = ~n6191 & ~n6193 ;
  assign n6195 = n2039 & ~n6194 ;
  assign n6196 = ~n6190 & ~n6195 ;
  assign n6197 = ~n6186 & n6196 ;
  assign n6198 = n2682 & ~n6197 ;
  assign n6199 = n99 & n1835 ;
  assign n6200 = n1355 & n6199 ;
  assign n6201 = n6109 & n6200 ;
  assign n6202 = n3193 & n5880 ;
  assign n6203 = n1666 & ~n2440 ;
  assign n6204 = ~x11 & n6203 ;
  assign n6205 = ~n2406 & ~n6204 ;
  assign n6206 = n1808 & ~n6205 ;
  assign n6207 = ~n6202 & ~n6206 ;
  assign n6208 = n5042 & ~n6207 ;
  assign n6209 = ~x4 & n198 ;
  assign n6210 = n2781 & n6209 ;
  assign n6211 = ~n6208 & ~n6210 ;
  assign n6212 = ~n6201 & n6211 ;
  assign n6213 = n6212 ^ x0 ;
  assign n6214 = n6213 ^ n6212 ;
  assign n6215 = n1160 & n2817 ;
  assign n6216 = x9 & n6215 ;
  assign n6217 = n141 & n4907 ;
  assign n6218 = ~n3219 & n6217 ;
  assign n6219 = ~n1632 & n1939 ;
  assign n6220 = n137 & n6219 ;
  assign n6221 = n883 & n6220 ;
  assign n6222 = ~n6218 & ~n6221 ;
  assign n6223 = ~n6216 & n6222 ;
  assign n6224 = n60 & ~n6223 ;
  assign n6225 = ~n91 & n1865 ;
  assign n6226 = ~n1632 & n6225 ;
  assign n6227 = ~n4522 & ~n6226 ;
  assign n6228 = n51 & ~n6227 ;
  assign n6229 = n812 & n1898 ;
  assign n6230 = x11 & ~n6229 ;
  assign n6231 = ~n3068 & ~n6230 ;
  assign n6232 = ~n6228 & ~n6231 ;
  assign n6233 = n141 & n2040 ;
  assign n6234 = ~x11 & ~n6233 ;
  assign n6235 = n23 & ~n969 ;
  assign n6236 = ~n6234 & n6235 ;
  assign n6237 = ~n6232 & n6236 ;
  assign n6238 = ~n6224 & ~n6237 ;
  assign n6239 = n6238 ^ n6212 ;
  assign n6240 = ~n6214 & n6239 ;
  assign n6241 = n6240 ^ n6212 ;
  assign n6242 = ~n6198 & n6241 ;
  assign n6243 = n992 & ~n6242 ;
  assign n6244 = n1336 & n1960 ;
  assign n6245 = ~n1835 & ~n6244 ;
  assign n6246 = n3684 & ~n6245 ;
  assign n6247 = n2113 & n5418 ;
  assign n6248 = n3978 & n6247 ;
  assign n6249 = ~n6246 & ~n6248 ;
  assign n6250 = n2236 & ~n6249 ;
  assign n6251 = n2641 & n5189 ;
  assign n6252 = n2331 & n3876 ;
  assign n6253 = ~n6251 & ~n6252 ;
  assign n6254 = ~n6250 & n6253 ;
  assign n6255 = ~n1000 & ~n6254 ;
  assign n6256 = n764 & n3193 ;
  assign n6257 = n777 & n799 ;
  assign n6258 = ~n2043 & ~n6257 ;
  assign n6259 = n84 & ~n6258 ;
  assign n6260 = ~n6256 & ~n6259 ;
  assign n6261 = n3923 & ~n6260 ;
  assign n6262 = n1007 & n6233 ;
  assign n6263 = n142 & n1535 ;
  assign n6264 = ~n4255 & ~n6263 ;
  assign n6265 = x8 ^ x0 ;
  assign n6266 = n2789 & n6265 ;
  assign n6267 = n6266 ^ x0 ;
  assign n6268 = x4 & n6267 ;
  assign n6269 = ~n6264 & n6268 ;
  assign n6270 = ~n6262 & ~n6269 ;
  assign n6271 = ~n6261 & n6270 ;
  assign n6272 = x2 & ~n6271 ;
  assign n6273 = ~n6255 & ~n6272 ;
  assign n6274 = n859 & n1147 ;
  assign n6275 = n1101 & n6274 ;
  assign n6276 = n4210 & n6275 ;
  assign n6277 = ~n1207 & ~n5678 ;
  assign n6278 = ~n1808 & n2685 ;
  assign n6279 = ~n6277 & n6278 ;
  assign n6280 = n1718 & n2682 ;
  assign n6281 = ~n6279 & ~n6280 ;
  assign n6282 = n1112 & ~n6281 ;
  assign n6283 = n614 & n4210 ;
  assign n6284 = n988 & n6283 ;
  assign n6285 = ~n6282 & ~n6284 ;
  assign n6286 = n25 & ~n6285 ;
  assign n6287 = x7 & n529 ;
  assign n6288 = n2686 & n6287 ;
  assign n6289 = n1946 & n6120 ;
  assign n6290 = n6288 & n6289 ;
  assign n6291 = ~n6286 & ~n6290 ;
  assign n6445 = n753 & n2242 ;
  assign n6446 = ~n3572 & ~n6445 ;
  assign n6447 = n70 & n2704 ;
  assign n6448 = ~n998 & ~n6447 ;
  assign n6449 = n4260 & ~n6448 ;
  assign n6450 = ~n6446 & n6449 ;
  assign n6292 = n831 & n1351 ;
  assign n6293 = n141 & n3408 ;
  assign n6294 = n753 & n812 ;
  assign n6295 = n5567 & n6294 ;
  assign n6296 = ~n6293 & ~n6295 ;
  assign n6297 = ~n6292 & n6296 ;
  assign n6298 = n277 & ~n6297 ;
  assign n6299 = n2692 & n4726 ;
  assign n6300 = ~n125 & ~n5063 ;
  assign n6301 = n534 & ~n6300 ;
  assign n6302 = ~n91 & n6301 ;
  assign n6303 = ~n6299 & ~n6302 ;
  assign n6304 = x9 & ~n6303 ;
  assign n6305 = ~n6298 & ~n6304 ;
  assign n6306 = n5075 ^ n4044 ;
  assign n6307 = x7 ^ x3 ;
  assign n6308 = x7 ^ x5 ;
  assign n6309 = n6307 & n6308 ;
  assign n6310 = n6309 ^ x7 ;
  assign n6311 = n6310 ^ n4044 ;
  assign n6312 = n6306 & n6311 ;
  assign n6313 = n6312 ^ n6309 ;
  assign n6314 = n6313 ^ x7 ;
  assign n6315 = n6314 ^ n5075 ;
  assign n6316 = n4044 & n6315 ;
  assign n6317 = n6316 ^ n4044 ;
  assign n6318 = n6305 & ~n6317 ;
  assign n6319 = n1865 & ~n6318 ;
  assign n6320 = ~n1102 & n3685 ;
  assign n6321 = ~n99 & ~n230 ;
  assign n6322 = ~n100 & ~n281 ;
  assign n6323 = n6322 ^ n6321 ;
  assign n6324 = n3162 ^ x5 ;
  assign n6325 = n6324 ^ n3162 ;
  assign n6326 = n3582 & n6325 ;
  assign n6327 = n6326 ^ n3162 ;
  assign n6328 = n6327 ^ n6321 ;
  assign n6329 = n6323 & ~n6328 ;
  assign n6330 = n6329 ^ n6326 ;
  assign n6331 = n6330 ^ n3162 ;
  assign n6332 = n6331 ^ n6322 ;
  assign n6333 = ~n6321 & ~n6332 ;
  assign n6334 = n6333 ^ n6321 ;
  assign n6335 = ~n6320 & n6334 ;
  assign n6336 = ~x9 & ~n6335 ;
  assign n6337 = n663 & ~n5777 ;
  assign n6338 = n4336 & n6337 ;
  assign n6339 = n203 & n4744 ;
  assign n6340 = x7 & ~n6339 ;
  assign n6341 = n499 & n4726 ;
  assign n6342 = n6341 ^ n6339 ;
  assign n6343 = n6340 ^ n573 ;
  assign n6344 = n6342 & n6343 ;
  assign n6345 = n6344 ^ n573 ;
  assign n6346 = n6340 & n6345 ;
  assign n6347 = n6346 ^ n6339 ;
  assign n6348 = n1351 & n6347 ;
  assign n6349 = ~n6338 & ~n6348 ;
  assign n6350 = ~n6336 & n6349 ;
  assign n6351 = n1939 & ~n6350 ;
  assign n6352 = ~n6319 & ~n6351 ;
  assign n6353 = n988 & n1891 ;
  assign n6354 = n167 & ~n1198 ;
  assign n6355 = ~n6353 & ~n6354 ;
  assign n6356 = ~x0 & n6355 ;
  assign n6357 = ~n529 & n3408 ;
  assign n6358 = n60 & ~n6357 ;
  assign n6359 = n286 & n6358 ;
  assign n6360 = ~n6356 & n6359 ;
  assign n6361 = n658 & n1759 ;
  assign n6362 = ~n1698 & ~n6361 ;
  assign n6363 = n5585 & ~n6362 ;
  assign n6364 = n571 & ~n1198 ;
  assign n6365 = ~n3408 & ~n6364 ;
  assign n6366 = n614 & n3684 ;
  assign n6367 = ~n6365 & n6366 ;
  assign n6368 = ~n6363 & ~n6367 ;
  assign n6369 = ~n6360 & n6368 ;
  assign n6370 = n1835 & ~n6369 ;
  assign n6371 = n499 & n5924 ;
  assign n6372 = x2 & ~n743 ;
  assign n6373 = ~n604 & n6372 ;
  assign n6374 = ~n6371 & ~n6373 ;
  assign n6375 = n84 & ~n6374 ;
  assign n6376 = n1698 ^ n940 ;
  assign n6377 = n1698 ^ n106 ;
  assign n6378 = n6377 ^ n106 ;
  assign n6379 = ~x14 & ~n47 ;
  assign n6380 = n658 & ~n6379 ;
  assign n6381 = n6380 ^ n106 ;
  assign n6382 = ~n6378 & ~n6381 ;
  assign n6383 = n6382 ^ n106 ;
  assign n6384 = n6376 & n6383 ;
  assign n6385 = n6384 ^ n940 ;
  assign n6386 = ~n6375 & ~n6385 ;
  assign n6387 = n3923 & ~n6386 ;
  assign n6388 = n128 & n2719 ;
  assign n6389 = x5 & n6388 ;
  assign n6390 = ~n6387 & ~n6389 ;
  assign n6391 = ~n6370 & n6390 ;
  assign n6392 = n6352 & n6391 ;
  assign n6451 = n6450 ^ n6392 ;
  assign n6452 = n6451 ^ n6392 ;
  assign n6393 = n920 & ~n3144 ;
  assign n6396 = n3011 ^ x2 ;
  assign n6397 = n6396 ^ n3011 ;
  assign n6394 = n3011 ^ n281 ;
  assign n6395 = n6394 ^ n3011 ;
  assign n6398 = n6397 ^ n6395 ;
  assign n6399 = n3140 ^ n3011 ;
  assign n6400 = n6399 ^ n3011 ;
  assign n6401 = n6400 ^ n6397 ;
  assign n6402 = n6397 & ~n6401 ;
  assign n6403 = n6402 ^ n6397 ;
  assign n6404 = ~n6398 & n6403 ;
  assign n6405 = n6404 ^ n6402 ;
  assign n6406 = n6405 ^ n3011 ;
  assign n6407 = n6406 ^ n6397 ;
  assign n6408 = ~x0 & n6407 ;
  assign n6409 = n6408 ^ n3011 ;
  assign n6410 = ~n6393 & ~n6409 ;
  assign n6411 = n2242 & ~n6410 ;
  assign n6412 = n100 & n3627 ;
  assign n6413 = n1759 & n6412 ;
  assign n6414 = ~n1227 & ~n2440 ;
  assign n6415 = ~n2706 & ~n6414 ;
  assign n6416 = ~x0 & ~n6415 ;
  assign n6417 = n125 & ~n6104 ;
  assign n6418 = ~n6416 & n6417 ;
  assign n6419 = ~n6413 & ~n6418 ;
  assign n6420 = n2954 & ~n6419 ;
  assign n6421 = ~n499 & n1808 ;
  assign n6422 = n5979 & n6421 ;
  assign n6423 = ~x3 & ~n6422 ;
  assign n6424 = n753 & ~n1105 ;
  assign n6425 = ~n6423 & ~n6424 ;
  assign n6426 = ~n6420 & ~n6425 ;
  assign n6427 = ~n6411 & n6426 ;
  assign n6428 = ~x10 & n190 ;
  assign n6429 = n322 & n529 ;
  assign n6430 = n6428 & n6429 ;
  assign n6431 = ~n2696 & ~n6430 ;
  assign n6432 = n2198 & ~n6431 ;
  assign n6433 = n988 & n1698 ;
  assign n6434 = n5943 & n6433 ;
  assign n6435 = x3 & ~n6434 ;
  assign n6436 = ~n1000 & n2247 ;
  assign n6437 = n2682 & n5706 ;
  assign n6438 = ~n6436 & ~n6437 ;
  assign n6439 = x4 & ~n6438 ;
  assign n6440 = n6435 & ~n6439 ;
  assign n6441 = ~n6432 & n6440 ;
  assign n6442 = ~n6427 & ~n6441 ;
  assign n6443 = n6442 ^ n6392 ;
  assign n6444 = n6443 ^ n6392 ;
  assign n6453 = n6452 ^ n6444 ;
  assign n6454 = n230 & n659 ;
  assign n6455 = ~n2719 & ~n6454 ;
  assign n6456 = n84 & ~n6455 ;
  assign n6457 = ~n4005 & ~n4781 ;
  assign n6458 = ~x10 & ~n6457 ;
  assign n6459 = ~n126 & ~n6458 ;
  assign n6460 = n180 & ~n6459 ;
  assign n6461 = n556 & n1577 ;
  assign n6462 = n6109 & n6461 ;
  assign n6463 = ~n6460 & ~n6462 ;
  assign n6464 = ~n6456 & n6463 ;
  assign n6465 = n3154 & ~n6464 ;
  assign n6466 = n4167 & n4597 ;
  assign n6467 = ~x8 & n6466 ;
  assign n6468 = x0 & ~n6467 ;
  assign n6469 = ~n6262 & n6468 ;
  assign n6470 = ~n6465 & n6469 ;
  assign n6471 = x3 & n3781 ;
  assign n6472 = n4059 ^ x3 ;
  assign n6473 = n6472 ^ n4059 ;
  assign n6474 = n6473 ^ x14 ;
  assign n6475 = n432 ^ n205 ;
  assign n6476 = ~n432 & n6475 ;
  assign n6477 = n6476 ^ n4059 ;
  assign n6478 = n6477 ^ n432 ;
  assign n6479 = ~n6474 & ~n6478 ;
  assign n6480 = n6479 ^ n6476 ;
  assign n6481 = n6480 ^ n432 ;
  assign n6482 = x14 & ~n6481 ;
  assign n6483 = ~n6471 & ~n6482 ;
  assign n6484 = n86 & n2954 ;
  assign n6485 = ~n6483 & n6484 ;
  assign n6486 = n3154 & n5725 ;
  assign n6487 = ~n1535 & n5425 ;
  assign n6488 = ~n125 & n3590 ;
  assign n6489 = n6487 & n6488 ;
  assign n6490 = ~n6486 & ~n6489 ;
  assign n6491 = ~x13 & ~n6490 ;
  assign n6492 = x5 & ~n4162 ;
  assign n6493 = n5410 & ~n6492 ;
  assign n6494 = ~x0 & ~n6493 ;
  assign n6495 = ~n6491 & n6494 ;
  assign n6496 = ~n6485 & n6495 ;
  assign n6497 = ~x2 & ~n6496 ;
  assign n6498 = ~n6470 & n6497 ;
  assign n6499 = n6498 ^ n6392 ;
  assign n6500 = n6499 ^ n6392 ;
  assign n6501 = n6500 ^ n6452 ;
  assign n6502 = ~n6452 & n6501 ;
  assign n6503 = n6502 ^ n6452 ;
  assign n6504 = n6453 & ~n6503 ;
  assign n6505 = n6504 ^ n6502 ;
  assign n6506 = n6505 ^ n6392 ;
  assign n6507 = n6506 ^ n6452 ;
  assign n6508 = ~x11 & ~n6507 ;
  assign n6509 = n6508 ^ n6392 ;
  assign n6510 = n6291 & n6509 ;
  assign n6511 = ~n6276 & n6510 ;
  assign n6512 = n6511 ^ x12 ;
  assign n6513 = n6512 ^ n6511 ;
  assign n6514 = n3482 & n3488 ;
  assign n6515 = n2447 & n4349 ;
  assign n6516 = ~n6514 & ~n6515 ;
  assign n6517 = n3521 & ~n6516 ;
  assign n6518 = n2331 & n3510 ;
  assign n6519 = ~n6517 & ~n6518 ;
  assign n6520 = n281 & ~n6519 ;
  assign n6521 = n6520 ^ n6511 ;
  assign n6522 = ~n6513 & ~n6521 ;
  assign n6523 = n6522 ^ n6511 ;
  assign n6524 = n6273 & n6523 ;
  assign n6525 = ~n6243 & n6524 ;
  assign n6526 = n6525 ^ x6 ;
  assign n6527 = n6526 ^ n6525 ;
  assign n6528 = n442 & n4191 ;
  assign n6529 = n2943 & n6528 ;
  assign n6530 = ~n71 & ~n4910 ;
  assign n6531 = n4904 & ~n6530 ;
  assign n6532 = n100 & n5216 ;
  assign n6533 = n2136 & n6532 ;
  assign n6534 = ~n6531 & ~n6533 ;
  assign n6535 = n525 & ~n6534 ;
  assign n6536 = n1101 & n5075 ;
  assign n6537 = ~n4744 & ~n6536 ;
  assign n6538 = n1705 & n3308 ;
  assign n6539 = ~n6537 & n6538 ;
  assign n6540 = ~n6535 & ~n6539 ;
  assign n6541 = ~n6529 & n6540 ;
  assign n6542 = n560 & ~n6541 ;
  assign n6543 = n969 & n3228 ;
  assign n6544 = n556 & n4044 ;
  assign n6545 = n6543 & n6544 ;
  assign n6546 = ~n6542 & ~n6545 ;
  assign n6547 = n499 & n1808 ;
  assign n6548 = n2719 & n6547 ;
  assign n6549 = n431 & n6548 ;
  assign n6550 = n343 & n4191 ;
  assign n6551 = n202 & n431 ;
  assign n6552 = ~n277 & ~n6551 ;
  assign n6553 = n3626 & ~n6552 ;
  assign n6554 = x9 & ~n3219 ;
  assign n6555 = n2120 ^ x14 ;
  assign n6556 = n2120 ^ x7 ;
  assign n6557 = n6556 ^ x7 ;
  assign n6558 = n6557 ^ n6555 ;
  assign n6559 = n6555 ^ n1944 ;
  assign n6560 = ~x11 & ~n6559 ;
  assign n6561 = n6560 ^ x7 ;
  assign n6562 = ~n6558 & n6561 ;
  assign n6563 = n6562 ^ n6560 ;
  assign n6564 = ~n6555 & n6563 ;
  assign n6565 = n6564 ^ n6560 ;
  assign n6566 = n6565 ^ n6562 ;
  assign n6567 = n6566 ^ n2120 ;
  assign n6568 = n6554 & n6567 ;
  assign n6569 = n743 & n1376 ;
  assign n6570 = ~n712 & ~n6569 ;
  assign n6571 = ~n6568 & n6570 ;
  assign n6572 = ~x8 & ~n6571 ;
  assign n6573 = ~n4713 & ~n5702 ;
  assign n6574 = n913 & ~n6573 ;
  assign n6575 = ~n6572 & ~n6574 ;
  assign n6576 = ~x10 & ~n6575 ;
  assign n6577 = ~n6553 & ~n6576 ;
  assign n6578 = ~n6550 & n6577 ;
  assign n6579 = n5880 & ~n6578 ;
  assign n6580 = n442 & n2696 ;
  assign n6581 = ~x0 & ~n1000 ;
  assign n6582 = n605 & n2686 ;
  assign n6583 = ~n6581 & ~n6582 ;
  assign n6584 = n969 & ~n6583 ;
  assign n6585 = ~n1193 & n6584 ;
  assign n6586 = ~n6580 & ~n6585 ;
  assign n6587 = ~n3023 & ~n6586 ;
  assign n6588 = ~n416 & n624 ;
  assign n6589 = ~n277 & n6588 ;
  assign n6590 = ~n1014 & ~n6589 ;
  assign n6591 = n3578 & ~n6590 ;
  assign n6592 = ~n405 & n642 ;
  assign n6593 = n1101 & ~n6592 ;
  assign n6594 = n343 & n525 ;
  assign n6595 = n202 & ~n6594 ;
  assign n6596 = x0 & n6595 ;
  assign n6597 = ~n6593 & ~n6596 ;
  assign n6598 = n2242 & n6597 ;
  assign n6599 = x9 ^ x8 ;
  assign n6600 = n6599 ^ x8 ;
  assign n6601 = n3363 ^ x8 ;
  assign n6602 = ~n6600 & n6601 ;
  assign n6603 = n6602 ^ x8 ;
  assign n6604 = n743 & ~n6603 ;
  assign n6605 = n6598 & ~n6604 ;
  assign n6606 = ~n6591 & ~n6605 ;
  assign n6607 = n6606 ^ x2 ;
  assign n6608 = n6607 ^ n6606 ;
  assign n6609 = n105 & n2384 ;
  assign n6610 = n3154 & n6609 ;
  assign n6611 = ~n1872 & ~n1935 ;
  assign n6612 = n1400 & ~n6611 ;
  assign n6613 = n605 & n1252 ;
  assign n6614 = ~n2927 & ~n6613 ;
  assign n6615 = ~n5965 & n6614 ;
  assign n6616 = n3569 & ~n6615 ;
  assign n6617 = ~n6612 & ~n6616 ;
  assign n6618 = ~n6610 & n6617 ;
  assign n6619 = n624 & ~n6618 ;
  assign n6620 = ~n3897 & ~n5213 ;
  assign n6621 = ~x5 & ~n2652 ;
  assign n6622 = n2934 & ~n6621 ;
  assign n6623 = n6620 & n6622 ;
  assign n6624 = x0 & n105 ;
  assign n6625 = n6624 ^ x4 ;
  assign n6626 = n6625 ^ n6624 ;
  assign n6627 = n6626 ^ n6623 ;
  assign n6628 = n1505 ^ x9 ;
  assign n6629 = ~x9 & n6628 ;
  assign n6630 = n6629 ^ n6624 ;
  assign n6631 = n6630 ^ x9 ;
  assign n6632 = n6627 & n6631 ;
  assign n6633 = n6632 ^ n6629 ;
  assign n6634 = n6633 ^ x9 ;
  assign n6635 = n6623 & ~n6634 ;
  assign n6636 = n6635 ^ n6623 ;
  assign n6637 = ~n6619 & ~n6636 ;
  assign n6638 = n6637 ^ n6606 ;
  assign n6639 = ~n6608 & n6638 ;
  assign n6640 = n6639 ^ n6606 ;
  assign n6641 = ~n6587 & n6640 ;
  assign n6642 = ~n6579 & n6641 ;
  assign n6643 = x3 & ~n6642 ;
  assign n6644 = n443 & n993 ;
  assign n6645 = n534 & ~n1232 ;
  assign n6646 = ~n60 & ~n105 ;
  assign n6647 = n6645 & ~n6646 ;
  assign n6648 = x12 & n6647 ;
  assign n6649 = ~n6644 & ~n6648 ;
  assign n6650 = n1731 & ~n6649 ;
  assign n6651 = n1336 & n5367 ;
  assign n6652 = ~n404 & ~n6651 ;
  assign n6653 = n512 & ~n6652 ;
  assign n6654 = n1255 & n2298 ;
  assign n6655 = ~x0 & n6654 ;
  assign n6656 = ~n5028 & ~n6655 ;
  assign n6657 = ~n6653 & n6656 ;
  assign n6658 = n6657 ^ n4876 ;
  assign n6659 = n6658 ^ x9 ;
  assign n6666 = n6659 ^ n6658 ;
  assign n6660 = n6659 ^ n3263 ;
  assign n6661 = n6660 ^ n6658 ;
  assign n6662 = n6659 ^ n6657 ;
  assign n6663 = n6662 ^ n3263 ;
  assign n6664 = n6663 ^ n6661 ;
  assign n6665 = ~n6661 & n6664 ;
  assign n6667 = n6666 ^ n6665 ;
  assign n6668 = n6667 ^ n6661 ;
  assign n6669 = n6658 ^ x0 ;
  assign n6670 = n6665 ^ n6661 ;
  assign n6671 = ~n6669 & ~n6670 ;
  assign n6672 = n6671 ^ n6658 ;
  assign n6673 = ~n6668 & n6672 ;
  assign n6674 = n6673 ^ n6658 ;
  assign n6675 = n6674 ^ n4876 ;
  assign n6676 = n6675 ^ n6658 ;
  assign n6677 = n1011 & ~n6676 ;
  assign n6678 = ~n6650 & ~n6677 ;
  assign n6679 = n709 & n2685 ;
  assign n6680 = n2236 ^ x9 ;
  assign n6681 = n105 ^ x8 ;
  assign n6682 = n2236 ^ x8 ;
  assign n6683 = n6682 ^ x8 ;
  assign n6684 = ~n6681 & ~n6683 ;
  assign n6685 = n6684 ^ x8 ;
  assign n6686 = ~n6680 & n6685 ;
  assign n6687 = n6686 ^ x9 ;
  assign n6688 = ~x10 & ~n6687 ;
  assign n6689 = ~n6679 & ~n6688 ;
  assign n6690 = n1865 & ~n6689 ;
  assign n6691 = ~n6104 & ~n6151 ;
  assign n6692 = ~n2236 & ~n4490 ;
  assign n6693 = ~n6691 & ~n6692 ;
  assign n6694 = n989 & n2136 ;
  assign n6695 = ~n6693 & ~n6694 ;
  assign n6696 = n452 & ~n6695 ;
  assign n6697 = ~n6690 & ~n6696 ;
  assign n6698 = n2446 & ~n6697 ;
  assign n6699 = n4627 & n5213 ;
  assign n6700 = ~n614 & ~n6699 ;
  assign n6701 = n1054 & ~n6700 ;
  assign n6702 = x10 & n1233 ;
  assign n6703 = n3750 & n6702 ;
  assign n6704 = n124 & n963 ;
  assign n6705 = n199 & n253 ;
  assign n6706 = n1439 & n6705 ;
  assign n6707 = ~n6704 & ~n6706 ;
  assign n6708 = n3626 & ~n6707 ;
  assign n6709 = ~n6703 & ~n6708 ;
  assign n6710 = ~n6701 & n6709 ;
  assign n6711 = n2652 & ~n6710 ;
  assign n6712 = ~x2 & n1101 ;
  assign n6713 = n3406 & n6712 ;
  assign n6715 = n19 & ~n723 ;
  assign n6716 = n6715 ^ n642 ;
  assign n6724 = n6716 ^ n642 ;
  assign n6714 = n642 ^ n191 ;
  assign n6717 = n6716 ^ n6714 ;
  assign n6718 = n6717 ^ n6716 ;
  assign n6719 = n6718 ^ n642 ;
  assign n6720 = n6717 ^ x9 ;
  assign n6721 = n6720 ^ n6717 ;
  assign n6722 = n6721 ^ n6719 ;
  assign n6723 = n6719 & ~n6722 ;
  assign n6725 = n6724 ^ n6723 ;
  assign n6726 = n6725 ^ n6719 ;
  assign n6727 = n1944 ^ n642 ;
  assign n6728 = n6723 ^ n6719 ;
  assign n6729 = n6727 & n6728 ;
  assign n6730 = n6729 ^ n642 ;
  assign n6731 = n6726 & ~n6730 ;
  assign n6732 = n6731 ^ n642 ;
  assign n6733 = n6732 ^ n6715 ;
  assign n6734 = n6733 ^ n642 ;
  assign n6735 = n6713 & n6734 ;
  assign n6736 = x11 ^ x8 ;
  assign n6737 = n59 ^ x11 ;
  assign n6738 = n6737 ^ n59 ;
  assign n6739 = n1052 ^ n59 ;
  assign n6740 = n6738 & n6739 ;
  assign n6741 = n6740 ^ n59 ;
  assign n6742 = ~n6736 & n6741 ;
  assign n6743 = n2198 & n6742 ;
  assign n6744 = ~x9 & n6743 ;
  assign n6745 = ~n6735 & ~n6744 ;
  assign n6746 = n499 & n3355 ;
  assign n6747 = n990 & n6746 ;
  assign n6748 = n6745 & ~n6747 ;
  assign n6749 = ~n6711 & n6748 ;
  assign n6750 = ~n6698 & n6749 ;
  assign n6751 = n6678 & n6750 ;
  assign n6752 = n1705 & n3616 ;
  assign n6753 = ~n1695 & ~n6752 ;
  assign n6754 = n2236 & ~n6753 ;
  assign n6755 = n969 & n2120 ;
  assign n6756 = n362 ^ x14 ;
  assign n6757 = x14 ^ x12 ;
  assign n6758 = n6756 & n6757 ;
  assign n6759 = n6758 ^ x14 ;
  assign n6760 = n1933 & n6759 ;
  assign n6761 = ~n6755 & ~n6760 ;
  assign n6762 = ~x9 & ~n6761 ;
  assign n6763 = x2 & n5368 ;
  assign n6764 = ~n912 & n992 ;
  assign n6765 = ~n1705 & n3626 ;
  assign n6766 = n6764 & n6765 ;
  assign n6767 = ~n6763 & n6766 ;
  assign n6768 = ~n6543 & ~n6767 ;
  assign n6769 = ~n6762 & n6768 ;
  assign n6770 = ~n6754 & n6769 ;
  assign n6771 = n230 & ~n6770 ;
  assign n6772 = ~x7 & n6771 ;
  assign n6773 = n20 & n379 ;
  assign n6774 = n1336 & n6773 ;
  assign n6775 = x10 & n181 ;
  assign n6776 = ~n1959 & n6775 ;
  assign n6777 = n1336 & n1579 ;
  assign n6778 = ~n404 & ~n6777 ;
  assign n6779 = n203 & ~n6778 ;
  assign n6780 = ~n6776 & ~n6779 ;
  assign n6781 = ~n6774 & n6780 ;
  assign n6782 = n2136 & ~n6781 ;
  assign n6783 = ~n1193 & n4271 ;
  assign n6784 = ~n167 & ~n6783 ;
  assign n6785 = n3521 & ~n6784 ;
  assign n6786 = ~n2434 & n6592 ;
  assign n6787 = ~n1112 & ~n6786 ;
  assign n6788 = x0 & ~n4876 ;
  assign n6789 = ~n6787 & n6788 ;
  assign n6790 = ~n6785 & ~n6789 ;
  assign n6791 = ~n6782 & n6790 ;
  assign n6792 = n190 & ~n6791 ;
  assign n6793 = ~n6772 & ~n6792 ;
  assign n6794 = n6751 & n6793 ;
  assign n6795 = n142 & ~n6794 ;
  assign n6796 = ~n6643 & ~n6795 ;
  assign n6797 = ~n6549 & n6796 ;
  assign n6798 = n6546 & n6797 ;
  assign n6799 = n6798 ^ n6525 ;
  assign n6800 = n6527 & n6799 ;
  assign n6801 = n6800 ^ n6525 ;
  assign n6802 = n6801 ^ n5948 ;
  assign n6803 = ~n6173 & n6802 ;
  assign n6804 = n6803 ^ n6800 ;
  assign n6805 = n6804 ^ n6525 ;
  assign n6806 = n6805 ^ n6172 ;
  assign n6807 = n5948 & ~n6806 ;
  assign n6808 = n6807 ^ n5948 ;
  assign n6809 = ~n5912 & n6808 ;
  assign n6810 = n6809 ^ n5877 ;
  assign n6811 = n5879 & n6810 ;
  assign n6812 = n6811 ^ n5877 ;
  assign n6813 = n6812 ^ n4227 ;
  assign n6814 = ~n5409 & ~n6813 ;
  assign n6815 = n6814 ^ n6811 ;
  assign n6816 = n6815 ^ n5877 ;
  assign n6817 = n6816 ^ n5408 ;
  assign n6818 = ~n4227 & n6817 ;
  assign n6819 = n6818 ^ n4227 ;
  assign n6820 = n3714 & ~n6819 ;
  assign y0 = ~n6820 ;
endmodule
