module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 ;
  assign n9 = ~x0 & x4 ;
  assign n10 = x3 ^ x2 ;
  assign n11 = ~x6 & x7 ;
  assign n12 = n11 ^ x3 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = x6 & ~x7 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = ~n13 & n15 ;
  assign n17 = n16 ^ n11 ;
  assign n18 = ~n10 & n17 ;
  assign n19 = n9 & n18 ;
  assign n20 = x5 & n19 ;
  assign n26 = ~x6 & ~x7 ;
  assign n84 = ~x5 & n26 ;
  assign n85 = ~x3 & ~n84 ;
  assign n86 = ~x0 & ~n85 ;
  assign n87 = x2 & ~n86 ;
  assign n45 = x4 & x7 ;
  assign n46 = x5 & n45 ;
  assign n88 = x2 & x3 ;
  assign n21 = ~x4 & n11 ;
  assign n22 = x4 & ~x5 ;
  assign n30 = n14 & n22 ;
  assign n89 = ~n21 & ~n30 ;
  assign n90 = n88 & n89 ;
  assign n91 = ~n46 & n90 ;
  assign n92 = ~n87 & ~n91 ;
  assign n39 = x0 & ~x4 ;
  assign n93 = n26 ^ x3 ;
  assign n94 = n93 ^ n26 ;
  assign n95 = x6 & x7 ;
  assign n96 = x5 & n95 ;
  assign n97 = n96 ^ n26 ;
  assign n98 = ~n94 & n97 ;
  assign n99 = n98 ^ n26 ;
  assign n100 = n39 & n99 ;
  assign n101 = ~n92 & ~n100 ;
  assign n102 = ~x2 & x3 ;
  assign n48 = ~x4 & x6 ;
  assign n103 = n48 ^ n26 ;
  assign n104 = x5 & n103 ;
  assign n105 = n104 ^ n26 ;
  assign n106 = n105 ^ x0 ;
  assign n107 = n106 ^ n105 ;
  assign n108 = n107 ^ n102 ;
  assign n109 = n95 ^ x5 ;
  assign n110 = n95 & ~n109 ;
  assign n111 = n110 ^ n105 ;
  assign n112 = n111 ^ n95 ;
  assign n113 = n108 & n112 ;
  assign n114 = n113 ^ n110 ;
  assign n115 = n114 ^ n95 ;
  assign n116 = n102 & n115 ;
  assign n117 = n116 ^ n102 ;
  assign n118 = ~n101 & ~n117 ;
  assign n119 = ~x2 & ~x3 ;
  assign n120 = x6 ^ x5 ;
  assign n128 = n120 ^ x0 ;
  assign n122 = n120 ^ x7 ;
  assign n121 = n120 ^ x4 ;
  assign n123 = n122 ^ n121 ;
  assign n124 = n123 ^ x6 ;
  assign n125 = n124 ^ n120 ;
  assign n126 = n125 ^ x0 ;
  assign n135 = n126 ^ x0 ;
  assign n127 = n126 ^ n122 ;
  assign n136 = n135 ^ n127 ;
  assign n137 = n128 & n136 ;
  assign n129 = n123 ^ n122 ;
  assign n130 = n129 ^ n128 ;
  assign n131 = ~n127 & ~n130 ;
  assign n143 = n137 ^ n131 ;
  assign n132 = n131 ^ n126 ;
  assign n133 = n132 ^ n128 ;
  assign n134 = n133 ^ n127 ;
  assign n138 = n137 ^ n126 ;
  assign n139 = n138 ^ n128 ;
  assign n140 = n139 ^ n127 ;
  assign n141 = n140 ^ n119 ;
  assign n142 = n134 & n141 ;
  assign n144 = n143 ^ n142 ;
  assign n145 = n119 & n144 ;
  assign n146 = n145 ^ n119 ;
  assign n147 = n118 & ~n146 ;
  assign n38 = x5 & n26 ;
  assign n40 = n38 & n39 ;
  assign n41 = ~x3 & ~n40 ;
  assign n27 = n22 & n26 ;
  assign n23 = x6 & n22 ;
  assign n24 = ~n21 & ~n23 ;
  assign n25 = x2 & ~n24 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n28 ^ n27 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = ~n29 & ~n32 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = x0 & ~n34 ;
  assign n36 = n35 ^ n27 ;
  assign n37 = x3 & ~n36 ;
  assign n42 = n41 ^ n37 ;
  assign n43 = n37 ^ x2 ;
  assign n44 = n43 ^ n42 ;
  assign n53 = x0 & ~x5 ;
  assign n54 = n11 & n53 ;
  assign n55 = x4 ^ x0 ;
  assign n63 = n55 ^ x4 ;
  assign n64 = n63 ^ x4 ;
  assign n65 = ~n63 & n64 ;
  assign n56 = n55 ^ x5 ;
  assign n57 = n56 ^ x7 ;
  assign n58 = n57 ^ n56 ;
  assign n59 = n56 ^ n55 ;
  assign n60 = n59 ^ x4 ;
  assign n61 = ~n58 & ~n60 ;
  assign n68 = n65 ^ n61 ;
  assign n62 = n61 ^ x6 ;
  assign n66 = n65 ^ n63 ;
  assign n67 = ~n62 & ~n66 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = ~x6 & n69 ;
  assign n71 = n70 ^ n61 ;
  assign n72 = n71 ^ n65 ;
  assign n73 = n72 ^ n67 ;
  assign n74 = ~n54 & ~n73 ;
  assign n47 = x6 & n46 ;
  assign n49 = x5 & ~n48 ;
  assign n50 = ~n45 & n49 ;
  assign n51 = ~x0 & n50 ;
  assign n52 = ~n47 & ~n51 ;
  assign n75 = n74 ^ n52 ;
  assign n76 = x2 & n75 ;
  assign n77 = n76 ^ n52 ;
  assign n78 = n44 & n77 ;
  assign n79 = n78 ^ n76 ;
  assign n80 = n79 ^ n52 ;
  assign n81 = n80 ^ x2 ;
  assign n82 = n42 & n81 ;
  assign n83 = n82 ^ n41 ;
  assign n148 = n147 ^ n83 ;
  assign n149 = n148 ^ n147 ;
  assign n150 = ~x0 & n96 ;
  assign n151 = ~n27 & ~n150 ;
  assign n152 = ~n9 & n119 ;
  assign n153 = ~n151 & n152 ;
  assign n154 = n153 ^ n147 ;
  assign n155 = n154 ^ n147 ;
  assign n156 = n149 & ~n155 ;
  assign n157 = n156 ^ n147 ;
  assign n158 = x1 & ~n157 ;
  assign n159 = n158 ^ n147 ;
  assign n160 = ~n20 & ~n159 ;
  assign y0 = ~n160 ;
endmodule
