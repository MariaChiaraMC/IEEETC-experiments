module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 ;
  assign n23 = x0 & ~x2 ;
  assign n24 = ~x6 & ~x7 ;
  assign n25 = x5 & n24 ;
  assign n26 = n25 ^ x5 ;
  assign n27 = ~x4 & ~n26 ;
  assign n28 = n23 & ~n27 ;
  assign n30 = n28 ^ x3 ;
  assign n43 = n30 ^ n28 ;
  assign n10 = x3 ^ x2 ;
  assign n11 = x5 & x6 ;
  assign n12 = x7 & n11 ;
  assign n13 = x4 & n12 ;
  assign n14 = n13 ^ x2 ;
  assign n15 = ~n10 & ~n14 ;
  assign n16 = n15 ^ x2 ;
  assign n17 = ~x1 & x2 ;
  assign n18 = n17 ^ x0 ;
  assign n19 = n16 & ~n18 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = ~x0 & n20 ;
  assign n22 = n21 ^ x0 ;
  assign n29 = n28 ^ n22 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = n32 ^ n28 ;
  assign n34 = x4 & x5 ;
  assign n35 = ~x3 & ~n34 ;
  assign n36 = x0 & ~n35 ;
  assign n37 = x2 & ~n36 ;
  assign n38 = ~x1 & ~n37 ;
  assign n39 = n38 ^ n31 ;
  assign n40 = n39 ^ n31 ;
  assign n41 = n40 ^ n33 ;
  assign n42 = n33 & ~n41 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = n44 ^ n33 ;
  assign n50 = x4 ^ x2 ;
  assign n46 = ~x1 & ~n11 ;
  assign n47 = n46 ^ x0 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = n48 ^ n46 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = n48 ^ x2 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n51 & n53 ;
  assign n55 = n54 ^ n50 ;
  assign n56 = n50 ^ n48 ;
  assign n57 = n56 ^ n52 ;
  assign n62 = n52 ^ n49 ;
  assign n63 = ~x5 & n24 ;
  assign n64 = ~x8 & n63 ;
  assign n65 = n64 ^ n46 ;
  assign n66 = n62 & n65 ;
  assign n58 = x8 & n11 ;
  assign n59 = x7 & n58 ;
  assign n60 = n59 ^ n50 ;
  assign n61 = n56 & n60 ;
  assign n67 = n66 ^ n61 ;
  assign n68 = n67 ^ n46 ;
  assign n69 = n68 ^ n48 ;
  assign n70 = n69 ^ n52 ;
  assign n71 = n57 & n70 ;
  assign n72 = n71 ^ n61 ;
  assign n73 = n72 ^ n48 ;
  assign n74 = n73 ^ n52 ;
  assign n75 = n55 & n74 ;
  assign n76 = n75 ^ n61 ;
  assign n77 = n76 ^ n54 ;
  assign n78 = n77 ^ n71 ;
  assign n79 = n78 ^ n48 ;
  assign n80 = n79 ^ n50 ;
  assign n81 = n80 ^ n52 ;
  assign n82 = n81 ^ x0 ;
  assign n83 = n82 ^ n28 ;
  assign n84 = n42 ^ n33 ;
  assign n85 = n83 & n84 ;
  assign n86 = n85 ^ n28 ;
  assign n87 = n45 & ~n86 ;
  assign n88 = n87 ^ n28 ;
  assign n89 = n88 ^ x3 ;
  assign n90 = n89 ^ n28 ;
  assign y0 = n90 ;
endmodule
