module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 ;
  assign n8 = ~x4 & x5 ;
  assign n9 = n8 ^ x2 ;
  assign n10 = n9 ^ n8 ;
  assign n11 = x4 & ~x5 ;
  assign n12 = n11 ^ n8 ;
  assign n13 = n10 & n12 ;
  assign n14 = n13 ^ n8 ;
  assign n15 = ~x3 & n14 ;
  assign n31 = x5 ^ x4 ;
  assign n32 = n31 ^ x5 ;
  assign n37 = n32 ^ n31 ;
  assign n38 = n37 ^ x3 ;
  assign n39 = n38 ^ x3 ;
  assign n40 = n31 ^ x2 ;
  assign n41 = n40 ^ x3 ;
  assign n42 = ~n39 & ~n41 ;
  assign n33 = n31 ^ x6 ;
  assign n34 = n33 ^ n32 ;
  assign n35 = n34 ^ x3 ;
  assign n36 = n32 & n35 ;
  assign n43 = n42 ^ n36 ;
  assign n44 = n43 ^ n32 ;
  assign n45 = n36 ^ x3 ;
  assign n46 = n45 ^ n38 ;
  assign n47 = ~x3 & ~n46 ;
  assign n48 = n47 ^ n36 ;
  assign n49 = n44 & n48 ;
  assign n50 = n49 ^ n42 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = n51 ^ n32 ;
  assign n53 = n52 ^ x3 ;
  assign n54 = n53 ^ n38 ;
  assign n55 = ~x0 & ~n54 ;
  assign n16 = x2 ^ x0 ;
  assign n17 = n16 ^ x4 ;
  assign n18 = n17 ^ x2 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = n17 ^ x5 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = n19 & n21 ;
  assign n23 = n22 ^ n17 ;
  assign n24 = n23 ^ n19 ;
  assign n25 = n17 ^ x3 ;
  assign n26 = ~n18 & ~n25 ;
  assign n27 = n26 ^ n17 ;
  assign n28 = ~n24 & ~n27 ;
  assign n29 = n28 ^ n17 ;
  assign n30 = n29 ^ n16 ;
  assign n56 = n55 ^ n30 ;
  assign n57 = n56 ^ n30 ;
  assign n58 = ~x3 & ~x4 ;
  assign n59 = x0 & n58 ;
  assign n60 = x4 & x5 ;
  assign n61 = x2 & n60 ;
  assign n62 = ~n59 & ~n61 ;
  assign n63 = n62 ^ n30 ;
  assign n64 = n63 ^ n30 ;
  assign n65 = ~n57 & n64 ;
  assign n66 = n65 ^ n30 ;
  assign n67 = ~x1 & n66 ;
  assign n68 = n67 ^ n30 ;
  assign n69 = ~n15 & n68 ;
  assign y0 = ~n69 ;
endmodule
