module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 ;
  assign n9 = ~x5 & ~x6 ;
  assign n10 = x4 ^ x3 ;
  assign n11 = x7 ^ x4 ;
  assign n12 = ~n10 & ~n11 ;
  assign n13 = n12 ^ x4 ;
  assign n14 = n9 & n13 ;
  assign n15 = x3 ^ x2 ;
  assign n16 = n15 ^ x6 ;
  assign n17 = n16 ^ x7 ;
  assign n18 = ~x3 & ~n17 ;
  assign n19 = x6 ^ x3 ;
  assign n20 = x7 ^ x3 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n19 & ~n21 ;
  assign n23 = n22 ^ x5 ;
  assign n24 = n18 & n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = x5 & n25 ;
  assign n27 = n26 ^ n15 ;
  assign n28 = n27 ^ x4 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ n14 ;
  assign n31 = ~x2 & x6 ;
  assign n32 = n31 ^ x5 ;
  assign n33 = x5 & n32 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = n34 ^ x5 ;
  assign n36 = ~n30 & ~n35 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ x5 ;
  assign n39 = ~n14 & n38 ;
  assign n40 = n39 ^ n14 ;
  assign n41 = ~x1 & n40 ;
  assign n42 = x5 & x6 ;
  assign n43 = ~x4 & ~n42 ;
  assign n44 = x1 & ~n43 ;
  assign n45 = x4 & ~x7 ;
  assign n46 = x5 & n45 ;
  assign n47 = ~x3 & ~n46 ;
  assign n48 = ~n44 & n47 ;
  assign n49 = x6 ^ x1 ;
  assign n50 = x7 ^ x1 ;
  assign n51 = n50 ^ x1 ;
  assign n52 = ~n49 & n51 ;
  assign n53 = n52 ^ x1 ;
  assign n54 = x4 & x5 ;
  assign n55 = x1 & ~n54 ;
  assign n56 = n55 ^ x3 ;
  assign n57 = n53 & n56 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = x3 & n58 ;
  assign n60 = n59 ^ x3 ;
  assign n61 = ~n48 & ~n60 ;
  assign n62 = ~x2 & n61 ;
  assign n63 = ~n41 & ~n62 ;
  assign n64 = ~x0 & ~n63 ;
  assign y0 = n64 ;
endmodule
