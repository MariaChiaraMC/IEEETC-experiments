module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 ;
  assign n41 = x7 & x8 ;
  assign n42 = ~x4 & ~n41 ;
  assign n43 = x5 & ~n42 ;
  assign n10 = ~x4 & ~x5 ;
  assign n11 = ~x6 & ~n10 ;
  assign n12 = ~x5 & x8 ;
  assign n13 = n11 & n12 ;
  assign n14 = ~x4 & x6 ;
  assign n15 = n14 ^ x3 ;
  assign n16 = x5 & n15 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = ~x7 & ~x8 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n14 & n19 ;
  assign n21 = n20 ^ n14 ;
  assign n22 = n21 ^ x3 ;
  assign n23 = n17 & n22 ;
  assign n24 = ~n13 & ~n23 ;
  assign n25 = ~x2 & ~n24 ;
  assign n26 = x6 ^ x4 ;
  assign n27 = x0 & x3 ;
  assign n28 = n27 ^ x6 ;
  assign n29 = n27 ^ x5 ;
  assign n30 = ~n27 & n29 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n28 & ~n31 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = n34 ^ x5 ;
  assign n36 = ~n26 & n35 ;
  assign n37 = n18 & n36 ;
  assign n38 = ~n25 & ~n37 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = n44 ^ n38 ;
  assign n39 = n38 ^ x2 ;
  assign n40 = n39 ^ n38 ;
  assign n46 = n45 ^ n40 ;
  assign n47 = n10 ^ x6 ;
  assign n48 = n10 & ~n18 ;
  assign n49 = n47 & n48 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = n50 ^ n38 ;
  assign n52 = n51 ^ n38 ;
  assign n53 = n52 ^ n45 ;
  assign n54 = ~n45 & n53 ;
  assign n55 = n54 ^ n45 ;
  assign n56 = ~n46 & ~n55 ;
  assign n57 = n56 ^ n54 ;
  assign n58 = n57 ^ n38 ;
  assign n59 = n58 ^ n45 ;
  assign n60 = x1 & n59 ;
  assign n61 = n60 ^ n38 ;
  assign y0 = ~n61 ;
endmodule
