module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 ;
  assign n22 = x1 ^ x0 ;
  assign n23 = x2 ^ x1 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = x5 ^ x3 ;
  assign n27 = x5 ^ x1 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = ~n26 & ~n28 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = n30 ^ n26 ;
  assign n32 = n25 & ~n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ n26 ;
  assign n35 = n22 & ~n34 ;
  assign n36 = ~x4 & n35 ;
  assign n37 = ~x19 & ~x20 ;
  assign n38 = n37 ^ x18 ;
  assign n39 = n38 ^ x18 ;
  assign n40 = x1 & x13 ;
  assign n41 = ~x0 & x1 ;
  assign n42 = x4 & ~n41 ;
  assign n43 = ~n40 & n42 ;
  assign n44 = ~x9 & ~x10 ;
  assign n45 = x11 ^ x8 ;
  assign n46 = ~x7 & x16 ;
  assign n47 = x11 & n46 ;
  assign n48 = n45 & n47 ;
  assign n49 = n48 ^ n45 ;
  assign n50 = n44 & n49 ;
  assign n51 = ~x6 & ~x17 ;
  assign n55 = ~x8 & x9 ;
  assign n56 = ~x11 & n55 ;
  assign n52 = ~x11 & x12 ;
  assign n53 = x13 & ~n52 ;
  assign n54 = x8 & ~n53 ;
  assign n57 = n56 ^ n54 ;
  assign n58 = n56 ^ x10 ;
  assign n59 = n58 ^ n56 ;
  assign n60 = n59 ^ n51 ;
  assign n61 = n60 ^ x17 ;
  assign n62 = n57 & n61 ;
  assign n63 = n62 ^ n56 ;
  assign n64 = n51 & n63 ;
  assign n65 = n64 ^ n51 ;
  assign n66 = x10 & ~x13 ;
  assign n67 = ~n52 & ~n66 ;
  assign n68 = n67 ^ x15 ;
  assign n69 = n68 ^ x9 ;
  assign n70 = ~x9 & n69 ;
  assign n71 = n70 ^ x15 ;
  assign n72 = n71 ^ x9 ;
  assign n73 = x11 & ~x12 ;
  assign n74 = n73 ^ x15 ;
  assign n75 = ~x13 & ~n74 ;
  assign n76 = n75 ^ x15 ;
  assign n77 = n72 & ~n76 ;
  assign n78 = n77 ^ x15 ;
  assign n79 = n78 ^ x15 ;
  assign n80 = n65 & n79 ;
  assign n81 = ~n50 & n80 ;
  assign n82 = n81 ^ x2 ;
  assign n83 = n82 ^ n81 ;
  assign n84 = x13 ^ x12 ;
  assign n85 = n84 ^ x12 ;
  assign n86 = x12 ^ x10 ;
  assign n87 = n85 & n86 ;
  assign n88 = n87 ^ x10 ;
  assign n89 = x12 ^ x9 ;
  assign n90 = n89 ^ n84 ;
  assign n91 = n90 ^ n73 ;
  assign n92 = n91 ^ n90 ;
  assign n93 = n90 ^ n84 ;
  assign n94 = n93 ^ x12 ;
  assign n95 = n94 ^ n87 ;
  assign n96 = n92 & n95 ;
  assign n97 = n96 ^ n56 ;
  assign n98 = ~x10 & n97 ;
  assign n99 = n98 ^ n96 ;
  assign n100 = n99 ^ n85 ;
  assign n101 = ~n88 & n100 ;
  assign n102 = n101 ^ n96 ;
  assign n103 = n102 ^ n98 ;
  assign n104 = n103 ^ n85 ;
  assign n105 = n104 ^ x13 ;
  assign n106 = n105 ^ n81 ;
  assign n107 = ~n83 & ~n106 ;
  assign n108 = n107 ^ n81 ;
  assign n109 = n43 & n108 ;
  assign n110 = x5 & ~n109 ;
  assign n111 = x0 & ~x1 ;
  assign n112 = n111 ^ x4 ;
  assign n113 = n112 ^ n111 ;
  assign n114 = ~x0 & ~x2 ;
  assign n115 = n114 ^ n111 ;
  assign n116 = ~n113 & n115 ;
  assign n117 = n116 ^ n111 ;
  assign n118 = ~x10 & x11 ;
  assign n119 = ~x8 & ~x9 ;
  assign n120 = n118 & n119 ;
  assign n121 = x2 & n120 ;
  assign n122 = n111 & n121 ;
  assign n123 = n122 ^ n110 ;
  assign n124 = n117 & ~n123 ;
  assign n125 = n124 ^ n122 ;
  assign n126 = ~n110 & n125 ;
  assign n127 = n126 ^ n110 ;
  assign n128 = ~x3 & n127 ;
  assign n129 = ~x0 & ~x1 ;
  assign n130 = ~x9 & ~n129 ;
  assign n131 = ~x1 & x3 ;
  assign n132 = ~x2 & n131 ;
  assign n133 = ~n114 & ~n132 ;
  assign n134 = ~n130 & ~n133 ;
  assign n135 = ~x5 & ~n134 ;
  assign n136 = ~x6 & ~x7 ;
  assign n137 = ~x12 & n136 ;
  assign n138 = ~x13 & ~n137 ;
  assign n139 = ~x8 & ~n138 ;
  assign n140 = n44 ^ x11 ;
  assign n141 = n44 ^ x5 ;
  assign n142 = n141 ^ x5 ;
  assign n143 = x13 ^ x5 ;
  assign n144 = ~n142 & ~n143 ;
  assign n145 = n144 ^ x5 ;
  assign n146 = ~n140 & n145 ;
  assign n147 = n139 & n146 ;
  assign n148 = ~n135 & n147 ;
  assign n149 = ~x12 & ~x13 ;
  assign n150 = ~x2 & x5 ;
  assign n151 = n118 & n136 ;
  assign n152 = ~n114 & ~n131 ;
  assign n153 = n151 & ~n152 ;
  assign n154 = x10 & ~x11 ;
  assign n155 = ~x5 & ~n132 ;
  assign n156 = n154 & ~n155 ;
  assign n157 = ~n153 & ~n156 ;
  assign n158 = x8 & ~n157 ;
  assign n159 = ~n150 & ~n158 ;
  assign n160 = n149 & ~n159 ;
  assign n161 = x9 & n160 ;
  assign n162 = ~n148 & ~n161 ;
  assign n163 = ~x4 & ~n162 ;
  assign n164 = x3 & ~x5 ;
  assign n165 = n164 ^ x4 ;
  assign n166 = n165 ^ n164 ;
  assign n167 = ~x3 & n149 ;
  assign n168 = x2 & n167 ;
  assign n170 = ~x8 & ~x11 ;
  assign n171 = ~n44 & n170 ;
  assign n173 = n171 ^ n136 ;
  assign n182 = n173 ^ n171 ;
  assign n169 = x8 & x9 ;
  assign n172 = n171 ^ n169 ;
  assign n174 = n173 ^ n172 ;
  assign n175 = n174 ^ n173 ;
  assign n176 = n175 ^ n171 ;
  assign n177 = n174 ^ x10 ;
  assign n178 = n177 ^ x11 ;
  assign n179 = n178 ^ n174 ;
  assign n180 = n179 ^ n176 ;
  assign n181 = n176 & n180 ;
  assign n183 = n182 ^ n181 ;
  assign n184 = n183 ^ n176 ;
  assign n185 = n171 ^ x11 ;
  assign n186 = n181 ^ n176 ;
  assign n187 = n185 & n186 ;
  assign n188 = n187 ^ n171 ;
  assign n189 = n184 & ~n188 ;
  assign n190 = n189 ^ n171 ;
  assign n191 = n190 ^ n136 ;
  assign n192 = n191 ^ n171 ;
  assign n193 = n168 & n192 ;
  assign n194 = n193 ^ n164 ;
  assign n195 = ~n166 & n194 ;
  assign n196 = n195 ^ n164 ;
  assign n197 = ~n129 & n196 ;
  assign n198 = x5 ^ x2 ;
  assign n199 = n198 ^ n23 ;
  assign n201 = n55 & n73 ;
  assign n202 = ~x3 & ~n201 ;
  assign n200 = ~x0 & x4 ;
  assign n203 = n202 ^ n200 ;
  assign n204 = x2 & n203 ;
  assign n205 = n204 ^ n202 ;
  assign n206 = ~n199 & ~n205 ;
  assign n207 = n206 ^ n204 ;
  assign n208 = n207 ^ n202 ;
  assign n209 = n208 ^ x2 ;
  assign n210 = ~n23 & ~n209 ;
  assign n211 = ~n197 & ~n210 ;
  assign n212 = ~n163 & n211 ;
  assign n213 = ~n128 & n212 ;
  assign n214 = n213 ^ x18 ;
  assign n215 = n39 & n214 ;
  assign n216 = n215 ^ x18 ;
  assign n217 = x14 & n216 ;
  assign n218 = ~n36 & n217 ;
  assign y0 = ~n218 ;
endmodule
