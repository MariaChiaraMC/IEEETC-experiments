module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 ;
  assign n9 = x1 & ~x3 ;
  assign n10 = ~x5 & ~x6 ;
  assign n11 = ~x0 & n10 ;
  assign n12 = n9 & n11 ;
  assign n54 = ~x6 & x7 ;
  assign n22 = x0 & x3 ;
  assign n55 = ~x1 & n22 ;
  assign n56 = x0 & n9 ;
  assign n57 = n56 ^ x5 ;
  assign n58 = n57 ^ n56 ;
  assign n17 = ~x1 & ~x3 ;
  assign n59 = n56 ^ n17 ;
  assign n60 = ~n58 & n59 ;
  assign n61 = n60 ^ n56 ;
  assign n62 = ~n55 & ~n61 ;
  assign n63 = n54 & ~n62 ;
  assign n18 = x5 & x6 ;
  assign n64 = x1 & x3 ;
  assign n65 = n18 & n64 ;
  assign n66 = x3 & ~n10 ;
  assign n67 = ~x3 & ~x6 ;
  assign n68 = ~x1 & ~x7 ;
  assign n69 = ~n67 & n68 ;
  assign n70 = ~n66 & n69 ;
  assign n71 = ~n65 & ~n70 ;
  assign n72 = ~x0 & ~n71 ;
  assign n73 = x1 & x6 ;
  assign n74 = x5 ^ x3 ;
  assign n75 = n74 ^ x6 ;
  assign n39 = ~x0 & x5 ;
  assign n76 = n73 ^ n39 ;
  assign n77 = n75 & n76 ;
  assign n78 = n77 ^ n39 ;
  assign n79 = n73 & n78 ;
  assign n80 = x7 & n79 ;
  assign n81 = ~n72 & ~n80 ;
  assign n82 = ~n63 & n81 ;
  assign n13 = x0 & ~x5 ;
  assign n14 = ~x6 & ~x7 ;
  assign n15 = ~x3 & n14 ;
  assign n16 = n13 & n15 ;
  assign n19 = n17 & n18 ;
  assign n20 = n19 ^ x1 ;
  assign n21 = n20 ^ x7 ;
  assign n32 = n21 ^ n20 ;
  assign n23 = ~x5 & x7 ;
  assign n24 = x6 & n23 ;
  assign n25 = n22 & n24 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = n26 ^ n20 ;
  assign n28 = n21 ^ n19 ;
  assign n29 = n28 ^ n25 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = ~n27 & ~n30 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = x6 ^ x3 ;
  assign n36 = n35 ^ n13 ;
  assign n37 = n13 ^ x6 ;
  assign n38 = n37 ^ x6 ;
  assign n40 = n39 ^ x6 ;
  assign n41 = ~n38 & n40 ;
  assign n42 = n41 ^ x6 ;
  assign n43 = n36 & n42 ;
  assign n44 = n43 ^ n13 ;
  assign n45 = n44 ^ n20 ;
  assign n46 = n31 ^ n27 ;
  assign n47 = ~n45 & ~n46 ;
  assign n48 = n47 ^ n20 ;
  assign n49 = ~n34 & n48 ;
  assign n50 = n49 ^ n20 ;
  assign n51 = n50 ^ x1 ;
  assign n52 = n51 ^ n20 ;
  assign n53 = ~n16 & ~n52 ;
  assign n83 = n82 ^ n53 ;
  assign n84 = ~x2 & n83 ;
  assign n85 = n84 ^ n82 ;
  assign n86 = ~n12 & n85 ;
  assign n87 = ~x4 & ~n86 ;
  assign n88 = x6 ^ x5 ;
  assign n89 = x7 ^ x1 ;
  assign n90 = n89 ^ x6 ;
  assign n91 = n90 ^ x1 ;
  assign n92 = n9 ^ x1 ;
  assign n93 = n91 & ~n92 ;
  assign n94 = n93 ^ x1 ;
  assign n95 = n88 & ~n94 ;
  assign n96 = n95 ^ n9 ;
  assign n97 = n96 ^ n95 ;
  assign n98 = x5 & n14 ;
  assign n99 = n98 ^ n95 ;
  assign n100 = n99 ^ n95 ;
  assign n101 = n97 & n100 ;
  assign n102 = n101 ^ n95 ;
  assign n103 = x0 & n102 ;
  assign n104 = n103 ^ n95 ;
  assign n105 = n104 ^ x2 ;
  assign n106 = n105 ^ n104 ;
  assign n107 = x5 & ~n54 ;
  assign n108 = n55 & n107 ;
  assign n109 = x6 ^ x1 ;
  assign n110 = x7 ^ x3 ;
  assign n111 = n110 ^ x7 ;
  assign n112 = x7 ^ x6 ;
  assign n113 = n112 ^ x7 ;
  assign n114 = n111 & n113 ;
  assign n115 = n114 ^ x7 ;
  assign n116 = ~n109 & n115 ;
  assign n117 = n116 ^ x0 ;
  assign n118 = n117 ^ n116 ;
  assign n119 = n54 & n64 ;
  assign n120 = x6 & n17 ;
  assign n121 = ~n119 & ~n120 ;
  assign n122 = n121 ^ n116 ;
  assign n123 = ~n118 & ~n122 ;
  assign n124 = n123 ^ n116 ;
  assign n125 = ~x5 & n124 ;
  assign n126 = ~n108 & ~n125 ;
  assign n127 = n126 ^ n104 ;
  assign n128 = ~n106 & ~n127 ;
  assign n129 = n128 ^ n104 ;
  assign n130 = x4 & n129 ;
  assign n131 = n12 ^ x2 ;
  assign n132 = n131 ^ n12 ;
  assign n133 = n18 & n55 ;
  assign n134 = n133 ^ n12 ;
  assign n135 = n132 & n134 ;
  assign n136 = n135 ^ n12 ;
  assign n137 = ~x7 & n136 ;
  assign n138 = ~n130 & ~n137 ;
  assign n139 = ~n87 & n138 ;
  assign y0 = ~n139 ;
endmodule
