module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 ;
  assign n9 = ~x1 & ~x5 ;
  assign n10 = ~x4 & ~n9 ;
  assign n11 = x5 ^ x2 ;
  assign n12 = x6 ^ x5 ;
  assign n13 = n12 ^ x6 ;
  assign n14 = ~x1 & x7 ;
  assign n15 = x3 & ~x6 ;
  assign n16 = ~n14 & ~n15 ;
  assign n17 = n16 ^ x6 ;
  assign n18 = n13 & ~n17 ;
  assign n19 = n18 ^ x6 ;
  assign n20 = ~n11 & n19 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = n10 & ~n21 ;
  assign n23 = ~x0 & ~n22 ;
  assign n24 = x6 & ~n10 ;
  assign n25 = x5 ^ x3 ;
  assign n26 = ~x1 & ~n25 ;
  assign n27 = n26 ^ x3 ;
  assign n28 = n24 & n27 ;
  assign n29 = x5 ^ x4 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n29 ^ x1 ;
  assign n33 = n31 & n32 ;
  assign n34 = n33 ^ n29 ;
  assign n35 = ~x2 & x6 ;
  assign n36 = ~n29 & ~n35 ;
  assign n37 = n36 ^ n25 ;
  assign n38 = ~n34 & n37 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n25 & n39 ;
  assign n41 = n40 ^ x3 ;
  assign n42 = n41 ^ n25 ;
  assign n43 = ~n28 & n42 ;
  assign n44 = n23 & n43 ;
  assign y0 = n44 ;
endmodule
