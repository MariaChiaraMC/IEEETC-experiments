// Benchmark "./pla/m1.pla_1" written by ABC on Mon Apr 20 15:44:06 2020

module \./pla/m1.pla_1  ( 
    x0, x1, x2, x3, x4, x5,
    z0  );
  input  x0, x1, x2, x3, x4, x5;
  output z0;
  assign z0 = ~x0;
endmodule


