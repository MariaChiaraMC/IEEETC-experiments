module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n10 = x7 ^ x0 ;
  assign n11 = ~x2 & x6 ;
  assign n12 = n11 ^ x7 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = ~x1 & ~x2 ;
  assign n15 = ~x3 & x5 ;
  assign n16 = n14 & n15 ;
  assign n17 = n16 ^ n11 ;
  assign n18 = n17 ^ n10 ;
  assign n19 = ~n13 & n18 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = ~x4 & ~x8 ;
  assign n22 = n16 & n21 ;
  assign n23 = n22 ^ n10 ;
  assign n24 = n20 & ~n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = ~n10 & n25 ;
  assign n27 = n26 ^ n19 ;
  assign n28 = n27 ^ n16 ;
  assign y0 = n28 ;
endmodule
