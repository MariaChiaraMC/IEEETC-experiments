module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 ;
  assign n10 = ~x7 & ~x8 ;
  assign n11 = x6 & ~n10 ;
  assign n12 = ~x3 & x5 ;
  assign n13 = ~x0 & x1 ;
  assign n14 = ~n12 & n13 ;
  assign n15 = x2 & x3 ;
  assign n16 = n15 ^ x5 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = x5 ^ x1 ;
  assign n19 = n18 ^ x5 ;
  assign n20 = n17 & ~n19 ;
  assign n21 = n20 ^ x5 ;
  assign n22 = x4 & ~n21 ;
  assign n23 = n22 ^ x5 ;
  assign n24 = ~n14 & n23 ;
  assign n25 = ~n11 & ~n24 ;
  assign y0 = n25 ;
endmodule
