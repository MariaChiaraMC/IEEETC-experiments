module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 ;
  assign n10 = x1 ^ x0 ;
  assign n11 = ~x2 & ~x3 ;
  assign n12 = ~x4 & ~x6 ;
  assign n13 = x7 & x8 ;
  assign n14 = n12 & n13 ;
  assign n15 = x6 ^ x4 ;
  assign n16 = n15 ^ x8 ;
  assign n17 = n16 ^ x6 ;
  assign n18 = n17 ^ x8 ;
  assign n20 = n18 ^ x5 ;
  assign n21 = n20 ^ n16 ;
  assign n34 = n21 ^ n16 ;
  assign n23 = n18 ^ x7 ;
  assign n24 = n23 ^ x5 ;
  assign n28 = n24 ^ x5 ;
  assign n29 = n28 ^ n18 ;
  assign n30 = n29 ^ x0 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n35 ^ n21 ;
  assign n32 = n30 ^ x0 ;
  assign n40 = n36 ^ n32 ;
  assign n41 = n30 ^ n21 ;
  assign n19 = n18 ^ x0 ;
  assign n42 = n41 ^ n19 ;
  assign n43 = n40 & ~n42 ;
  assign n22 = n16 ^ x8 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n26 ^ n21 ;
  assign n31 = n30 ^ n27 ;
  assign n33 = n32 ^ n31 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n37 ^ n19 ;
  assign n39 = n19 & ~n38 ;
  assign n44 = n43 ^ n39 ;
  assign n45 = n44 ^ n21 ;
  assign n46 = n45 ^ n30 ;
  assign n47 = n46 ^ n32 ;
  assign n48 = n47 ^ n19 ;
  assign n49 = n39 ^ n21 ;
  assign n50 = n49 ^ n30 ;
  assign n51 = n32 ^ n30 ;
  assign n52 = n51 ^ n19 ;
  assign n53 = n32 ^ n21 ;
  assign n54 = n53 ^ n36 ;
  assign n55 = ~n52 & ~n54 ;
  assign n56 = n55 ^ n32 ;
  assign n57 = n56 ^ n36 ;
  assign n58 = n57 ^ n19 ;
  assign n59 = ~n50 & n58 ;
  assign n60 = n59 ^ n30 ;
  assign n61 = n48 & n60 ;
  assign n62 = n61 ^ n55 ;
  assign n63 = n62 ^ n43 ;
  assign n64 = n63 ^ n59 ;
  assign n65 = n64 ^ n21 ;
  assign n66 = n65 ^ n35 ;
  assign n67 = ~n14 & ~n66 ;
  assign n68 = n11 & ~n67 ;
  assign n69 = n68 ^ n10 ;
  assign n70 = n69 ^ x1 ;
  assign n71 = n70 ^ n69 ;
  assign n72 = x3 & ~x5 ;
  assign n73 = ~n13 & ~n72 ;
  assign n74 = x2 & x3 ;
  assign n75 = x1 & x6 ;
  assign n76 = ~n74 & n75 ;
  assign n77 = ~n73 & n76 ;
  assign n78 = x3 & x5 ;
  assign n79 = ~x6 & x7 ;
  assign n80 = x2 & n79 ;
  assign n81 = n78 & n80 ;
  assign n82 = x8 & n81 ;
  assign n83 = n82 ^ n77 ;
  assign n84 = ~x7 & x8 ;
  assign n85 = n84 ^ n79 ;
  assign n86 = ~x2 & n85 ;
  assign n87 = n86 ^ n79 ;
  assign n88 = n72 & n87 ;
  assign n89 = x2 & n84 ;
  assign n90 = x1 & n89 ;
  assign n91 = ~x3 & ~x6 ;
  assign n92 = n91 ^ x3 ;
  assign n93 = ~x5 & n92 ;
  assign n94 = n93 ^ x3 ;
  assign n95 = n90 & n94 ;
  assign n96 = ~x5 & ~x7 ;
  assign n97 = x2 & ~n91 ;
  assign n98 = n96 & n97 ;
  assign n99 = x5 & x7 ;
  assign n100 = ~n11 & ~n99 ;
  assign n101 = ~x6 & ~n100 ;
  assign n102 = ~n98 & ~n101 ;
  assign n103 = x1 & ~n102 ;
  assign n104 = x7 & n11 ;
  assign n105 = x6 ^ x3 ;
  assign n106 = n105 ^ x2 ;
  assign n107 = n106 ^ n105 ;
  assign n108 = n107 ^ n104 ;
  assign n109 = x3 & ~x7 ;
  assign n110 = n109 ^ x6 ;
  assign n111 = n109 & ~n110 ;
  assign n112 = n111 ^ n105 ;
  assign n113 = n112 ^ n109 ;
  assign n114 = n108 & ~n113 ;
  assign n115 = n114 ^ n111 ;
  assign n116 = n115 ^ n109 ;
  assign n117 = ~n104 & n116 ;
  assign n118 = n117 ^ n104 ;
  assign n119 = x5 & n118 ;
  assign n120 = ~n103 & ~n119 ;
  assign n121 = ~x8 & ~n120 ;
  assign n122 = ~n95 & ~n121 ;
  assign n123 = ~n88 & n122 ;
  assign n124 = n123 ^ x4 ;
  assign n125 = n124 ^ n123 ;
  assign n126 = ~x2 & ~x6 ;
  assign n127 = ~n109 & n126 ;
  assign n128 = ~x8 & ~n97 ;
  assign n129 = ~n127 & n128 ;
  assign n130 = ~x5 & n129 ;
  assign n132 = x3 & x6 ;
  assign n131 = x7 & ~x8 ;
  assign n133 = n132 ^ n131 ;
  assign n134 = n133 ^ n131 ;
  assign n135 = n134 ^ n130 ;
  assign n136 = x2 & x5 ;
  assign n137 = ~n78 & ~n136 ;
  assign n138 = ~x6 & ~n84 ;
  assign n139 = n138 ^ n137 ;
  assign n140 = ~n137 & n139 ;
  assign n141 = n140 ^ n131 ;
  assign n142 = n141 ^ n137 ;
  assign n143 = n135 & ~n142 ;
  assign n144 = n143 ^ n140 ;
  assign n145 = n144 ^ n137 ;
  assign n146 = ~n130 & ~n145 ;
  assign n147 = n146 ^ n130 ;
  assign n148 = x1 & n147 ;
  assign n162 = x3 & n89 ;
  assign n149 = n109 ^ n13 ;
  assign n150 = n149 ^ x3 ;
  assign n151 = n150 ^ n13 ;
  assign n152 = n13 & n151 ;
  assign n153 = n152 ^ n149 ;
  assign n154 = n153 ^ n13 ;
  assign n155 = n149 ^ x2 ;
  assign n156 = n155 ^ n13 ;
  assign n157 = x5 & ~n156 ;
  assign n158 = n157 ^ n149 ;
  assign n159 = n154 & n158 ;
  assign n160 = n159 ^ n149 ;
  assign n161 = n160 ^ n109 ;
  assign n163 = n162 ^ n161 ;
  assign n164 = ~x6 & n163 ;
  assign n165 = n164 ^ n161 ;
  assign n166 = ~n148 & ~n165 ;
  assign n167 = n166 ^ n123 ;
  assign n168 = ~n125 & n167 ;
  assign n169 = n168 ^ n123 ;
  assign n170 = n169 ^ n77 ;
  assign n171 = n83 & ~n170 ;
  assign n172 = n171 ^ n168 ;
  assign n173 = n172 ^ n123 ;
  assign n174 = n173 ^ n82 ;
  assign n175 = ~n77 & ~n174 ;
  assign n176 = n175 ^ n77 ;
  assign n177 = n176 ^ n69 ;
  assign n178 = n177 ^ n10 ;
  assign n179 = ~n71 & ~n178 ;
  assign n180 = n179 ^ n176 ;
  assign n181 = ~n12 & ~n99 ;
  assign n182 = ~n96 & ~n181 ;
  assign n183 = n182 ^ x2 ;
  assign n184 = n183 ^ n182 ;
  assign n185 = ~x5 & x8 ;
  assign n186 = ~x4 & n185 ;
  assign n187 = ~x6 & ~x7 ;
  assign n188 = ~x8 & n187 ;
  assign n189 = ~n186 & ~n188 ;
  assign n190 = n189 ^ n182 ;
  assign n191 = n184 & ~n190 ;
  assign n192 = n191 ^ n182 ;
  assign n193 = ~x3 & n192 ;
  assign n194 = n12 & n78 ;
  assign n195 = x8 ^ x5 ;
  assign n196 = n195 ^ x8 ;
  assign n197 = x6 & x8 ;
  assign n198 = n197 ^ x8 ;
  assign n199 = n196 & ~n198 ;
  assign n200 = n199 ^ x8 ;
  assign n201 = x4 & ~n200 ;
  assign n202 = ~n194 & ~n201 ;
  assign n203 = x7 & ~n202 ;
  assign n204 = ~x8 & n72 ;
  assign n205 = ~n186 & ~n204 ;
  assign n206 = x6 & ~n205 ;
  assign n207 = ~n203 & ~n206 ;
  assign n208 = x2 & ~n207 ;
  assign n209 = n208 ^ n193 ;
  assign n210 = n72 & n84 ;
  assign n211 = x6 & ~x8 ;
  assign n212 = n109 & n211 ;
  assign n213 = ~n210 & ~n212 ;
  assign n214 = n213 ^ x4 ;
  assign n215 = n214 ^ n213 ;
  assign n216 = n79 & n185 ;
  assign n217 = n211 ^ n84 ;
  assign n218 = ~x2 & n217 ;
  assign n219 = n218 ^ n84 ;
  assign n220 = x5 & n219 ;
  assign n221 = ~x3 & n220 ;
  assign n222 = ~n216 & ~n221 ;
  assign n223 = n222 ^ n213 ;
  assign n224 = n215 & n223 ;
  assign n225 = n224 ^ n213 ;
  assign n226 = n225 ^ n193 ;
  assign n227 = n209 & ~n226 ;
  assign n228 = n227 ^ n224 ;
  assign n229 = n228 ^ n213 ;
  assign n230 = n229 ^ n208 ;
  assign n231 = ~n193 & ~n230 ;
  assign n232 = n231 ^ n193 ;
  assign n233 = ~n176 & ~n232 ;
  assign n234 = n233 ^ n10 ;
  assign n235 = ~n180 & ~n234 ;
  assign n236 = n235 ^ n233 ;
  assign n237 = ~n10 & n236 ;
  assign n238 = n237 ^ n179 ;
  assign n239 = n238 ^ x0 ;
  assign n240 = n239 ^ n176 ;
  assign y0 = n240 ;
endmodule
