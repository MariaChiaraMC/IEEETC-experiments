module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 ;
  assign n16 = ~x4 & ~x5 ;
  assign n17 = ~x11 & x12 ;
  assign n18 = x13 & x14 ;
  assign n19 = ~x6 & x8 ;
  assign n20 = n18 & n19 ;
  assign n21 = n17 & n20 ;
  assign n22 = x11 & ~x13 ;
  assign n23 = ~x12 & n22 ;
  assign n24 = ~x0 & n23 ;
  assign n25 = ~x6 & ~x8 ;
  assign n26 = x9 & ~n25 ;
  assign n27 = n24 & n26 ;
  assign n28 = ~n21 & ~n27 ;
  assign n29 = n16 & ~n28 ;
  assign n30 = n29 ^ x9 ;
  assign n31 = n30 ^ x7 ;
  assign n96 = n31 ^ n30 ;
  assign n35 = ~x1 & ~x6 ;
  assign n33 = ~x12 & x14 ;
  assign n34 = x4 & n33 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = n34 ^ x11 ;
  assign n38 = n37 ^ x11 ;
  assign n39 = x11 & x12 ;
  assign n40 = ~x2 & n39 ;
  assign n41 = n40 ^ x11 ;
  assign n42 = ~n38 & ~n41 ;
  assign n43 = n42 ^ x11 ;
  assign n44 = ~n36 & n43 ;
  assign n45 = n44 ^ n35 ;
  assign n46 = x5 & ~n45 ;
  assign n32 = x13 ^ x4 ;
  assign n47 = n46 ^ n32 ;
  assign n48 = n47 ^ x13 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = n49 ^ n32 ;
  assign n52 = x7 & ~x14 ;
  assign n53 = x12 & ~x13 ;
  assign n54 = n52 & ~n53 ;
  assign n55 = x12 ^ x11 ;
  assign n56 = x1 & ~n55 ;
  assign n57 = n54 & n56 ;
  assign n58 = ~x5 & n57 ;
  assign n51 = n47 ^ n32 ;
  assign n59 = n58 ^ n51 ;
  assign n60 = ~n50 & ~n59 ;
  assign n61 = n60 ^ n58 ;
  assign n65 = ~x11 & ~x12 ;
  assign n66 = x5 & ~x7 ;
  assign n67 = n65 & ~n66 ;
  assign n62 = n32 ^ x14 ;
  assign n63 = n62 ^ n51 ;
  assign n64 = n63 ^ n49 ;
  assign n68 = n67 ^ n64 ;
  assign n69 = n62 ^ n58 ;
  assign n70 = ~n68 & ~n69 ;
  assign n71 = n70 ^ n62 ;
  assign n72 = n71 ^ n49 ;
  assign n73 = n72 ^ n67 ;
  assign n74 = n62 ^ n49 ;
  assign n75 = n63 ^ n58 ;
  assign n76 = n75 ^ n50 ;
  assign n77 = ~n74 & ~n76 ;
  assign n78 = n77 ^ n51 ;
  assign n79 = n78 ^ n49 ;
  assign n80 = n79 ^ n58 ;
  assign n81 = n73 & ~n80 ;
  assign n82 = n81 ^ n49 ;
  assign n83 = n82 ^ n50 ;
  assign n84 = n61 & ~n83 ;
  assign n85 = n84 ^ n81 ;
  assign n86 = n85 ^ n49 ;
  assign n87 = n86 ^ n50 ;
  assign n88 = n87 ^ x4 ;
  assign n89 = ~x0 & ~n88 ;
  assign n90 = n89 ^ n31 ;
  assign n91 = n90 ^ n30 ;
  assign n92 = n31 ^ n29 ;
  assign n93 = n92 ^ n89 ;
  assign n94 = n93 ^ n91 ;
  assign n95 = n91 & n94 ;
  assign n97 = n96 ^ n95 ;
  assign n98 = n97 ^ n91 ;
  assign n99 = x4 & n65 ;
  assign n100 = x5 & x6 ;
  assign n101 = ~x13 & ~x14 ;
  assign n102 = ~n18 & ~n101 ;
  assign n103 = n100 & ~n102 ;
  assign n104 = n99 & n103 ;
  assign n105 = n16 & n19 ;
  assign n106 = n101 & n105 ;
  assign n107 = x11 & n106 ;
  assign n108 = ~n104 & ~n107 ;
  assign n109 = n108 ^ n30 ;
  assign n110 = n95 ^ n91 ;
  assign n111 = ~n109 & n110 ;
  assign n112 = n111 ^ n30 ;
  assign n113 = ~n98 & ~n112 ;
  assign n114 = n113 ^ n30 ;
  assign n115 = n114 ^ x9 ;
  assign n116 = n115 ^ n30 ;
  assign n117 = x10 & ~n116 ;
  assign n118 = n25 & n53 ;
  assign n119 = x7 & ~x9 ;
  assign n120 = ~x11 & x14 ;
  assign n121 = n119 & n120 ;
  assign n122 = n16 & n121 ;
  assign n123 = n118 & n122 ;
  assign n124 = ~n117 & ~n123 ;
  assign n125 = x3 & ~n124 ;
  assign n129 = ~x9 & ~n120 ;
  assign n130 = x3 & ~x13 ;
  assign n131 = ~n52 & ~n130 ;
  assign n132 = ~n129 & n131 ;
  assign n133 = n17 & ~n132 ;
  assign n134 = ~x7 & x8 ;
  assign n135 = x6 & n134 ;
  assign n136 = n135 ^ x12 ;
  assign n137 = n135 ^ x13 ;
  assign n138 = n137 ^ x13 ;
  assign n139 = n16 & n130 ;
  assign n140 = n139 ^ x13 ;
  assign n141 = n138 & n140 ;
  assign n142 = n141 ^ x13 ;
  assign n143 = n136 & n142 ;
  assign n144 = n143 ^ x12 ;
  assign n145 = ~x11 & ~n144 ;
  assign n146 = n23 ^ x14 ;
  assign n147 = n146 ^ x0 ;
  assign n156 = n147 ^ n146 ;
  assign n148 = ~x1 & n23 ;
  assign n149 = n148 ^ n22 ;
  assign n150 = n149 ^ n147 ;
  assign n151 = n150 ^ n146 ;
  assign n152 = n147 ^ n23 ;
  assign n153 = n152 ^ n149 ;
  assign n154 = n153 ^ n151 ;
  assign n155 = n151 & ~n154 ;
  assign n157 = n156 ^ n155 ;
  assign n158 = n157 ^ n151 ;
  assign n159 = n146 ^ n65 ;
  assign n160 = n155 ^ n151 ;
  assign n161 = ~n159 & n160 ;
  assign n162 = n161 ^ n146 ;
  assign n163 = ~n158 & n162 ;
  assign n164 = n163 ^ n146 ;
  assign n165 = n164 ^ x14 ;
  assign n166 = n165 ^ n146 ;
  assign n167 = ~n145 & ~n166 ;
  assign n168 = n167 ^ x9 ;
  assign n176 = n168 ^ n120 ;
  assign n177 = ~x9 & n176 ;
  assign n169 = x12 ^ x9 ;
  assign n170 = n169 ^ n168 ;
  assign n171 = n170 ^ x3 ;
  assign n172 = n171 ^ n170 ;
  assign n173 = n170 ^ n168 ;
  assign n174 = n173 ^ x9 ;
  assign n175 = ~n172 & ~n174 ;
  assign n178 = n177 ^ n175 ;
  assign n179 = n178 ^ n168 ;
  assign n180 = n177 ^ n168 ;
  assign n126 = ~x4 & ~x9 ;
  assign n181 = ~x13 & n126 ;
  assign n182 = n181 ^ n170 ;
  assign n183 = n182 ^ n168 ;
  assign n184 = n183 ^ n175 ;
  assign n185 = n184 ^ n172 ;
  assign n186 = n180 & n185 ;
  assign n187 = n186 ^ x9 ;
  assign n188 = n179 & ~n187 ;
  assign n189 = n188 ^ n177 ;
  assign n190 = n189 ^ n186 ;
  assign n191 = n190 ^ n167 ;
  assign n192 = ~n133 & ~n191 ;
  assign n127 = n53 & n126 ;
  assign n128 = x11 & n127 ;
  assign n193 = n192 ^ n128 ;
  assign n194 = x10 & ~n193 ;
  assign n195 = n194 ^ n192 ;
  assign n196 = ~n125 & n195 ;
  assign y0 = ~n196 ;
endmodule
