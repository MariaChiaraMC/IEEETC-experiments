module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 ;
  assign n53 = x1 & ~x4 ;
  assign n24 = x5 & ~x6 ;
  assign n54 = x2 & n24 ;
  assign n55 = n53 & n54 ;
  assign n9 = ~x4 & x5 ;
  assign n56 = x1 & ~x2 ;
  assign n57 = x3 & ~x6 ;
  assign n58 = n56 & n57 ;
  assign n59 = ~n9 & n58 ;
  assign n60 = ~n55 & ~n59 ;
  assign n61 = ~x0 & ~n60 ;
  assign n10 = ~x4 & x6 ;
  assign n62 = ~x0 & ~n10 ;
  assign n63 = x3 & x4 ;
  assign n64 = ~x1 & x2 ;
  assign n65 = ~n63 & n64 ;
  assign n66 = n62 & n65 ;
  assign n67 = ~x3 & x6 ;
  assign n68 = n56 & n67 ;
  assign n69 = ~x4 & n68 ;
  assign n70 = ~n66 & ~n69 ;
  assign n71 = ~x5 & ~n70 ;
  assign n72 = x5 & x6 ;
  assign n73 = x3 & n72 ;
  assign n74 = ~x4 & ~n73 ;
  assign n19 = x4 & x5 ;
  assign n20 = x0 & ~n19 ;
  assign n39 = x4 & ~x6 ;
  assign n75 = ~x2 & ~n39 ;
  assign n76 = x1 & ~n75 ;
  assign n77 = n20 & n76 ;
  assign n78 = ~n74 & n77 ;
  assign n79 = ~n71 & ~n78 ;
  assign n80 = ~n61 & n79 ;
  assign n81 = n24 & n63 ;
  assign n82 = n64 & n81 ;
  assign n83 = x0 & ~x3 ;
  assign n13 = x1 & ~x5 ;
  assign n84 = n13 ^ x2 ;
  assign n85 = n84 ^ n13 ;
  assign n86 = ~x5 & n10 ;
  assign n87 = ~x1 & x4 ;
  assign n88 = n24 & n87 ;
  assign n89 = ~n86 & ~n88 ;
  assign n90 = n89 ^ n13 ;
  assign n91 = ~n85 & ~n90 ;
  assign n92 = n91 ^ n13 ;
  assign n93 = n83 & n92 ;
  assign n94 = ~n82 & ~n93 ;
  assign n95 = ~x7 & n94 ;
  assign n96 = n80 & n95 ;
  assign n34 = x4 & ~x5 ;
  assign n35 = ~n9 & ~n34 ;
  assign n11 = ~n9 & ~n10 ;
  assign n12 = ~x0 & ~n11 ;
  assign n14 = x6 & ~n13 ;
  assign n15 = n12 & ~n14 ;
  assign n16 = x1 & x6 ;
  assign n17 = ~x0 & ~n16 ;
  assign n18 = ~n10 & n17 ;
  assign n21 = x6 & n20 ;
  assign n22 = ~n18 & ~n21 ;
  assign n23 = x1 & x5 ;
  assign n25 = ~n23 & ~n24 ;
  assign n26 = x4 ^ x1 ;
  assign n27 = ~x6 & ~n26 ;
  assign n28 = n25 & ~n27 ;
  assign n29 = x7 & n28 ;
  assign n30 = n22 & n29 ;
  assign n31 = ~n15 & ~n30 ;
  assign n36 = n35 ^ n31 ;
  assign n37 = n36 ^ n31 ;
  assign n32 = n31 ^ x0 ;
  assign n33 = n32 ^ n31 ;
  assign n38 = n37 ^ n33 ;
  assign n40 = ~n16 & ~n39 ;
  assign n41 = x7 & n40 ;
  assign n42 = n41 ^ n31 ;
  assign n43 = n42 ^ n31 ;
  assign n44 = n43 ^ n37 ;
  assign n45 = ~n37 & ~n44 ;
  assign n46 = n45 ^ n37 ;
  assign n47 = ~n38 & ~n46 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = n48 ^ n31 ;
  assign n50 = n49 ^ n37 ;
  assign n51 = ~x3 & n50 ;
  assign n52 = n51 ^ n31 ;
  assign n97 = n96 ^ n52 ;
  assign n98 = n97 ^ x2 ;
  assign n109 = n98 ^ n97 ;
  assign n99 = x0 & x3 ;
  assign n100 = n86 & n99 ;
  assign n101 = ~x1 & n100 ;
  assign n102 = x7 & ~n101 ;
  assign n103 = n102 ^ n98 ;
  assign n104 = n103 ^ n97 ;
  assign n105 = n102 ^ n96 ;
  assign n106 = n105 ^ n102 ;
  assign n107 = n106 ^ n104 ;
  assign n108 = n104 & ~n107 ;
  assign n110 = n109 ^ n108 ;
  assign n111 = n110 ^ n104 ;
  assign n112 = x6 ^ x3 ;
  assign n113 = n112 ^ x4 ;
  assign n114 = n113 ^ x6 ;
  assign n115 = n114 ^ n113 ;
  assign n116 = n112 ^ x0 ;
  assign n117 = n116 ^ x1 ;
  assign n118 = n117 ^ x5 ;
  assign n119 = n118 ^ n113 ;
  assign n120 = n119 ^ n112 ;
  assign n121 = n120 ^ n115 ;
  assign n122 = n115 & n121 ;
  assign n123 = n122 ^ n113 ;
  assign n124 = n123 ^ n115 ;
  assign n126 = x5 ^ x1 ;
  assign n125 = n118 ^ x1 ;
  assign n127 = n126 ^ n125 ;
  assign n128 = n127 ^ n126 ;
  assign n129 = n128 ^ n120 ;
  assign n131 = n128 ^ n113 ;
  assign n132 = n131 ^ n112 ;
  assign n133 = n129 & n132 ;
  assign n130 = n120 & n129 ;
  assign n134 = n133 ^ n130 ;
  assign n135 = n134 ^ n126 ;
  assign n136 = n135 ^ n128 ;
  assign n137 = n136 ^ n113 ;
  assign n138 = n137 ^ n120 ;
  assign n139 = ~n112 & n138 ;
  assign n140 = n139 ^ n130 ;
  assign n141 = n140 ^ n126 ;
  assign n142 = n141 ^ n120 ;
  assign n143 = ~n124 & ~n142 ;
  assign n144 = n143 ^ n122 ;
  assign n145 = n144 ^ n126 ;
  assign n146 = n145 ^ n113 ;
  assign n147 = n146 ^ n115 ;
  assign n148 = n147 ^ n126 ;
  assign n149 = n148 ^ n97 ;
  assign n150 = n108 ^ n104 ;
  assign n151 = n149 & n150 ;
  assign n152 = n151 ^ n97 ;
  assign n153 = n111 & n152 ;
  assign n154 = n153 ^ n97 ;
  assign n155 = n154 ^ n96 ;
  assign n156 = n155 ^ n97 ;
  assign y0 = ~n156 ;
endmodule
