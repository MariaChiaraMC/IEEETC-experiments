module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n11 = x8 ^ x1 ;
  assign n12 = n11 ^ x4 ;
  assign n13 = x7 ^ x5 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = x8 ^ x5 ;
  assign n16 = n14 & n15 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = n17 ^ n11 ;
  assign n19 = n12 & n18 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = n20 ^ x5 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = ~n11 & n22 ;
  assign n24 = n23 ^ n11 ;
  assign y0 = n24 ;
endmodule
