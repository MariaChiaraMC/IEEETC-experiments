module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 ;
  assign n17 = x9 & x15 ;
  assign n18 = x12 & ~x14 ;
  assign n19 = ~x11 & ~n18 ;
  assign n20 = x13 & ~n19 ;
  assign n21 = x2 ^ x0 ;
  assign n22 = n21 ^ x1 ;
  assign n23 = x7 ^ x3 ;
  assign n24 = x3 ^ x2 ;
  assign n25 = n24 ^ x3 ;
  assign n26 = ~n23 & n25 ;
  assign n27 = n26 ^ x3 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = ~n22 & ~n28 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n30 ^ x3 ;
  assign n32 = n31 ^ x1 ;
  assign n33 = n21 & n32 ;
  assign n34 = n33 ^ n21 ;
  assign n35 = ~n20 & n34 ;
  assign n36 = x11 & x13 ;
  assign n37 = x12 & n36 ;
  assign n38 = x15 & ~n37 ;
  assign n39 = ~x14 & n37 ;
  assign n40 = n39 ^ x2 ;
  assign n41 = x3 & ~x6 ;
  assign n42 = n41 ^ x1 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = ~x0 & x7 ;
  assign n45 = x8 & n44 ;
  assign n46 = n45 ^ n41 ;
  assign n47 = n43 & n46 ;
  assign n48 = n47 ^ n41 ;
  assign n49 = n48 ^ n39 ;
  assign n50 = n40 & ~n49 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = n51 ^ n41 ;
  assign n53 = n52 ^ x2 ;
  assign n54 = ~n39 & ~n53 ;
  assign n55 = n54 ^ n39 ;
  assign n56 = ~n38 & ~n55 ;
  assign n57 = ~n35 & ~n56 ;
  assign n58 = x4 & x10 ;
  assign n59 = ~x5 & n58 ;
  assign n60 = ~n57 & n59 ;
  assign n61 = ~n17 & ~n60 ;
  assign y0 = ~n61 ;
endmodule
