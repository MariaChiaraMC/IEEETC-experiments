module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n11 = ~x6 & x9 ;
  assign n12 = ~x0 & ~x7 ;
  assign n13 = ~x3 & n12 ;
  assign n14 = ~n11 & ~n13 ;
  assign n15 = ~x0 & ~x8 ;
  assign n16 = x7 & ~n15 ;
  assign n17 = ~x2 & ~x4 ;
  assign n18 = ~n16 & n17 ;
  assign n19 = ~n14 & n18 ;
  assign n20 = ~x1 & ~x5 ;
  assign n21 = n12 ^ x3 ;
  assign n22 = n21 ^ n12 ;
  assign n23 = ~x7 & ~x8 ;
  assign n24 = x6 & ~x9 ;
  assign n25 = n12 & ~n24 ;
  assign n26 = ~n23 & ~n25 ;
  assign n27 = n26 ^ n12 ;
  assign n28 = ~n22 & n27 ;
  assign n29 = n28 ^ n12 ;
  assign n30 = n20 & n29 ;
  assign n31 = n19 & n30 ;
  assign y0 = n31 ;
endmodule
