module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n18 = x0 & x9 ;
  assign n19 = x14 & x16 ;
  assign n20 = x5 & n19 ;
  assign n21 = n18 & n20 ;
  assign n22 = x10 & ~x11 ;
  assign n23 = x12 & x15 ;
  assign n24 = n22 & n23 ;
  assign n25 = ~x7 & ~x8 ;
  assign n26 = x13 & n25 ;
  assign n27 = n24 & n26 ;
  assign n28 = ~x1 & ~x4 ;
  assign n29 = ~x2 & n28 ;
  assign n30 = x3 & x6 ;
  assign n31 = n29 & n30 ;
  assign n32 = n27 & n31 ;
  assign n33 = n21 & n32 ;
  assign y0 = n33 ;
endmodule
