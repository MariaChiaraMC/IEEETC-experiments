module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 ;
  assign n7 = ~x0 & ~x2 ;
  assign n8 = ~x4 & ~x5 ;
  assign n9 = n7 & n8 ;
  assign n10 = ~x3 & n9 ;
  assign n11 = ~x4 & ~n7 ;
  assign n12 = ~n8 & ~n11 ;
  assign n13 = ~x1 & n12 ;
  assign n14 = x5 ^ x0 ;
  assign n15 = x2 & x3 ;
  assign n16 = n15 ^ x5 ;
  assign n17 = ~n14 & n16 ;
  assign n18 = x4 & n17 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = n13 & ~n19 ;
  assign n21 = x4 & x5 ;
  assign n22 = ~x2 & ~n21 ;
  assign n23 = x0 & x5 ;
  assign n24 = x2 & x4 ;
  assign n25 = ~n23 & ~n24 ;
  assign n26 = ~n22 & n25 ;
  assign n27 = n26 ^ x3 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = x4 ^ x2 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = x2 ^ x0 ;
  assign n32 = n31 ^ x5 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = n31 ^ x4 ;
  assign n35 = ~n33 & ~n34 ;
  assign n36 = n35 ^ n31 ;
  assign n37 = ~n30 & n36 ;
  assign n38 = n37 ^ n31 ;
  assign n39 = n38 ^ n26 ;
  assign n40 = ~n28 & n39 ;
  assign n41 = n40 ^ n26 ;
  assign n42 = x1 & n41 ;
  assign n43 = ~n20 & ~n42 ;
  assign n44 = ~n10 & n43 ;
  assign y0 = ~n44 ;
endmodule
