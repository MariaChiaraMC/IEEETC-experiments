module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 ;
  assign n10 = ~x4 & ~x7 ;
  assign n11 = x6 ^ x5 ;
  assign n12 = x1 & ~x2 ;
  assign n13 = ~x8 & n12 ;
  assign n14 = n13 ^ x6 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = x2 & x8 ;
  assign n17 = ~x1 & n16 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = n15 & n18 ;
  assign n20 = n19 ^ n13 ;
  assign n21 = ~n11 & n20 ;
  assign n22 = n10 & n21 ;
  assign n48 = x7 & x8 ;
  assign n49 = x5 & x6 ;
  assign n50 = x1 & x4 ;
  assign n51 = n49 & n50 ;
  assign n52 = ~x1 & ~x4 ;
  assign n53 = x5 & ~x6 ;
  assign n54 = n52 & n53 ;
  assign n55 = ~n51 & ~n54 ;
  assign n56 = n48 & ~n55 ;
  assign n57 = x5 & ~x8 ;
  assign n58 = ~x1 & n57 ;
  assign n59 = x4 & ~x6 ;
  assign n60 = n58 & n59 ;
  assign n61 = x7 & n60 ;
  assign n62 = ~x5 & x8 ;
  assign n63 = x1 & ~x4 ;
  assign n64 = n62 & n63 ;
  assign n65 = x7 ^ x6 ;
  assign n66 = n64 & n65 ;
  assign n67 = ~n61 & ~n66 ;
  assign n68 = ~n56 & n67 ;
  assign n29 = x8 ^ x5 ;
  assign n31 = n29 ^ x4 ;
  assign n32 = n31 ^ n29 ;
  assign n23 = x4 ^ x1 ;
  assign n25 = n23 ^ x6 ;
  assign n24 = n23 ^ x8 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = n27 ^ n23 ;
  assign n30 = n29 ^ n28 ;
  assign n33 = n32 ^ n30 ;
  assign n36 = n28 ^ n23 ;
  assign n34 = n25 ^ n23 ;
  assign n35 = n34 ^ n30 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = ~n33 & n37 ;
  assign n39 = n38 ^ n28 ;
  assign n40 = n39 ^ n34 ;
  assign n41 = n40 ^ n36 ;
  assign n42 = n35 ^ n32 ;
  assign n43 = n39 & n42 ;
  assign n44 = n43 ^ n28 ;
  assign n45 = n44 ^ n30 ;
  assign n46 = n45 ^ n32 ;
  assign n47 = n41 & ~n46 ;
  assign n69 = n68 ^ n47 ;
  assign n70 = n69 ^ n68 ;
  assign n71 = n68 ^ x7 ;
  assign n72 = n71 ^ n68 ;
  assign n73 = n70 & ~n72 ;
  assign n74 = n73 ^ n68 ;
  assign n75 = x2 & ~n74 ;
  assign n76 = n75 ^ n68 ;
  assign n77 = n76 ^ x0 ;
  assign n78 = n77 ^ n76 ;
  assign n79 = n10 & n13 ;
  assign n80 = x6 & x7 ;
  assign n82 = n50 ^ x2 ;
  assign n81 = n52 ^ x8 ;
  assign n83 = n82 ^ n81 ;
  assign n84 = n83 ^ n80 ;
  assign n85 = n81 ^ x2 ;
  assign n86 = n85 ^ n52 ;
  assign n87 = n52 & ~n86 ;
  assign n88 = n87 ^ n81 ;
  assign n89 = n88 ^ n52 ;
  assign n90 = n84 & n89 ;
  assign n91 = n90 ^ n87 ;
  assign n92 = n91 ^ n52 ;
  assign n93 = n80 & n92 ;
  assign n94 = ~n79 & ~n93 ;
  assign n95 = ~x5 & ~n94 ;
  assign n96 = n48 & n50 ;
  assign n97 = ~x2 & n53 ;
  assign n98 = n96 & n97 ;
  assign n99 = ~n58 & ~n62 ;
  assign n100 = x2 & ~x6 ;
  assign n101 = n10 & n100 ;
  assign n102 = ~n99 & n101 ;
  assign n103 = ~n98 & ~n102 ;
  assign n104 = ~n95 & n103 ;
  assign n105 = n104 ^ n76 ;
  assign n106 = n78 & n105 ;
  assign n107 = n106 ^ n76 ;
  assign n108 = ~n22 & n107 ;
  assign n109 = x3 & ~n108 ;
  assign n110 = ~x1 & ~x5 ;
  assign n111 = ~x7 & x8 ;
  assign n112 = ~x0 & n111 ;
  assign n113 = x4 & n100 ;
  assign n114 = n112 & n113 ;
  assign n115 = n110 & n114 ;
  assign n116 = n49 ^ x0 ;
  assign n117 = n49 ^ n12 ;
  assign n118 = n117 ^ n12 ;
  assign n119 = n118 ^ n116 ;
  assign n120 = x2 & ~x5 ;
  assign n121 = n120 ^ x1 ;
  assign n122 = ~x1 & n121 ;
  assign n123 = n122 ^ n12 ;
  assign n124 = n123 ^ x1 ;
  assign n125 = ~n119 & ~n124 ;
  assign n126 = n125 ^ n122 ;
  assign n127 = n126 ^ x1 ;
  assign n128 = n116 & ~n127 ;
  assign n129 = n48 & n128 ;
  assign n130 = ~x0 & ~x5 ;
  assign n131 = n13 & n130 ;
  assign n132 = x6 & n131 ;
  assign n133 = ~n129 & ~n132 ;
  assign n134 = n133 ^ x4 ;
  assign n135 = n134 ^ n133 ;
  assign n136 = n135 ^ x3 ;
  assign n137 = ~x6 & x7 ;
  assign n138 = x8 ^ x7 ;
  assign n139 = x2 & ~n138 ;
  assign n140 = ~n137 & ~n139 ;
  assign n141 = x0 & ~x1 ;
  assign n142 = x5 & ~n100 ;
  assign n143 = n141 & n142 ;
  assign n144 = ~n140 & n143 ;
  assign n145 = x8 & n80 ;
  assign n146 = n120 & n145 ;
  assign n147 = ~x2 & x8 ;
  assign n149 = n110 & n137 ;
  assign n148 = x1 & ~n57 ;
  assign n150 = n149 ^ n148 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = ~x6 & ~x7 ;
  assign n153 = ~n120 & n152 ;
  assign n154 = n153 ^ n149 ;
  assign n155 = n154 ^ n149 ;
  assign n156 = n151 & n155 ;
  assign n157 = n156 ^ n149 ;
  assign n158 = ~n147 & n157 ;
  assign n159 = n158 ^ n149 ;
  assign n160 = ~n146 & ~n159 ;
  assign n161 = ~x0 & ~n160 ;
  assign n162 = n161 ^ n144 ;
  assign n163 = ~n144 & n162 ;
  assign n164 = n163 ^ n133 ;
  assign n165 = n164 ^ n144 ;
  assign n166 = ~n136 & ~n165 ;
  assign n167 = n166 ^ n163 ;
  assign n168 = n167 ^ n144 ;
  assign n169 = ~x3 & ~n168 ;
  assign n170 = n169 ^ x3 ;
  assign n171 = ~n115 & n170 ;
  assign n172 = ~n109 & n171 ;
  assign y0 = ~n172 ;
endmodule
