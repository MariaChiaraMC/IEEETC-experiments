module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 ;
  assign n16 = x2 & ~x3 ;
  assign n17 = n16 ^ x0 ;
  assign n18 = n16 ^ x2 ;
  assign n19 = n16 ^ x4 ;
  assign n20 = ~n16 & ~n19 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = ~n18 & ~n21 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n23 ^ n16 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = n17 & ~n25 ;
  assign n27 = n26 ^ x0 ;
  assign n28 = x6 ^ x5 ;
  assign n29 = n28 ^ x6 ;
  assign n30 = n29 ^ x2 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = x3 ^ x2 ;
  assign n34 = n33 ^ x2 ;
  assign n35 = ~n28 & n34 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = n32 & n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = n38 ^ n33 ;
  assign n40 = n39 ^ n28 ;
  assign n41 = n27 & ~n40 ;
  assign n42 = x1 & ~n41 ;
  assign n43 = ~x11 & ~x13 ;
  assign n44 = ~x10 & n43 ;
  assign n45 = ~x9 & n44 ;
  assign n46 = ~x12 & n45 ;
  assign n47 = ~x2 & x3 ;
  assign n48 = n47 ^ x0 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = x5 & x6 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = ~n49 & n51 ;
  assign n53 = n52 ^ n47 ;
  assign n54 = ~x1 & n53 ;
  assign n55 = n46 & ~n54 ;
  assign n56 = ~n42 & n55 ;
  assign y0 = n56 ;
endmodule
