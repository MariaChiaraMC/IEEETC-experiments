module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 ;
  assign n23 = ~x1 & x3 ;
  assign n22 = x1 ^ x0 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = x2 ^ x1 ;
  assign n27 = n26 ^ x1 ;
  assign n28 = n23 & ~n27 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = n25 & n29 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n31 ^ n26 ;
  assign n33 = n32 ^ n23 ;
  assign n34 = x5 & n33 ;
  assign n35 = ~x4 & n34 ;
  assign n36 = ~x3 & ~x4 ;
  assign n37 = ~x0 & ~x2 ;
  assign n38 = x1 & n37 ;
  assign n39 = n36 & n38 ;
  assign n40 = x14 & ~n39 ;
  assign n236 = ~x19 & ~x20 ;
  assign n41 = ~x12 & ~x13 ;
  assign n42 = x9 & n41 ;
  assign n54 = ~n23 & ~n37 ;
  assign n55 = ~x10 & x11 ;
  assign n56 = ~x6 & ~x7 ;
  assign n57 = n55 & n56 ;
  assign n58 = ~n54 & n57 ;
  assign n43 = x8 ^ x5 ;
  assign n45 = n43 ^ x2 ;
  assign n44 = n43 ^ x8 ;
  assign n46 = n45 ^ n44 ;
  assign n59 = n58 ^ n46 ;
  assign n63 = n59 ^ n45 ;
  assign n64 = n63 ^ n43 ;
  assign n47 = n46 ^ n45 ;
  assign n48 = n47 ^ n43 ;
  assign n49 = n48 ^ n43 ;
  assign n50 = ~x2 & n23 ;
  assign n51 = n50 ^ n45 ;
  assign n52 = n51 ^ n43 ;
  assign n53 = ~n49 & ~n52 ;
  assign n60 = n59 ^ n53 ;
  assign n61 = n60 ^ n43 ;
  assign n62 = ~n48 & ~n61 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = n65 ^ n48 ;
  assign n67 = x10 & ~x11 ;
  assign n68 = n67 ^ n43 ;
  assign n69 = n64 ^ n61 ;
  assign n70 = n69 ^ n48 ;
  assign n71 = ~n68 & ~n70 ;
  assign n72 = n71 ^ n43 ;
  assign n73 = n66 & n72 ;
  assign n74 = n73 ^ n71 ;
  assign n75 = n74 ^ n43 ;
  assign n76 = n75 ^ x8 ;
  assign n77 = n42 & n76 ;
  assign n78 = ~x5 & ~n37 ;
  assign n79 = ~x3 & ~n78 ;
  assign n80 = ~x12 & n56 ;
  assign n81 = ~x13 & ~n80 ;
  assign n82 = ~x9 & ~x10 ;
  assign n84 = ~x0 & ~x1 ;
  assign n85 = ~x9 & ~n84 ;
  assign n86 = ~n37 & ~n50 ;
  assign n87 = ~n85 & ~n86 ;
  assign n88 = ~x5 & ~n87 ;
  assign n83 = x5 & x11 ;
  assign n89 = n88 ^ n83 ;
  assign n90 = n89 ^ n83 ;
  assign n91 = ~x11 & ~x13 ;
  assign n92 = n91 ^ n83 ;
  assign n93 = n92 ^ n83 ;
  assign n94 = ~n90 & n93 ;
  assign n95 = n94 ^ n83 ;
  assign n96 = ~n82 & n95 ;
  assign n97 = n96 ^ n83 ;
  assign n98 = ~n81 & n97 ;
  assign n99 = ~x8 & n98 ;
  assign n100 = ~n79 & ~n99 ;
  assign n101 = ~n77 & n100 ;
  assign n102 = ~x4 & ~n101 ;
  assign n103 = ~x2 & x5 ;
  assign n104 = n103 ^ x2 ;
  assign n105 = n104 ^ n23 ;
  assign n137 = n105 ^ n104 ;
  assign n106 = n41 & ~n84 ;
  assign n107 = n36 & n106 ;
  assign n113 = x11 ^ x10 ;
  assign n114 = n113 ^ n56 ;
  assign n108 = x11 ^ x8 ;
  assign n109 = n108 ^ n56 ;
  assign n110 = n109 ^ x11 ;
  assign n111 = n110 ^ x9 ;
  assign n112 = n111 ^ n56 ;
  assign n115 = n114 ^ n112 ;
  assign n118 = n111 ^ x9 ;
  assign n116 = x11 ^ x9 ;
  assign n117 = n116 ^ n112 ;
  assign n119 = n118 ^ n117 ;
  assign n120 = ~n115 & ~n119 ;
  assign n121 = n120 ^ n111 ;
  assign n122 = n121 ^ n116 ;
  assign n123 = n122 ^ n118 ;
  assign n124 = n117 ^ n114 ;
  assign n125 = ~n121 & n124 ;
  assign n126 = n125 ^ n111 ;
  assign n127 = n126 ^ n112 ;
  assign n128 = n127 ^ n114 ;
  assign n129 = ~n123 & n128 ;
  assign n130 = n107 & n129 ;
  assign n131 = n130 ^ n105 ;
  assign n132 = n131 ^ n104 ;
  assign n133 = n105 ^ n103 ;
  assign n134 = n133 ^ n130 ;
  assign n135 = n134 ^ n132 ;
  assign n136 = ~n132 & ~n135 ;
  assign n138 = n137 ^ n136 ;
  assign n139 = n138 ^ n132 ;
  assign n140 = ~x8 & ~x10 ;
  assign n141 = ~x8 & ~x11 ;
  assign n142 = ~x10 & ~x13 ;
  assign n143 = ~n141 & ~n142 ;
  assign n144 = ~n140 & ~n143 ;
  assign n145 = x11 & ~x12 ;
  assign n146 = ~x13 & ~n145 ;
  assign n147 = x15 & ~n142 ;
  assign n148 = ~x6 & ~x17 ;
  assign n149 = ~x1 & n148 ;
  assign n150 = ~n147 & n149 ;
  assign n151 = ~n146 & n150 ;
  assign n152 = x13 ^ x10 ;
  assign n153 = n152 ^ x13 ;
  assign n154 = n153 ^ x11 ;
  assign n155 = ~x7 & x16 ;
  assign n156 = n155 ^ x8 ;
  assign n157 = ~x8 & n156 ;
  assign n158 = n157 ^ x13 ;
  assign n159 = n158 ^ x8 ;
  assign n160 = ~n154 & n159 ;
  assign n161 = n160 ^ n157 ;
  assign n162 = n161 ^ x8 ;
  assign n163 = x11 & ~n162 ;
  assign n164 = n163 ^ x11 ;
  assign n165 = ~x9 & ~n164 ;
  assign n166 = n151 & ~n165 ;
  assign n167 = ~n144 & n166 ;
  assign n168 = x5 & ~n167 ;
  assign n169 = n168 ^ n104 ;
  assign n170 = n136 ^ n132 ;
  assign n171 = ~n169 & ~n170 ;
  assign n172 = n171 ^ n104 ;
  assign n173 = ~n139 & n172 ;
  assign n174 = n173 ^ n104 ;
  assign n175 = n174 ^ x2 ;
  assign n176 = n175 ^ n104 ;
  assign n213 = x4 & ~n84 ;
  assign n177 = ~x8 & ~x9 ;
  assign n178 = n55 & n177 ;
  assign n179 = x2 & n178 ;
  assign n180 = ~x4 & ~n179 ;
  assign n181 = x0 & ~n180 ;
  assign n182 = n42 & n83 ;
  assign n183 = n140 & n182 ;
  assign n184 = ~n181 & ~n183 ;
  assign n185 = ~x1 & ~n184 ;
  assign n186 = ~x12 & x13 ;
  assign n187 = n145 ^ x10 ;
  assign n188 = n187 ^ n145 ;
  assign n189 = x13 & n141 ;
  assign n190 = n189 ^ n145 ;
  assign n191 = ~n188 & n190 ;
  assign n192 = n191 ^ n145 ;
  assign n193 = x9 & n192 ;
  assign n194 = ~n186 & ~n193 ;
  assign n195 = ~x2 & ~n194 ;
  assign n196 = x13 ^ x1 ;
  assign n197 = x13 ^ x0 ;
  assign n198 = n197 ^ x0 ;
  assign n199 = n198 ^ n196 ;
  assign n200 = ~x10 & ~x11 ;
  assign n201 = n200 ^ x12 ;
  assign n202 = ~x12 & ~n201 ;
  assign n203 = n202 ^ x0 ;
  assign n204 = n203 ^ x12 ;
  assign n205 = n199 & ~n204 ;
  assign n206 = n205 ^ n202 ;
  assign n207 = n206 ^ x12 ;
  assign n208 = n196 & ~n207 ;
  assign n209 = n208 ^ x1 ;
  assign n210 = ~n195 & ~n209 ;
  assign n211 = x5 & ~n210 ;
  assign n212 = ~n185 & ~n211 ;
  assign n214 = n213 ^ n212 ;
  assign n215 = n214 ^ x3 ;
  assign n223 = n215 ^ n214 ;
  assign n216 = ~x0 & x2 ;
  assign n217 = n216 ^ n215 ;
  assign n218 = n217 ^ n214 ;
  assign n219 = n215 ^ n212 ;
  assign n220 = n219 ^ n216 ;
  assign n221 = n220 ^ n218 ;
  assign n222 = n218 & ~n221 ;
  assign n224 = n223 ^ n222 ;
  assign n225 = n224 ^ n218 ;
  assign n226 = n214 ^ x5 ;
  assign n227 = n222 ^ n218 ;
  assign n228 = ~n226 & n227 ;
  assign n229 = n228 ^ n214 ;
  assign n230 = ~n225 & ~n229 ;
  assign n231 = n230 ^ n214 ;
  assign n232 = n231 ^ n213 ;
  assign n233 = n232 ^ n214 ;
  assign n234 = ~n176 & ~n233 ;
  assign n235 = ~n102 & n234 ;
  assign n237 = n236 ^ n235 ;
  assign n238 = n237 ^ n235 ;
  assign n239 = n235 ^ x18 ;
  assign n240 = ~n238 & n239 ;
  assign n241 = n240 ^ n235 ;
  assign n242 = n40 & n241 ;
  assign n243 = ~n35 & n242 ;
  assign y0 = ~n243 ;
endmodule
