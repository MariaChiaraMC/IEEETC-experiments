module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 ;
  assign n13 = ~x7 & ~x11 ;
  assign n14 = ~x8 & ~x10 ;
  assign n15 = ~x9 & n14 ;
  assign n16 = n13 & n15 ;
  assign n17 = x2 & ~x3 ;
  assign n18 = n17 ^ x0 ;
  assign n19 = n17 ^ x2 ;
  assign n20 = n17 ^ x4 ;
  assign n21 = ~n17 & ~n20 ;
  assign n22 = n21 ^ n17 ;
  assign n23 = ~n19 & ~n22 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n24 ^ n17 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = n18 & ~n26 ;
  assign n28 = n27 ^ x0 ;
  assign n29 = x5 ^ x2 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = n30 ^ x6 ;
  assign n32 = x5 ^ x3 ;
  assign n33 = n32 ^ x5 ;
  assign n34 = x6 ^ x5 ;
  assign n35 = ~n33 & n34 ;
  assign n36 = n35 ^ x5 ;
  assign n37 = n31 & n36 ;
  assign n38 = n37 ^ n29 ;
  assign n39 = n28 & ~n38 ;
  assign n40 = n39 ^ x1 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = ~x0 & x5 ;
  assign n43 = x6 & n42 ;
  assign n44 = x0 & x3 ;
  assign n45 = ~x2 & n44 ;
  assign n46 = ~n43 & ~n45 ;
  assign n47 = n46 ^ n39 ;
  assign n48 = ~n41 & n47 ;
  assign n49 = n48 ^ n39 ;
  assign n50 = n16 & n49 ;
  assign y0 = n50 ;
endmodule
