module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 ;
  assign n11 = x4 & ~x8 ;
  assign n12 = x6 & x7 ;
  assign n13 = x1 & x9 ;
  assign n14 = ~x3 & ~x5 ;
  assign n15 = n13 & n14 ;
  assign n16 = n12 & n15 ;
  assign n17 = x3 & ~x9 ;
  assign n18 = ~x1 & x5 ;
  assign n19 = ~x6 & ~x7 ;
  assign n20 = n18 & n19 ;
  assign n21 = n17 & n20 ;
  assign n22 = ~n16 & ~n21 ;
  assign n23 = x0 & ~n22 ;
  assign n24 = x1 & x3 ;
  assign n25 = x7 & ~x9 ;
  assign n26 = ~x0 & ~x6 ;
  assign n27 = n25 & n26 ;
  assign n28 = n24 & n27 ;
  assign n29 = ~x5 & n28 ;
  assign n30 = ~n23 & ~n29 ;
  assign n31 = n11 & ~n30 ;
  assign n114 = x6 & ~x7 ;
  assign n199 = n11 & n114 ;
  assign n259 = n18 & n199 ;
  assign n44 = x7 & x8 ;
  assign n122 = ~x6 & n44 ;
  assign n260 = n19 ^ x1 ;
  assign n261 = n260 ^ n19 ;
  assign n62 = x5 & ~x8 ;
  assign n262 = n62 & n114 ;
  assign n263 = n262 ^ n19 ;
  assign n264 = n261 & n263 ;
  assign n265 = n264 ^ n19 ;
  assign n266 = ~x4 & n265 ;
  assign n267 = ~n122 & ~n266 ;
  assign n268 = ~x4 & x5 ;
  assign n269 = x1 & n268 ;
  assign n270 = n269 ^ x5 ;
  assign n271 = ~n267 & ~n270 ;
  assign n272 = ~n259 & ~n271 ;
  assign n273 = x0 & ~n272 ;
  assign n42 = ~x0 & ~x1 ;
  assign n33 = x7 & ~x8 ;
  assign n274 = ~x4 & ~n33 ;
  assign n277 = x6 ^ x4 ;
  assign n275 = x6 ^ x5 ;
  assign n283 = n277 ^ n275 ;
  assign n276 = n275 ^ n12 ;
  assign n278 = n277 ^ n276 ;
  assign n279 = n275 ^ x6 ;
  assign n280 = n279 ^ n12 ;
  assign n281 = n280 ^ n278 ;
  assign n282 = ~n278 & ~n281 ;
  assign n284 = n283 ^ n282 ;
  assign n285 = n284 ^ n278 ;
  assign n286 = n277 ^ n44 ;
  assign n287 = n282 ^ n278 ;
  assign n288 = ~n286 & ~n287 ;
  assign n289 = n288 ^ n277 ;
  assign n290 = ~n285 & ~n289 ;
  assign n291 = n290 ^ n277 ;
  assign n292 = n291 ^ n277 ;
  assign n293 = ~n274 & n292 ;
  assign n294 = n42 & n293 ;
  assign n202 = ~x8 & n114 ;
  assign n203 = ~x4 & n202 ;
  assign n295 = ~x0 & ~x5 ;
  assign n296 = n203 & n295 ;
  assign n297 = x1 & n296 ;
  assign n298 = x3 & ~n297 ;
  assign n299 = ~n294 & n298 ;
  assign n300 = ~n273 & n299 ;
  assign n301 = x0 & x7 ;
  assign n102 = ~x1 & x8 ;
  assign n302 = n102 ^ x8 ;
  assign n303 = ~x4 & ~n302 ;
  assign n304 = n303 ^ x8 ;
  assign n305 = n301 & ~n304 ;
  assign n306 = n305 ^ x6 ;
  assign n314 = n306 ^ n305 ;
  assign n217 = ~x7 & x8 ;
  assign n307 = ~x4 & n217 ;
  assign n308 = n307 ^ n306 ;
  assign n309 = n308 ^ n305 ;
  assign n310 = n307 ^ n42 ;
  assign n311 = n310 ^ n307 ;
  assign n312 = n311 ^ n309 ;
  assign n313 = ~n309 & ~n312 ;
  assign n315 = n314 ^ n313 ;
  assign n316 = n315 ^ n309 ;
  assign n317 = ~n217 & ~n274 ;
  assign n318 = n317 ^ n305 ;
  assign n319 = n313 ^ n309 ;
  assign n320 = n318 & ~n319 ;
  assign n321 = n320 ^ n305 ;
  assign n322 = ~n316 & ~n321 ;
  assign n323 = n322 ^ n305 ;
  assign n324 = n323 ^ x6 ;
  assign n325 = n324 ^ n305 ;
  assign n326 = ~x5 & n325 ;
  assign n146 = ~x6 & n42 ;
  assign n327 = n33 & n146 ;
  assign n328 = x4 & n327 ;
  assign n329 = ~x3 & ~n328 ;
  assign n330 = ~n326 & n329 ;
  assign n331 = ~n300 & ~n330 ;
  assign n32 = x0 & x3 ;
  assign n34 = ~x5 & ~x6 ;
  assign n35 = n33 & n34 ;
  assign n36 = ~n32 & n35 ;
  assign n37 = ~x0 & ~x3 ;
  assign n38 = n13 ^ x1 ;
  assign n39 = ~n37 & ~n38 ;
  assign n40 = n39 ^ x1 ;
  assign n41 = n36 & ~n40 ;
  assign n43 = x3 & n42 ;
  assign n45 = x9 & n44 ;
  assign n46 = n43 & n45 ;
  assign n47 = ~x5 & n46 ;
  assign n48 = ~x0 & x5 ;
  assign n49 = ~x8 & ~x9 ;
  assign n50 = n48 & ~n49 ;
  assign n51 = ~x1 & ~x3 ;
  assign n52 = n51 ^ n24 ;
  assign n53 = ~x8 & n52 ;
  assign n54 = n53 ^ n24 ;
  assign n55 = n50 & n54 ;
  assign n56 = n55 ^ x7 ;
  assign n57 = n56 ^ n55 ;
  assign n58 = n57 ^ n47 ;
  assign n59 = ~x5 & x8 ;
  assign n60 = ~x1 & n59 ;
  assign n61 = ~n42 & n60 ;
  assign n63 = ~n42 & n62 ;
  assign n66 = n63 ^ n48 ;
  assign n67 = n66 ^ n63 ;
  assign n64 = n63 ^ x8 ;
  assign n65 = n64 ^ n63 ;
  assign n68 = n67 ^ n65 ;
  assign n69 = n63 ^ x1 ;
  assign n70 = n69 ^ n63 ;
  assign n71 = n70 ^ n67 ;
  assign n72 = n67 & ~n71 ;
  assign n73 = n72 ^ n67 ;
  assign n74 = n68 & n73 ;
  assign n75 = n74 ^ n72 ;
  assign n76 = n75 ^ n63 ;
  assign n77 = n76 ^ n67 ;
  assign n78 = ~x3 & n77 ;
  assign n79 = n78 ^ n63 ;
  assign n80 = ~n61 & ~n79 ;
  assign n81 = n80 ^ x9 ;
  assign n82 = ~n80 & n81 ;
  assign n83 = n82 ^ n55 ;
  assign n84 = n83 ^ n80 ;
  assign n85 = ~n58 & ~n84 ;
  assign n86 = n85 ^ n82 ;
  assign n87 = n86 ^ n80 ;
  assign n88 = ~n47 & ~n87 ;
  assign n89 = n88 ^ n47 ;
  assign n90 = x6 & n89 ;
  assign n91 = ~n41 & ~n90 ;
  assign n92 = ~x0 & n59 ;
  assign n93 = x0 & ~x3 ;
  assign n94 = x5 & n93 ;
  assign n95 = ~n92 & ~n94 ;
  assign n96 = n13 & ~n95 ;
  assign n97 = x5 & x9 ;
  assign n98 = x8 & n97 ;
  assign n99 = n43 & n98 ;
  assign n100 = n62 ^ n42 ;
  assign n101 = n100 ^ n42 ;
  assign n103 = x0 & ~n102 ;
  assign n104 = ~n59 & n103 ;
  assign n105 = n104 ^ n42 ;
  assign n106 = ~n101 & n105 ;
  assign n107 = n106 ^ n42 ;
  assign n108 = n17 & n107 ;
  assign n109 = ~n99 & ~n108 ;
  assign n110 = ~n96 & n109 ;
  assign n111 = n19 & ~n110 ;
  assign n112 = ~x4 & ~n111 ;
  assign n113 = n91 & n112 ;
  assign n115 = n97 & n102 ;
  assign n116 = ~n114 & n115 ;
  assign n118 = ~x5 & ~x9 ;
  assign n117 = x1 & n114 ;
  assign n119 = n118 ^ n117 ;
  assign n120 = n117 ^ n98 ;
  assign n121 = n120 ^ n98 ;
  assign n123 = n122 ^ n98 ;
  assign n124 = ~n121 & ~n123 ;
  assign n125 = n124 ^ n98 ;
  assign n126 = n119 & n125 ;
  assign n127 = n126 ^ n118 ;
  assign n128 = ~n116 & ~n127 ;
  assign n129 = n32 & ~n128 ;
  assign n130 = n129 ^ x4 ;
  assign n131 = x9 ^ x1 ;
  assign n132 = n92 ^ x9 ;
  assign n133 = n132 ^ n92 ;
  assign n134 = n133 ^ n131 ;
  assign n135 = x8 ^ x5 ;
  assign n136 = ~x8 & ~n135 ;
  assign n137 = n136 ^ n92 ;
  assign n138 = n137 ^ x8 ;
  assign n139 = n134 & ~n138 ;
  assign n140 = n139 ^ n136 ;
  assign n141 = n140 ^ x8 ;
  assign n142 = n131 & ~n141 ;
  assign n143 = n12 & n142 ;
  assign n144 = n143 ^ x3 ;
  assign n145 = n144 ^ n143 ;
  assign n147 = n45 & n146 ;
  assign n148 = x5 & n147 ;
  assign n152 = x6 ^ x1 ;
  assign n153 = n152 ^ x7 ;
  assign n149 = x6 ^ x0 ;
  assign n150 = n149 ^ x7 ;
  assign n160 = n153 ^ n150 ;
  assign n151 = n150 ^ x7 ;
  assign n154 = n153 ^ n151 ;
  assign n155 = n154 ^ n150 ;
  assign n156 = n151 ^ x6 ;
  assign n157 = n156 ^ n151 ;
  assign n158 = n157 ^ n155 ;
  assign n159 = n155 & ~n158 ;
  assign n161 = n160 ^ n159 ;
  assign n162 = n161 ^ n155 ;
  assign n163 = n150 ^ n25 ;
  assign n164 = n159 ^ n155 ;
  assign n165 = ~n163 & n164 ;
  assign n166 = n165 ^ n150 ;
  assign n167 = ~n162 & ~n166 ;
  assign n168 = n167 ^ n150 ;
  assign n169 = n168 ^ n150 ;
  assign n170 = n62 & n169 ;
  assign n171 = ~n148 & ~n170 ;
  assign n172 = n171 ^ n143 ;
  assign n173 = ~n145 & ~n172 ;
  assign n174 = n173 ^ n143 ;
  assign n175 = n174 ^ n129 ;
  assign n176 = ~n130 & n175 ;
  assign n177 = n176 ^ n173 ;
  assign n178 = n177 ^ n143 ;
  assign n179 = n178 ^ x4 ;
  assign n180 = ~n129 & ~n179 ;
  assign n181 = n180 ^ n129 ;
  assign n182 = ~n113 & n181 ;
  assign n183 = ~x1 & ~x6 ;
  assign n184 = n32 & n183 ;
  assign n185 = ~x7 & ~x8 ;
  assign n186 = n185 ^ n44 ;
  assign n187 = n186 ^ n184 ;
  assign n188 = n44 ^ x9 ;
  assign n189 = n44 ^ x5 ;
  assign n190 = n189 ^ n188 ;
  assign n191 = ~n188 & n190 ;
  assign n192 = n191 ^ n44 ;
  assign n193 = n192 ^ n188 ;
  assign n194 = n187 & ~n193 ;
  assign n195 = n194 ^ n191 ;
  assign n196 = n195 ^ n188 ;
  assign n197 = n184 & ~n196 ;
  assign n198 = ~n182 & ~n197 ;
  assign n332 = n331 ^ n198 ;
  assign n200 = n32 & n199 ;
  assign n201 = ~x5 & ~n200 ;
  assign n218 = n26 & n217 ;
  assign n219 = n44 ^ x6 ;
  assign n220 = n219 ^ n44 ;
  assign n221 = n186 & ~n220 ;
  assign n222 = n221 ^ n44 ;
  assign n223 = x0 & n222 ;
  assign n224 = ~n218 & ~n223 ;
  assign n225 = ~x4 & ~n224 ;
  assign n226 = ~x3 & n225 ;
  assign n204 = x4 & n44 ;
  assign n205 = ~n122 & ~n204 ;
  assign n206 = ~n203 & n205 ;
  assign n207 = n93 & ~n206 ;
  assign n208 = ~x0 & x3 ;
  assign n209 = n33 ^ x4 ;
  assign n210 = n209 ^ n33 ;
  assign n211 = n185 ^ n33 ;
  assign n212 = n210 & n211 ;
  assign n213 = n212 ^ n33 ;
  assign n214 = n208 & n213 ;
  assign n215 = ~x6 & n214 ;
  assign n216 = ~n207 & ~n215 ;
  assign n227 = n226 ^ n216 ;
  assign n228 = n227 ^ n216 ;
  assign n229 = x6 & n204 ;
  assign n230 = n37 & n229 ;
  assign n231 = n230 ^ n216 ;
  assign n232 = n231 ^ n216 ;
  assign n233 = ~n228 & ~n232 ;
  assign n234 = n233 ^ n216 ;
  assign n235 = x1 & n234 ;
  assign n236 = n235 ^ n216 ;
  assign n237 = n201 & n236 ;
  assign n238 = x7 & n26 ;
  assign n239 = n54 & n238 ;
  assign n240 = n239 ^ x4 ;
  assign n241 = n240 ^ n239 ;
  assign n242 = ~n37 & ~n51 ;
  assign n243 = n202 & ~n242 ;
  assign n244 = x0 & n24 ;
  assign n245 = n44 ^ x8 ;
  assign n246 = ~x6 & ~n245 ;
  assign n247 = n246 ^ x8 ;
  assign n248 = n244 & ~n247 ;
  assign n249 = ~n243 & ~n248 ;
  assign n250 = n249 ^ n239 ;
  assign n251 = n241 & ~n250 ;
  assign n252 = n251 ^ n239 ;
  assign n253 = x5 & ~n252 ;
  assign n254 = ~n237 & ~n253 ;
  assign n255 = n93 & n204 ;
  assign n256 = n183 & n255 ;
  assign n257 = ~n254 & ~n256 ;
  assign n258 = n257 ^ n198 ;
  assign n333 = n332 ^ n258 ;
  assign n334 = n332 ^ x9 ;
  assign n335 = n334 ^ n332 ;
  assign n336 = ~n333 & ~n335 ;
  assign n337 = n336 ^ n332 ;
  assign n338 = x2 & ~n337 ;
  assign n339 = n338 ^ n198 ;
  assign n340 = ~n31 & n339 ;
  assign y0 = ~n340 ;
endmodule
