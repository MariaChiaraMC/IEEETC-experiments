module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 ;
  assign n8 = ~x1 & x6 ;
  assign n9 = ~x4 & x5 ;
  assign n10 = x3 & n9 ;
  assign n11 = x2 & ~x4 ;
  assign n12 = n11 ^ x0 ;
  assign n13 = n12 ^ n10 ;
  assign n16 = ~x3 & ~x5 ;
  assign n14 = ~x2 & ~x3 ;
  assign n15 = ~x5 & ~n14 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = ~n11 & n17 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = n13 & ~n19 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n21 ^ n16 ;
  assign n23 = n22 ^ n11 ;
  assign n24 = ~n10 & n23 ;
  assign n25 = n8 & ~n24 ;
  assign n26 = x2 & ~x6 ;
  assign n27 = x5 & n26 ;
  assign n28 = x3 & n27 ;
  assign n29 = x0 & n28 ;
  assign n30 = ~n25 & ~n29 ;
  assign n31 = x3 & x6 ;
  assign n32 = x4 & n31 ;
  assign n33 = n9 & n14 ;
  assign n34 = ~n32 & ~n33 ;
  assign n35 = x0 & ~n34 ;
  assign n36 = x3 ^ x2 ;
  assign n37 = x3 ^ x0 ;
  assign n38 = ~x5 & x6 ;
  assign n39 = n38 ^ x0 ;
  assign n40 = x0 & n39 ;
  assign n41 = n40 ^ x0 ;
  assign n42 = ~n37 & n41 ;
  assign n43 = n42 ^ n40 ;
  assign n44 = n43 ^ x0 ;
  assign n45 = n44 ^ n38 ;
  assign n46 = n36 & n45 ;
  assign n47 = ~n27 & ~n46 ;
  assign n48 = ~n35 & n47 ;
  assign n49 = x1 & ~n48 ;
  assign n50 = x5 ^ x4 ;
  assign n51 = ~x1 & ~x2 ;
  assign n52 = n51 ^ x3 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n53 ^ n50 ;
  assign n55 = ~x0 & ~x2 ;
  assign n56 = n55 ^ x5 ;
  assign n57 = n55 & ~n56 ;
  assign n58 = n57 ^ n51 ;
  assign n59 = n58 ^ n55 ;
  assign n60 = n54 & ~n59 ;
  assign n61 = n60 ^ n57 ;
  assign n62 = n61 ^ n55 ;
  assign n63 = n50 & n62 ;
  assign n64 = ~x6 & n63 ;
  assign n65 = x0 & n8 ;
  assign n66 = n65 ^ n51 ;
  assign n67 = n66 ^ x3 ;
  assign n74 = n67 ^ n66 ;
  assign n68 = n67 ^ x5 ;
  assign n69 = n68 ^ n66 ;
  assign n70 = n67 ^ n65 ;
  assign n71 = n70 ^ x5 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = n69 & ~n72 ;
  assign n75 = n74 ^ n73 ;
  assign n76 = n75 ^ n69 ;
  assign n77 = n66 ^ x6 ;
  assign n78 = n73 ^ n69 ;
  assign n79 = n77 & n78 ;
  assign n80 = n79 ^ n66 ;
  assign n81 = ~n76 & n80 ;
  assign n82 = n81 ^ n66 ;
  assign n83 = n82 ^ n51 ;
  assign n84 = n83 ^ n66 ;
  assign n85 = x4 & n84 ;
  assign n86 = ~n64 & ~n85 ;
  assign n87 = ~n49 & n86 ;
  assign n88 = n30 & n87 ;
  assign y0 = ~n88 ;
endmodule
