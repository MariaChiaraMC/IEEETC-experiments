module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n10 = ~x4 & x5 ;
  assign n11 = ~x6 & ~n10 ;
  assign n12 = x3 & ~x4 ;
  assign n13 = x2 & n12 ;
  assign n14 = x1 & n13 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n11 & ~n15 ;
  assign n17 = x5 ^ x1 ;
  assign n18 = n17 ^ x6 ;
  assign n19 = x3 ^ x2 ;
  assign n20 = x6 ^ x5 ;
  assign n21 = x4 ^ x3 ;
  assign n22 = n21 ^ x3 ;
  assign n23 = ~n20 & ~n22 ;
  assign n24 = n23 ^ x3 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = ~n19 & n25 ;
  assign n27 = n26 ^ x5 ;
  assign n28 = n18 & ~n27 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = x6 & n29 ;
  assign n31 = n30 ^ x6 ;
  assign n32 = ~n16 & ~n31 ;
  assign y0 = n32 ;
endmodule
