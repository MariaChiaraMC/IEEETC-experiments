module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 ;
  assign n28 = x2 & ~x3 ;
  assign n79 = ~x1 & x4 ;
  assign n159 = ~x5 & n79 ;
  assign n160 = ~x6 & ~x7 ;
  assign n161 = n159 & n160 ;
  assign n162 = n28 & n161 ;
  assign n163 = x0 & ~n162 ;
  assign n11 = ~x5 & x8 ;
  assign n12 = ~x2 & ~n11 ;
  assign n13 = x7 & x8 ;
  assign n14 = x5 & ~n13 ;
  assign n15 = n12 & ~n14 ;
  assign n16 = ~x3 & ~x4 ;
  assign n17 = ~x5 & ~x8 ;
  assign n18 = n16 & n17 ;
  assign n19 = ~n15 & ~n18 ;
  assign n20 = x0 & x6 ;
  assign n21 = ~x1 & n20 ;
  assign n22 = ~n19 & n21 ;
  assign n23 = x7 & n17 ;
  assign n24 = ~x3 & n23 ;
  assign n25 = ~n15 & ~n24 ;
  assign n26 = ~x6 & ~n25 ;
  assign n27 = x4 & x8 ;
  assign n29 = x6 & x7 ;
  assign n30 = x5 & n29 ;
  assign n31 = n28 & n30 ;
  assign n32 = n27 & n31 ;
  assign n33 = ~n26 & ~n32 ;
  assign n34 = n33 ^ x1 ;
  assign n35 = n34 ^ n33 ;
  assign n36 = n35 ^ x0 ;
  assign n37 = ~x4 & ~x6 ;
  assign n38 = x5 & n28 ;
  assign n39 = n13 & n38 ;
  assign n40 = n37 & n39 ;
  assign n41 = x5 & ~x8 ;
  assign n42 = ~n11 & ~n41 ;
  assign n43 = ~n27 & ~n42 ;
  assign n44 = x6 ^ x3 ;
  assign n45 = x7 & ~n44 ;
  assign n46 = n43 & n45 ;
  assign n47 = ~x4 & x6 ;
  assign n48 = x3 & n47 ;
  assign n49 = n41 & n48 ;
  assign n50 = ~x2 & ~n49 ;
  assign n51 = ~n46 & n50 ;
  assign n52 = x3 & x7 ;
  assign n53 = x8 ^ x5 ;
  assign n54 = x8 ^ x6 ;
  assign n55 = n54 ^ x6 ;
  assign n56 = n37 ^ x6 ;
  assign n57 = ~n55 & n56 ;
  assign n58 = n57 ^ x6 ;
  assign n59 = ~n53 & n58 ;
  assign n60 = n52 & n59 ;
  assign n61 = x4 & ~n44 ;
  assign n62 = n17 & n61 ;
  assign n63 = x2 & ~n62 ;
  assign n64 = ~n60 & n63 ;
  assign n65 = ~n51 & ~n64 ;
  assign n66 = n65 ^ n40 ;
  assign n67 = ~n40 & n66 ;
  assign n68 = n67 ^ n33 ;
  assign n69 = n68 ^ n40 ;
  assign n70 = ~n36 & ~n69 ;
  assign n71 = n70 ^ n67 ;
  assign n72 = n71 ^ n40 ;
  assign n73 = ~x0 & ~n72 ;
  assign n74 = n73 ^ x0 ;
  assign n75 = ~n22 & n74 ;
  assign n93 = ~x6 & ~n16 ;
  assign n94 = ~n42 & n93 ;
  assign n76 = n17 & n37 ;
  assign n77 = x1 & ~x4 ;
  assign n78 = x6 & ~n77 ;
  assign n80 = n79 ^ x8 ;
  assign n81 = n79 ^ x5 ;
  assign n82 = n80 & n81 ;
  assign n83 = n78 & n82 ;
  assign n84 = ~n76 & ~n83 ;
  assign n85 = n84 ^ n17 ;
  assign n86 = n85 ^ n84 ;
  assign n87 = n84 ^ n47 ;
  assign n88 = n87 ^ n84 ;
  assign n89 = n86 & n88 ;
  assign n90 = n89 ^ n84 ;
  assign n91 = x3 & ~n90 ;
  assign n92 = n91 ^ n84 ;
  assign n95 = n94 ^ n92 ;
  assign n96 = x3 & n79 ;
  assign n97 = n96 ^ n92 ;
  assign n98 = n92 ^ x0 ;
  assign n99 = n92 & ~n98 ;
  assign n100 = n99 ^ n92 ;
  assign n101 = n97 & n100 ;
  assign n102 = n101 ^ n99 ;
  assign n103 = n102 ^ n92 ;
  assign n104 = n103 ^ x0 ;
  assign n105 = ~n95 & ~n104 ;
  assign n106 = n105 ^ n94 ;
  assign n107 = n106 ^ x1 ;
  assign n108 = n107 ^ x2 ;
  assign n124 = n108 ^ n107 ;
  assign n109 = x6 ^ x0 ;
  assign n110 = n109 ^ x6 ;
  assign n111 = ~x3 & x6 ;
  assign n112 = ~x2 & x4 ;
  assign n113 = n111 & n112 ;
  assign n114 = n113 ^ x6 ;
  assign n115 = ~n110 & ~n114 ;
  assign n116 = n115 ^ x6 ;
  assign n117 = ~n42 & ~n116 ;
  assign n118 = n117 ^ n108 ;
  assign n119 = n118 ^ n107 ;
  assign n120 = n108 ^ n106 ;
  assign n121 = n120 ^ n117 ;
  assign n122 = n121 ^ n119 ;
  assign n123 = ~n119 & ~n122 ;
  assign n125 = n124 ^ n123 ;
  assign n126 = n125 ^ n119 ;
  assign n127 = x3 & n27 ;
  assign n128 = ~x0 & n127 ;
  assign n129 = x5 & n128 ;
  assign n130 = n16 & n41 ;
  assign n131 = ~n129 & ~n130 ;
  assign n132 = ~x6 & ~n131 ;
  assign n133 = n132 ^ n107 ;
  assign n134 = n123 ^ n119 ;
  assign n135 = ~n133 & ~n134 ;
  assign n136 = n135 ^ n107 ;
  assign n137 = ~n126 & n136 ;
  assign n138 = n137 ^ n107 ;
  assign n139 = n138 ^ x1 ;
  assign n140 = n139 ^ n107 ;
  assign n141 = n140 ^ x7 ;
  assign n142 = n141 ^ n140 ;
  assign n143 = n142 ^ n75 ;
  assign n144 = x2 & x3 ;
  assign n145 = x6 & n144 ;
  assign n146 = ~x1 & n145 ;
  assign n147 = ~n20 & ~n146 ;
  assign n148 = n147 ^ n17 ;
  assign n149 = ~n147 & ~n148 ;
  assign n150 = n149 ^ n140 ;
  assign n151 = n150 ^ n147 ;
  assign n152 = n143 & ~n151 ;
  assign n153 = n152 ^ n149 ;
  assign n154 = n153 ^ n147 ;
  assign n155 = n75 & ~n154 ;
  assign n156 = n155 ^ n75 ;
  assign n164 = n163 ^ n156 ;
  assign n165 = n164 ^ n156 ;
  assign n157 = n156 ^ x8 ;
  assign n158 = n157 ^ n156 ;
  assign n166 = n165 ^ n158 ;
  assign n167 = n30 & n77 ;
  assign n168 = ~n161 & ~n167 ;
  assign n169 = ~x0 & ~n144 ;
  assign n170 = ~n168 & ~n169 ;
  assign n171 = x6 ^ x4 ;
  assign n172 = x7 ^ x6 ;
  assign n173 = ~n171 & n172 ;
  assign n174 = ~x3 & ~n173 ;
  assign n175 = x1 & ~x2 ;
  assign n177 = ~x4 & n29 ;
  assign n178 = x3 & ~n177 ;
  assign n176 = x4 & n160 ;
  assign n179 = n178 ^ n176 ;
  assign n180 = x5 & ~n179 ;
  assign n181 = n180 ^ n178 ;
  assign n182 = n175 & ~n181 ;
  assign n183 = ~n174 & n182 ;
  assign n184 = ~n170 & ~n183 ;
  assign n185 = x7 ^ x4 ;
  assign n186 = n185 ^ x1 ;
  assign n187 = n186 ^ n38 ;
  assign n188 = x6 ^ x1 ;
  assign n189 = n188 ^ x6 ;
  assign n190 = n172 ^ x6 ;
  assign n191 = n189 & n190 ;
  assign n192 = n191 ^ x6 ;
  assign n193 = n192 ^ n186 ;
  assign n194 = ~n187 & ~n193 ;
  assign n195 = n194 ^ n191 ;
  assign n196 = n195 ^ x6 ;
  assign n197 = n196 ^ n38 ;
  assign n198 = ~n186 & n197 ;
  assign n199 = n198 ^ n186 ;
  assign n200 = n184 & n199 ;
  assign n201 = n200 ^ n156 ;
  assign n202 = n201 ^ n156 ;
  assign n203 = n202 ^ n165 ;
  assign n204 = ~n165 & n203 ;
  assign n205 = n204 ^ n165 ;
  assign n206 = n166 & ~n205 ;
  assign n207 = n206 ^ n204 ;
  assign n208 = n207 ^ n156 ;
  assign n209 = n208 ^ n165 ;
  assign n210 = x9 & n209 ;
  assign n211 = n210 ^ n156 ;
  assign y0 = ~n211 ;
endmodule
