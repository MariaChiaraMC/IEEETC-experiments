module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 ;
  assign n16 = x12 ^ x11 ;
  assign n17 = ~x3 & x4 ;
  assign n18 = x13 & ~n17 ;
  assign n19 = ~x2 & n18 ;
  assign n20 = ~x10 & ~x13 ;
  assign n21 = ~x1 & x5 ;
  assign n22 = n21 ^ x2 ;
  assign n23 = n21 ^ x3 ;
  assign n24 = n23 ^ x3 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = x3 ^ x1 ;
  assign n27 = ~x3 & x6 ;
  assign n28 = ~n26 & n27 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = x6 ^ x4 ;
  assign n31 = x5 & ~n30 ;
  assign n32 = n31 ^ x4 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = ~n29 & ~n33 ;
  assign n35 = n34 ^ x3 ;
  assign n36 = n35 ^ n29 ;
  assign n37 = ~n25 & n36 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = n38 ^ n29 ;
  assign n40 = n22 & ~n39 ;
  assign n41 = n40 ^ x0 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = x5 & ~x6 ;
  assign n44 = n43 ^ x2 ;
  assign n45 = ~x1 & ~n44 ;
  assign n46 = n45 ^ x2 ;
  assign n47 = n46 ^ n40 ;
  assign n48 = ~n42 & ~n47 ;
  assign n49 = n48 ^ n40 ;
  assign n50 = n20 & n49 ;
  assign n51 = ~n19 & ~n50 ;
  assign n52 = ~x9 & ~n51 ;
  assign n53 = x10 & ~x13 ;
  assign n54 = x14 ^ x13 ;
  assign n55 = ~x2 & ~x3 ;
  assign n56 = x0 & ~x1 ;
  assign n57 = ~n55 & n56 ;
  assign n58 = n57 ^ n53 ;
  assign n59 = ~n54 & n58 ;
  assign n60 = n59 ^ n57 ;
  assign n61 = n53 & n60 ;
  assign n62 = n61 ^ x10 ;
  assign n63 = ~n52 & ~n62 ;
  assign n64 = n63 ^ x12 ;
  assign n65 = n64 ^ n63 ;
  assign n66 = n65 ^ n16 ;
  assign n67 = n53 ^ x9 ;
  assign n68 = n53 & n67 ;
  assign n69 = n68 ^ n63 ;
  assign n70 = n69 ^ n53 ;
  assign n71 = ~n66 & ~n70 ;
  assign n72 = n71 ^ n68 ;
  assign n73 = n72 ^ n53 ;
  assign n74 = ~n16 & n73 ;
  assign y0 = n74 ;
endmodule
