module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 ;
  assign n25 = x1 & x2 ;
  assign n26 = x14 ^ x3 ;
  assign n27 = n25 & ~n26 ;
  assign n28 = x5 & ~n27 ;
  assign n29 = x15 & x16 ;
  assign n30 = x17 ^ x5 ;
  assign n31 = n30 ^ x17 ;
  assign n32 = ~x3 & ~x14 ;
  assign n33 = n32 ^ x17 ;
  assign n34 = n31 & n33 ;
  assign n35 = n34 ^ x17 ;
  assign n36 = x18 & ~n35 ;
  assign n37 = n29 & ~n36 ;
  assign n38 = ~n28 & n37 ;
  assign n39 = x14 & x16 ;
  assign n40 = x3 & ~x15 ;
  assign n41 = n39 & ~n40 ;
  assign n42 = x5 & x17 ;
  assign n43 = ~n41 & n42 ;
  assign n44 = n25 & n43 ;
  assign n45 = ~n38 & ~n44 ;
  assign n46 = ~x1 & ~x2 ;
  assign n47 = x3 & x14 ;
  assign n48 = ~x9 & n47 ;
  assign n49 = x0 & n32 ;
  assign n50 = ~n48 & ~n49 ;
  assign n51 = n46 & ~n50 ;
  assign n52 = ~x0 & x5 ;
  assign n53 = ~x0 & x10 ;
  assign n54 = n53 ^ n46 ;
  assign n55 = x14 ^ x1 ;
  assign n56 = n55 ^ x1 ;
  assign n57 = ~x2 & x11 ;
  assign n58 = n57 ^ x1 ;
  assign n59 = n56 & ~n58 ;
  assign n60 = n59 ^ x1 ;
  assign n61 = n60 ^ n53 ;
  assign n62 = ~n54 & ~n61 ;
  assign n63 = n62 ^ n59 ;
  assign n64 = n63 ^ x1 ;
  assign n65 = n64 ^ n46 ;
  assign n66 = n53 & n65 ;
  assign n67 = n66 ^ n53 ;
  assign n68 = ~n52 & ~n67 ;
  assign n69 = ~n51 & n68 ;
  assign n70 = x4 & ~n69 ;
  assign n71 = ~n45 & n70 ;
  assign n72 = x6 ^ x3 ;
  assign n73 = n72 ^ x6 ;
  assign n74 = x7 ^ x6 ;
  assign n75 = n73 & n74 ;
  assign n76 = n75 ^ x6 ;
  assign n77 = x17 & n76 ;
  assign n78 = n25 & n77 ;
  assign n79 = ~x18 & x23 ;
  assign n80 = n29 & n79 ;
  assign n81 = n27 & n80 ;
  assign n82 = ~n78 & ~n81 ;
  assign n83 = n52 & ~n82 ;
  assign n84 = ~n71 & ~n83 ;
  assign y0 = ~n84 ;
endmodule
