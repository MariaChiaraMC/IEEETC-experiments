module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 ;
  assign n17 = x4 & x5 ;
  assign n18 = ~x1 & n17 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = n19 ^ x0 ;
  assign n100 = n20 ^ n19 ;
  assign n21 = x14 & ~x15 ;
  assign n22 = x12 & ~x13 ;
  assign n23 = ~n21 & ~n22 ;
  assign n24 = ~x0 & ~x5 ;
  assign n25 = x4 & ~x6 ;
  assign n26 = n24 & n25 ;
  assign n27 = ~x0 & ~x4 ;
  assign n28 = n27 ^ n17 ;
  assign n29 = n28 ^ x7 ;
  assign n41 = n29 ^ n28 ;
  assign n30 = ~x5 & x6 ;
  assign n31 = ~x8 & ~x9 ;
  assign n32 = x11 ^ x10 ;
  assign n33 = n31 & n32 ;
  assign n34 = n30 & n33 ;
  assign n35 = n34 ^ n29 ;
  assign n36 = n35 ^ n28 ;
  assign n37 = n29 ^ n17 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = ~n36 & ~n39 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = n42 ^ n36 ;
  assign n44 = x5 & ~x6 ;
  assign n45 = ~n30 & ~n44 ;
  assign n46 = n45 ^ n28 ;
  assign n47 = n40 ^ n36 ;
  assign n48 = n46 & ~n47 ;
  assign n49 = n48 ^ n28 ;
  assign n50 = ~n43 & n49 ;
  assign n51 = n50 ^ n28 ;
  assign n52 = n51 ^ n27 ;
  assign n53 = n52 ^ n28 ;
  assign n54 = ~n26 & ~n53 ;
  assign n55 = ~n23 & ~n54 ;
  assign n56 = x6 & n17 ;
  assign n57 = x10 & ~x11 ;
  assign n58 = n22 & n57 ;
  assign n59 = n21 & n58 ;
  assign n60 = n56 & n59 ;
  assign n61 = x12 & x14 ;
  assign n62 = n56 & n61 ;
  assign n63 = ~x10 & x11 ;
  assign n64 = x15 ^ x13 ;
  assign n65 = n63 & n64 ;
  assign n66 = n62 & n65 ;
  assign n67 = ~x4 & x7 ;
  assign n68 = ~x13 & n21 ;
  assign n69 = ~x12 & n68 ;
  assign n70 = ~n67 & ~n69 ;
  assign n71 = n44 & ~n70 ;
  assign n72 = x14 & x15 ;
  assign n73 = x4 & x7 ;
  assign n74 = n22 & n73 ;
  assign n75 = n72 & n74 ;
  assign n76 = ~n71 & ~n75 ;
  assign n77 = ~x0 & ~n76 ;
  assign n78 = x6 & ~n23 ;
  assign n79 = n17 ^ x10 ;
  assign n80 = n79 ^ n17 ;
  assign n81 = ~x4 & n24 ;
  assign n82 = n81 ^ n17 ;
  assign n83 = ~n80 & n82 ;
  assign n84 = n83 ^ n17 ;
  assign n85 = n78 & n84 ;
  assign n86 = ~n77 & ~n85 ;
  assign n87 = ~x11 & ~n86 ;
  assign n88 = ~n66 & ~n87 ;
  assign n89 = x9 ^ x8 ;
  assign n90 = ~n88 & n89 ;
  assign n91 = ~n60 & ~n90 ;
  assign n92 = ~n55 & n91 ;
  assign n93 = ~x1 & ~n92 ;
  assign n94 = n93 ^ n20 ;
  assign n95 = n94 ^ n19 ;
  assign n96 = n20 ^ n18 ;
  assign n97 = n96 ^ n93 ;
  assign n98 = n97 ^ n95 ;
  assign n99 = ~n95 & n98 ;
  assign n101 = n100 ^ n99 ;
  assign n102 = n101 ^ n95 ;
  assign n103 = ~x9 & ~x10 ;
  assign n104 = ~x11 & ~x12 ;
  assign n105 = x14 ^ x13 ;
  assign n106 = n105 ^ x15 ;
  assign n107 = n106 ^ x13 ;
  assign n108 = n107 ^ n104 ;
  assign n109 = x15 ^ x8 ;
  assign n110 = ~x13 & n109 ;
  assign n111 = n110 ^ x15 ;
  assign n112 = ~n108 & ~n111 ;
  assign n113 = n112 ^ n110 ;
  assign n114 = n113 ^ x15 ;
  assign n115 = n114 ^ x13 ;
  assign n116 = n104 & n115 ;
  assign n117 = ~n103 & ~n116 ;
  assign n118 = ~x14 & ~x15 ;
  assign n119 = x10 ^ x9 ;
  assign n120 = n118 & n119 ;
  assign n121 = ~x13 & n120 ;
  assign n122 = x8 & ~n121 ;
  assign n123 = ~n117 & ~n122 ;
  assign n124 = ~x7 & ~n123 ;
  assign n125 = x1 & n30 ;
  assign n126 = x4 & n125 ;
  assign n127 = ~n124 & n126 ;
  assign n128 = n127 ^ n19 ;
  assign n129 = n99 ^ n95 ;
  assign n130 = n128 & ~n129 ;
  assign n131 = n130 ^ n19 ;
  assign n132 = ~n102 & ~n131 ;
  assign n133 = n132 ^ n19 ;
  assign n134 = n133 ^ x2 ;
  assign n135 = n134 ^ n19 ;
  assign n136 = ~x3 & ~n135 ;
  assign y0 = n136 ;
endmodule
