module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 ;
  assign n9 = x3 & x5 ;
  assign n10 = ~x3 & ~x5 ;
  assign n11 = ~x2 & x6 ;
  assign n12 = ~n10 & n11 ;
  assign n13 = ~n9 & n12 ;
  assign n14 = n13 ^ x2 ;
  assign n15 = ~x1 & n14 ;
  assign n16 = n15 ^ x2 ;
  assign n17 = ~x0 & n16 ;
  assign n33 = x0 & x1 ;
  assign n18 = ~x2 & x3 ;
  assign n19 = n18 ^ x0 ;
  assign n20 = x3 ^ x1 ;
  assign n21 = n20 ^ x1 ;
  assign n22 = ~x6 & ~x7 ;
  assign n23 = n22 ^ x1 ;
  assign n24 = n21 & n23 ;
  assign n25 = n24 ^ x1 ;
  assign n26 = n25 ^ n18 ;
  assign n27 = n19 & ~n26 ;
  assign n28 = n27 ^ n24 ;
  assign n29 = n28 ^ x1 ;
  assign n30 = n29 ^ x0 ;
  assign n31 = ~n18 & ~n30 ;
  assign n32 = n31 ^ n18 ;
  assign n34 = n33 ^ n32 ;
  assign n35 = ~n9 & ~n34 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = ~x0 & ~x5 ;
  assign n38 = ~x3 & ~n37 ;
  assign n39 = n38 ^ x5 ;
  assign n40 = n39 ^ x6 ;
  assign n47 = n40 ^ n39 ;
  assign n41 = n40 ^ n33 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = n38 ^ n33 ;
  assign n44 = n43 ^ n33 ;
  assign n45 = n44 ^ n42 ;
  assign n46 = n42 & ~n45 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = n48 ^ n42 ;
  assign n50 = n39 ^ x7 ;
  assign n51 = n46 ^ n42 ;
  assign n52 = ~n50 & n51 ;
  assign n53 = n52 ^ n39 ;
  assign n54 = n49 & ~n53 ;
  assign n55 = n54 ^ n39 ;
  assign n56 = n55 ^ n38 ;
  assign n57 = n56 ^ n39 ;
  assign n58 = ~x2 & n57 ;
  assign n59 = x2 & x5 ;
  assign n60 = n59 ^ x3 ;
  assign n61 = x7 ^ x5 ;
  assign n62 = n61 ^ x7 ;
  assign n63 = x6 & x7 ;
  assign n64 = n63 ^ x7 ;
  assign n65 = ~n62 & ~n64 ;
  assign n66 = n65 ^ x7 ;
  assign n67 = n66 ^ n59 ;
  assign n68 = n60 & n67 ;
  assign n69 = n68 ^ n65 ;
  assign n70 = n69 ^ x7 ;
  assign n71 = n70 ^ x3 ;
  assign n72 = ~n59 & n71 ;
  assign n73 = n72 ^ n59 ;
  assign n74 = n73 ^ n59 ;
  assign n75 = n74 ^ x1 ;
  assign n76 = n75 ^ n74 ;
  assign n77 = x3 ^ x2 ;
  assign n78 = x3 ^ x0 ;
  assign n79 = n78 ^ x0 ;
  assign n80 = n37 ^ x0 ;
  assign n81 = n79 & n80 ;
  assign n82 = n81 ^ x0 ;
  assign n83 = n77 & n82 ;
  assign n84 = n83 ^ n74 ;
  assign n85 = ~n76 & ~n84 ;
  assign n86 = n85 ^ n74 ;
  assign n87 = ~n58 & n86 ;
  assign n88 = ~n36 & n87 ;
  assign n89 = n88 ^ x4 ;
  assign n90 = n89 ^ n88 ;
  assign n91 = ~x1 & ~x3 ;
  assign n92 = n22 & n91 ;
  assign n93 = n37 & n92 ;
  assign n95 = n59 ^ x5 ;
  assign n96 = n95 ^ n59 ;
  assign n94 = n60 ^ n59 ;
  assign n97 = n96 ^ n94 ;
  assign n98 = n59 ^ x0 ;
  assign n99 = n98 ^ n59 ;
  assign n100 = n99 ^ n96 ;
  assign n101 = ~n96 & ~n100 ;
  assign n102 = n101 ^ n96 ;
  assign n103 = ~n97 & ~n102 ;
  assign n104 = n103 ^ n101 ;
  assign n105 = n104 ^ n59 ;
  assign n106 = n105 ^ n96 ;
  assign n107 = x1 & ~n106 ;
  assign n108 = n107 ^ n59 ;
  assign n109 = ~n63 & n108 ;
  assign n110 = ~x0 & n63 ;
  assign n111 = ~n10 & ~n110 ;
  assign n112 = x2 & ~n111 ;
  assign n113 = n9 & ~n33 ;
  assign n114 = x6 ^ x0 ;
  assign n115 = x6 ^ x1 ;
  assign n116 = n115 ^ x1 ;
  assign n117 = x7 ^ x1 ;
  assign n118 = n116 & n117 ;
  assign n119 = n118 ^ x1 ;
  assign n120 = ~n114 & n119 ;
  assign n121 = n120 ^ x0 ;
  assign n122 = n113 & ~n121 ;
  assign n123 = ~n112 & ~n122 ;
  assign n124 = ~n109 & n123 ;
  assign n125 = ~n93 & n124 ;
  assign n126 = n125 ^ n88 ;
  assign n127 = n90 & n126 ;
  assign n128 = n127 ^ n88 ;
  assign n129 = ~n17 & n128 ;
  assign y0 = ~n129 ;
endmodule
