module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 ;
  assign n9 = x4 & x6 ;
  assign n10 = x5 & x7 ;
  assign n11 = ~x5 & ~x7 ;
  assign n12 = ~n10 & ~n11 ;
  assign n13 = n9 & ~n12 ;
  assign n14 = x1 & ~x2 ;
  assign n15 = ~x2 & ~x7 ;
  assign n16 = ~x4 & n15 ;
  assign n17 = ~n14 & ~n16 ;
  assign n18 = x6 & ~x7 ;
  assign n19 = x5 & n18 ;
  assign n20 = x1 & n19 ;
  assign n21 = x7 ^ x4 ;
  assign n22 = x5 ^ x4 ;
  assign n23 = n22 ^ x4 ;
  assign n24 = n21 & ~n23 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = x2 & n25 ;
  assign n27 = ~n20 & ~n26 ;
  assign n28 = n17 & n27 ;
  assign n29 = ~n13 & n28 ;
  assign n30 = ~x3 & ~n29 ;
  assign n31 = ~x2 & x3 ;
  assign n32 = n31 ^ x1 ;
  assign n33 = ~x2 & x4 ;
  assign n34 = ~x5 & ~n33 ;
  assign n35 = ~n9 & n34 ;
  assign n36 = n35 ^ n31 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = x4 & n18 ;
  assign n39 = ~n10 & ~n38 ;
  assign n40 = n39 ^ n35 ;
  assign n41 = n37 & n40 ;
  assign n42 = n41 ^ n35 ;
  assign n43 = ~n32 & ~n42 ;
  assign n44 = n43 ^ x1 ;
  assign n45 = x5 & ~x7 ;
  assign n46 = ~x3 & ~x6 ;
  assign n47 = n45 & n46 ;
  assign n48 = n47 ^ x4 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = n49 ^ n44 ;
  assign n51 = ~x1 & ~x6 ;
  assign n52 = n10 & n51 ;
  assign n53 = x3 & ~n52 ;
  assign n54 = ~x2 & n45 ;
  assign n55 = n54 ^ n53 ;
  assign n56 = n53 & ~n55 ;
  assign n57 = n56 ^ n47 ;
  assign n58 = n57 ^ n53 ;
  assign n59 = ~n50 & n58 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = n60 ^ n53 ;
  assign n62 = n44 & n61 ;
  assign n63 = n62 ^ n44 ;
  assign n64 = ~n30 & n63 ;
  assign n65 = ~x0 & ~n64 ;
  assign n66 = x6 & n10 ;
  assign n67 = x0 & n66 ;
  assign n68 = n67 ^ x2 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = n69 ^ x1 ;
  assign n71 = n18 ^ x3 ;
  assign n72 = ~n18 & ~n71 ;
  assign n73 = n72 ^ n67 ;
  assign n74 = n73 ^ n18 ;
  assign n75 = n70 & n74 ;
  assign n76 = n75 ^ n72 ;
  assign n77 = n76 ^ n18 ;
  assign n78 = ~x1 & ~n77 ;
  assign n79 = n78 ^ x1 ;
  assign n82 = x4 ^ x3 ;
  assign n86 = n82 ^ x4 ;
  assign n80 = x5 ^ x2 ;
  assign n81 = n80 ^ x5 ;
  assign n83 = n82 ^ x5 ;
  assign n84 = n83 ^ x4 ;
  assign n85 = ~n81 & ~n84 ;
  assign n87 = n86 ^ n85 ;
  assign n88 = x6 ^ x4 ;
  assign n89 = x7 & n88 ;
  assign n90 = n89 ^ x4 ;
  assign n91 = n86 & n90 ;
  assign n92 = n91 ^ n89 ;
  assign n93 = n87 & n92 ;
  assign n94 = n93 ^ x4 ;
  assign n95 = n94 ^ x4 ;
  assign n96 = ~n79 & n95 ;
  assign n97 = ~x3 & n14 ;
  assign n98 = n11 ^ x4 ;
  assign n99 = n98 ^ n11 ;
  assign n100 = x6 & ~n10 ;
  assign n101 = n100 ^ n11 ;
  assign n102 = ~n99 & ~n101 ;
  assign n103 = n102 ^ n11 ;
  assign n104 = n97 & n103 ;
  assign n105 = ~n96 & ~n104 ;
  assign n106 = ~n65 & n105 ;
  assign y0 = ~n106 ;
endmodule
