module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 ;
  assign n49 = ~x0 & ~x4 ;
  assign n50 = x3 & n49 ;
  assign n51 = ~x5 & n50 ;
  assign n15 = x1 ^ x0 ;
  assign n16 = n15 ^ x1 ;
  assign n17 = ~x7 & ~x8 ;
  assign n18 = x11 & x13 ;
  assign n19 = ~x10 & ~n18 ;
  assign n20 = ~n17 & n19 ;
  assign n21 = ~x6 & ~x9 ;
  assign n22 = x7 & x8 ;
  assign n23 = x4 & ~n22 ;
  assign n24 = x5 & ~n23 ;
  assign n25 = n21 & ~n24 ;
  assign n26 = ~x11 & ~x13 ;
  assign n27 = n26 ^ x12 ;
  assign n28 = n25 & ~n27 ;
  assign n29 = n20 & n28 ;
  assign n37 = n29 ^ x3 ;
  assign n38 = n37 ^ x3 ;
  assign n39 = n37 & ~n38 ;
  assign n31 = x5 ^ x3 ;
  assign n30 = n29 ^ x1 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = n31 ^ n29 ;
  assign n34 = n33 ^ x3 ;
  assign n35 = n32 & ~n34 ;
  assign n42 = n39 ^ n35 ;
  assign n36 = n35 ^ n16 ;
  assign n40 = n39 ^ n37 ;
  assign n41 = n36 & n40 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = n16 & n43 ;
  assign n45 = n44 ^ n35 ;
  assign n46 = n45 ^ n39 ;
  assign n47 = n46 ^ n41 ;
  assign n48 = n47 ^ n15 ;
  assign n52 = n51 ^ n48 ;
  assign n53 = ~x2 & n52 ;
  assign n54 = n53 ^ n51 ;
  assign y0 = n54 ;
endmodule
