module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 ;
  output y0 ;
  wire n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 ;
  assign n23 = x1 ^ x0 ;
  assign n24 = x2 ^ x1 ;
  assign n25 = n24 ^ x5 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = x5 ^ x3 ;
  assign n28 = x5 ^ x1 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = ~n27 & ~n29 ;
  assign n31 = n30 ^ x5 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = n26 & ~n32 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ n27 ;
  assign n36 = n23 & ~n35 ;
  assign n37 = ~x4 & n36 ;
  assign n38 = ~x19 & ~x20 ;
  assign n39 = n38 ^ x18 ;
  assign n40 = n39 ^ x18 ;
  assign n41 = ~x1 & ~x8 ;
  assign n42 = ~x9 & ~x10 ;
  assign n43 = x11 & n42 ;
  assign n44 = x0 & x2 ;
  assign n45 = n43 & n44 ;
  assign n46 = n41 & n45 ;
  assign n47 = x5 ^ x4 ;
  assign n48 = ~x12 & ~x13 ;
  assign n49 = ~x0 & ~x1 ;
  assign n50 = n48 & ~n49 ;
  assign n57 = x11 ^ x10 ;
  assign n52 = ~x6 & ~x7 ;
  assign n58 = n57 ^ n52 ;
  assign n51 = x11 ^ x8 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n53 ^ x11 ;
  assign n55 = n54 ^ x9 ;
  assign n56 = n55 ^ n52 ;
  assign n59 = n58 ^ n56 ;
  assign n62 = n55 ^ x9 ;
  assign n60 = x11 ^ x9 ;
  assign n61 = n60 ^ n56 ;
  assign n63 = n62 ^ n61 ;
  assign n64 = ~n59 & ~n63 ;
  assign n65 = n64 ^ n55 ;
  assign n66 = n65 ^ n60 ;
  assign n67 = n66 ^ n62 ;
  assign n68 = n61 ^ n58 ;
  assign n69 = ~n65 & n68 ;
  assign n70 = n69 ^ n55 ;
  assign n71 = n70 ^ n56 ;
  assign n72 = n71 ^ n58 ;
  assign n73 = ~n67 & n72 ;
  assign n74 = n50 & n73 ;
  assign n75 = n74 ^ x0 ;
  assign n76 = x2 & ~n75 ;
  assign n77 = n76 ^ x0 ;
  assign n78 = n77 ^ x5 ;
  assign n79 = n78 ^ n77 ;
  assign n80 = x12 & ~x13 ;
  assign n81 = ~x6 & ~n80 ;
  assign n82 = ~x7 & ~n81 ;
  assign n83 = ~x17 & ~n82 ;
  assign n84 = x8 ^ x7 ;
  assign n85 = n84 ^ x7 ;
  assign n86 = x10 & ~x13 ;
  assign n87 = n86 ^ x7 ;
  assign n88 = n85 & ~n87 ;
  assign n89 = n88 ^ x7 ;
  assign n90 = x11 & ~n89 ;
  assign n91 = n90 ^ x13 ;
  assign n92 = n91 ^ n83 ;
  assign n93 = ~x15 & n42 ;
  assign n94 = n93 ^ x12 ;
  assign n95 = ~x13 & ~n94 ;
  assign n96 = n95 ^ n93 ;
  assign n97 = ~n92 & n96 ;
  assign n98 = n97 ^ n95 ;
  assign n99 = n98 ^ n93 ;
  assign n100 = n99 ^ x13 ;
  assign n101 = n83 & ~n100 ;
  assign n102 = ~x1 & ~n101 ;
  assign n103 = ~x8 & x10 ;
  assign n104 = ~x16 & ~n103 ;
  assign n105 = ~x7 & n104 ;
  assign n106 = ~n102 & ~n105 ;
  assign n107 = x2 & ~n106 ;
  assign n108 = x0 & ~x1 ;
  assign n109 = ~x0 & x1 ;
  assign n110 = ~x2 & x13 ;
  assign n111 = n110 ^ x12 ;
  assign n112 = x1 & x2 ;
  assign n113 = x9 & ~n112 ;
  assign n114 = ~x10 & ~n41 ;
  assign n115 = x11 & ~n114 ;
  assign n116 = n113 & n115 ;
  assign n117 = n116 ^ n110 ;
  assign n118 = n117 ^ n116 ;
  assign n119 = n118 ^ n111 ;
  assign n120 = ~x8 & ~x10 ;
  assign n121 = x9 & n120 ;
  assign n122 = ~x11 & n121 ;
  assign n123 = n122 ^ x0 ;
  assign n124 = ~x0 & n123 ;
  assign n125 = n124 ^ n116 ;
  assign n126 = n125 ^ x0 ;
  assign n127 = ~n119 & ~n126 ;
  assign n128 = n127 ^ n124 ;
  assign n129 = n128 ^ x0 ;
  assign n130 = ~n111 & ~n129 ;
  assign n131 = n130 ^ n110 ;
  assign n132 = ~n109 & ~n131 ;
  assign n133 = ~n108 & n132 ;
  assign n134 = ~n107 & n133 ;
  assign n135 = n134 ^ n77 ;
  assign n136 = n79 & ~n135 ;
  assign n137 = n136 ^ n77 ;
  assign n138 = ~n47 & n137 ;
  assign n139 = n138 ^ x4 ;
  assign n140 = ~n46 & n139 ;
  assign n141 = ~x3 & ~n140 ;
  assign n142 = ~x1 & x3 ;
  assign n143 = ~x2 & n142 ;
  assign n144 = x5 & n143 ;
  assign n145 = x4 & ~x5 ;
  assign n147 = x2 & ~x21 ;
  assign n146 = x1 & x3 ;
  assign n148 = n147 ^ n146 ;
  assign n149 = n146 ^ n108 ;
  assign n150 = n146 & ~n149 ;
  assign n151 = n150 ^ n146 ;
  assign n152 = ~n148 & n151 ;
  assign n153 = n152 ^ n150 ;
  assign n154 = n153 ^ n146 ;
  assign n155 = n154 ^ n108 ;
  assign n156 = n145 & ~n155 ;
  assign n157 = n156 ^ n145 ;
  assign n158 = ~n144 & ~n157 ;
  assign n159 = ~n141 & n158 ;
  assign n181 = x9 & n48 ;
  assign n160 = ~x13 & ~n52 ;
  assign n161 = ~n80 & ~n160 ;
  assign n162 = ~x11 & ~n42 ;
  assign n163 = ~x13 & n162 ;
  assign n164 = n163 ^ x5 ;
  assign n165 = n163 ^ n43 ;
  assign n166 = n165 ^ n43 ;
  assign n167 = n166 ^ n164 ;
  assign n168 = ~x0 & ~x2 ;
  assign n169 = ~n143 & ~n168 ;
  assign n170 = ~x9 & ~n49 ;
  assign n171 = n170 ^ n169 ;
  assign n172 = ~n169 & n171 ;
  assign n173 = n172 ^ n43 ;
  assign n174 = n173 ^ n169 ;
  assign n175 = n167 & n174 ;
  assign n176 = n175 ^ n172 ;
  assign n177 = n176 ^ n169 ;
  assign n178 = n164 & ~n177 ;
  assign n179 = n178 ^ x5 ;
  assign n180 = n161 & n179 ;
  assign n182 = n181 ^ n180 ;
  assign n183 = n182 ^ x8 ;
  assign n191 = n183 ^ n182 ;
  assign n184 = ~x2 & x5 ;
  assign n185 = n184 ^ n183 ;
  assign n186 = n185 ^ n182 ;
  assign n187 = n183 ^ n180 ;
  assign n188 = n187 ^ n184 ;
  assign n189 = n188 ^ n186 ;
  assign n190 = n186 & ~n189 ;
  assign n192 = n191 ^ n190 ;
  assign n193 = n192 ^ n186 ;
  assign n194 = x11 & n52 ;
  assign n195 = ~x10 & n194 ;
  assign n196 = ~n142 & ~n168 ;
  assign n197 = n195 & ~n196 ;
  assign n198 = x10 & ~x11 ;
  assign n199 = ~x5 & ~n143 ;
  assign n200 = n198 & ~n199 ;
  assign n201 = ~n197 & ~n200 ;
  assign n202 = n201 ^ n182 ;
  assign n203 = n190 ^ n186 ;
  assign n204 = n202 & n203 ;
  assign n205 = n204 ^ n182 ;
  assign n206 = ~n193 & n205 ;
  assign n207 = n206 ^ n182 ;
  assign n208 = n207 ^ n181 ;
  assign n209 = n208 ^ n182 ;
  assign n210 = n209 ^ n112 ;
  assign n211 = n210 ^ x4 ;
  assign n220 = n211 ^ n210 ;
  assign n212 = ~x3 & x16 ;
  assign n213 = x5 & ~n212 ;
  assign n214 = n213 ^ n211 ;
  assign n215 = n214 ^ n210 ;
  assign n216 = n213 ^ n112 ;
  assign n217 = n216 ^ n213 ;
  assign n218 = n217 ^ n215 ;
  assign n219 = n215 & n218 ;
  assign n221 = n220 ^ n219 ;
  assign n222 = n221 ^ n215 ;
  assign n223 = n210 ^ x0 ;
  assign n224 = n219 ^ n215 ;
  assign n225 = n223 & n224 ;
  assign n226 = n225 ^ n210 ;
  assign n227 = ~n222 & n226 ;
  assign n228 = n227 ^ n210 ;
  assign n229 = n228 ^ n112 ;
  assign n230 = n229 ^ n210 ;
  assign n231 = n159 & ~n230 ;
  assign n232 = n231 ^ x18 ;
  assign n233 = n40 & n232 ;
  assign n234 = n233 ^ x18 ;
  assign n235 = x14 & n234 ;
  assign n236 = ~n37 & n235 ;
  assign y0 = ~n236 ;
endmodule
