module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 ;
  assign n19 = x12 & ~x13 ;
  assign n20 = x14 & ~x15 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = x10 ^ x5 ;
  assign n23 = x10 ^ x6 ;
  assign n24 = n23 ^ x6 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = ~x8 & ~x9 ;
  assign n27 = x8 & x9 ;
  assign n28 = ~n26 & ~n27 ;
  assign n29 = n28 ^ x0 ;
  assign n30 = ~x0 & ~n29 ;
  assign n31 = n30 ^ x6 ;
  assign n32 = n31 ^ x0 ;
  assign n33 = n25 & ~n32 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ x0 ;
  assign n36 = ~n22 & ~n35 ;
  assign n37 = ~x11 & n36 ;
  assign n17 = ~x0 & ~x5 ;
  assign n38 = x6 & x7 ;
  assign n39 = n17 & ~n38 ;
  assign n40 = x5 & x7 ;
  assign n41 = ~n39 & ~n40 ;
  assign n42 = ~n37 & n41 ;
  assign n43 = ~n21 & ~n42 ;
  assign n44 = x6 & x12 ;
  assign n45 = ~x10 & x11 ;
  assign n46 = n44 & n45 ;
  assign n47 = x15 ^ x13 ;
  assign n48 = n46 & n47 ;
  assign n49 = x14 & n48 ;
  assign n50 = ~x0 & ~n49 ;
  assign n51 = x5 & ~n50 ;
  assign n52 = ~n43 & ~n51 ;
  assign n18 = x6 & n17 ;
  assign n53 = n52 ^ n18 ;
  assign n54 = n53 ^ x1 ;
  assign n92 = n54 ^ n53 ;
  assign n55 = ~x11 & ~x12 ;
  assign n56 = ~x13 & ~x15 ;
  assign n57 = n56 ^ x8 ;
  assign n58 = n57 ^ x14 ;
  assign n65 = n58 ^ n56 ;
  assign n59 = n58 ^ x1 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = x14 ^ x1 ;
  assign n62 = n61 ^ x1 ;
  assign n63 = n62 ^ n60 ;
  assign n64 = n60 & ~n63 ;
  assign n66 = n65 ^ n64 ;
  assign n67 = n66 ^ n60 ;
  assign n68 = n56 ^ n47 ;
  assign n69 = n64 ^ n60 ;
  assign n70 = n68 & n69 ;
  assign n71 = n70 ^ n56 ;
  assign n72 = n67 & n71 ;
  assign n73 = n72 ^ n56 ;
  assign n74 = n73 ^ n56 ;
  assign n75 = n55 & n74 ;
  assign n76 = x7 & x14 ;
  assign n77 = n76 ^ x9 ;
  assign n78 = n77 ^ x9 ;
  assign n79 = n27 ^ x9 ;
  assign n80 = n79 ^ x9 ;
  assign n81 = ~n78 & ~n80 ;
  assign n82 = n81 ^ x9 ;
  assign n83 = x10 & n82 ;
  assign n84 = n83 ^ x9 ;
  assign n85 = n75 & n84 ;
  assign n86 = n85 ^ n54 ;
  assign n87 = n86 ^ n53 ;
  assign n88 = n85 ^ n18 ;
  assign n89 = n88 ^ n85 ;
  assign n90 = n89 ^ n87 ;
  assign n91 = n87 & n90 ;
  assign n93 = n92 ^ n91 ;
  assign n94 = n93 ^ n87 ;
  assign n95 = n53 ^ x7 ;
  assign n96 = n91 ^ n87 ;
  assign n97 = n95 & n96 ;
  assign n98 = n97 ^ n53 ;
  assign n99 = ~n94 & ~n98 ;
  assign n100 = n99 ^ n53 ;
  assign n101 = n100 ^ n18 ;
  assign n102 = n101 ^ n53 ;
  assign n103 = x4 & n102 ;
  assign n104 = ~x4 & ~x7 ;
  assign n105 = ~x6 & x7 ;
  assign n106 = n26 & n105 ;
  assign n107 = n45 & n106 ;
  assign n108 = ~n104 & ~n107 ;
  assign n109 = x5 & ~n108 ;
  assign n110 = ~n21 & n109 ;
  assign n114 = ~x6 & ~n28 ;
  assign n115 = n40 & ~n114 ;
  assign n111 = ~x4 & ~x5 ;
  assign n112 = x7 ^ x6 ;
  assign n113 = n111 & n112 ;
  assign n116 = n115 ^ n113 ;
  assign n117 = n116 ^ x10 ;
  assign n124 = n117 ^ n116 ;
  assign n118 = n117 ^ n21 ;
  assign n119 = n118 ^ n116 ;
  assign n120 = n113 ^ n21 ;
  assign n121 = n120 ^ n21 ;
  assign n122 = n121 ^ n119 ;
  assign n123 = n119 & ~n122 ;
  assign n125 = n124 ^ n123 ;
  assign n126 = n125 ^ n119 ;
  assign n127 = n116 ^ n106 ;
  assign n128 = n123 ^ n119 ;
  assign n129 = n127 & n128 ;
  assign n130 = n129 ^ n116 ;
  assign n131 = ~n126 & n130 ;
  assign n132 = n131 ^ n116 ;
  assign n133 = n132 ^ n113 ;
  assign n134 = n133 ^ n116 ;
  assign n135 = ~x11 & n134 ;
  assign n136 = ~n110 & ~n135 ;
  assign n137 = ~x1 & ~n136 ;
  assign n138 = ~x0 & n137 ;
  assign n139 = ~n103 & ~n138 ;
  assign y0 = ~n139 ;
endmodule
