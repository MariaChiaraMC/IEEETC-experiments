module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 ;
  assign n16 = ~x8 & x9 ;
  assign n17 = ~x4 & ~x10 ;
  assign n18 = ~n16 & n17 ;
  assign n19 = x7 & ~x9 ;
  assign n20 = ~x5 & n19 ;
  assign n21 = n20 ^ x9 ;
  assign n22 = n18 & n21 ;
  assign n23 = ~x2 & ~x8 ;
  assign n24 = ~x1 & ~n23 ;
  assign n25 = x6 & x14 ;
  assign n26 = x0 & ~x3 ;
  assign n27 = n25 & n26 ;
  assign n28 = ~n24 & n27 ;
  assign n29 = n22 & n28 ;
  assign n30 = x2 & x7 ;
  assign n31 = n30 ^ x5 ;
  assign n32 = ~x9 & n30 ;
  assign n33 = n31 & n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n29 & ~n34 ;
  assign n36 = ~x10 & n16 ;
  assign n37 = x4 & n30 ;
  assign n38 = x8 & ~x9 ;
  assign n39 = ~x1 & ~n38 ;
  assign n40 = n37 & n39 ;
  assign n41 = ~n36 & n40 ;
  assign n42 = ~x7 & x9 ;
  assign n43 = x2 & n42 ;
  assign n44 = x1 & ~n43 ;
  assign n45 = x8 & ~n44 ;
  assign n46 = n45 ^ n19 ;
  assign n47 = n46 ^ n17 ;
  assign n48 = n42 ^ x2 ;
  assign n49 = n19 & ~n48 ;
  assign n50 = n49 ^ n42 ;
  assign n51 = n47 & n50 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = n52 ^ n42 ;
  assign n54 = n53 ^ n19 ;
  assign n55 = n17 & n54 ;
  assign n56 = ~n41 & ~n55 ;
  assign n57 = ~x5 & n25 ;
  assign n58 = ~n56 & n57 ;
  assign n59 = x0 & ~n58 ;
  assign n60 = ~x6 & ~x14 ;
  assign n61 = ~x10 & n60 ;
  assign n62 = ~n30 & ~n61 ;
  assign n63 = x5 & ~x9 ;
  assign n64 = ~x1 & ~x4 ;
  assign n65 = x2 & ~n25 ;
  assign n66 = n64 & ~n65 ;
  assign n67 = n66 ^ x2 ;
  assign n68 = n67 ^ n66 ;
  assign n69 = x1 & x4 ;
  assign n70 = n69 ^ n66 ;
  assign n71 = n70 ^ n66 ;
  assign n72 = ~n68 & n71 ;
  assign n73 = n72 ^ n66 ;
  assign n74 = ~x7 & n73 ;
  assign n75 = n74 ^ n66 ;
  assign n76 = n63 & n75 ;
  assign n77 = ~n62 & n76 ;
  assign n78 = x6 & x10 ;
  assign n79 = ~x14 & n69 ;
  assign n80 = n43 & n79 ;
  assign n81 = ~n78 & n80 ;
  assign n82 = ~n77 & ~n81 ;
  assign n83 = ~x8 & ~n82 ;
  assign n84 = x8 & x10 ;
  assign n85 = ~x2 & n19 ;
  assign n86 = n69 & n85 ;
  assign n87 = n84 & n86 ;
  assign n88 = ~x0 & ~n87 ;
  assign n89 = n57 & ~n88 ;
  assign n97 = ~x2 & ~x7 ;
  assign n98 = n61 & n97 ;
  assign n90 = x7 & x10 ;
  assign n91 = x6 & ~n90 ;
  assign n92 = x2 & n79 ;
  assign n93 = n16 & n92 ;
  assign n94 = ~n91 & n93 ;
  assign n99 = n98 ^ n94 ;
  assign n100 = n99 ^ n94 ;
  assign n95 = n94 ^ n64 ;
  assign n96 = n95 ^ n94 ;
  assign n101 = n100 ^ n96 ;
  assign n102 = n94 ^ n38 ;
  assign n103 = n102 ^ n94 ;
  assign n104 = n103 ^ n100 ;
  assign n105 = n100 & n104 ;
  assign n106 = n105 ^ n100 ;
  assign n107 = n101 & n106 ;
  assign n108 = n107 ^ n105 ;
  assign n109 = n108 ^ n94 ;
  assign n110 = n109 ^ n100 ;
  assign n111 = x5 & n110 ;
  assign n112 = n111 ^ n94 ;
  assign n113 = ~n89 & ~n112 ;
  assign n114 = ~n83 & n113 ;
  assign n115 = x3 & ~n114 ;
  assign n116 = ~n59 & n115 ;
  assign n117 = ~n35 & ~n116 ;
  assign n118 = ~x12 & ~x13 ;
  assign n119 = ~x11 & n118 ;
  assign n120 = ~n117 & n119 ;
  assign y0 = n120 ;
endmodule
