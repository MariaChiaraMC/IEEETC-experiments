module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 ;
  assign n16 = ~x3 & x4 ;
  assign n17 = x1 ^ x0 ;
  assign n18 = ~x10 & ~x11 ;
  assign n19 = x13 ^ x12 ;
  assign n20 = n19 ^ x14 ;
  assign n21 = n20 ^ x12 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = x14 ^ x7 ;
  assign n24 = ~x12 & n23 ;
  assign n25 = n24 ^ x14 ;
  assign n26 = ~n22 & ~n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n27 ^ x14 ;
  assign n29 = n28 ^ x12 ;
  assign n30 = n18 & n29 ;
  assign n31 = n30 ^ x7 ;
  assign n32 = x9 ^ x8 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = ~x13 & ~x14 ;
  assign n36 = ~x12 & n35 ;
  assign n37 = n36 ^ x8 ;
  assign n38 = ~n30 & ~n37 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n34 & n39 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n41 ^ n36 ;
  assign n43 = n42 ^ n30 ;
  assign n44 = ~n31 & ~n43 ;
  assign n45 = n44 ^ x7 ;
  assign n46 = ~x6 & n45 ;
  assign n47 = ~x2 & ~x5 ;
  assign n48 = ~n46 & n47 ;
  assign n49 = x1 & ~n48 ;
  assign n50 = n17 & n49 ;
  assign n51 = n50 ^ n17 ;
  assign n52 = n16 & n51 ;
  assign y0 = n52 ;
endmodule
