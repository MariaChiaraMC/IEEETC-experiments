module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 ;
  assign n16 = ~x11 & ~x12 ;
  assign n17 = x6 & ~x10 ;
  assign n22 = x5 & x7 ;
  assign n23 = x3 & ~x4 ;
  assign n24 = n22 & n23 ;
  assign n18 = ~x3 & ~x4 ;
  assign n19 = ~x7 & ~x8 ;
  assign n20 = ~x5 & n19 ;
  assign n21 = n18 & n20 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = ~x8 & ~x9 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = n28 ^ n21 ;
  assign n30 = n26 & n29 ;
  assign n31 = n30 ^ n21 ;
  assign n32 = x13 & n31 ;
  assign n33 = n32 ^ n21 ;
  assign n34 = n17 & n33 ;
  assign n35 = ~x6 & x10 ;
  assign n36 = x5 & n35 ;
  assign n37 = x13 ^ x3 ;
  assign n39 = ~x7 & ~x9 ;
  assign n38 = ~x8 & x9 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = n39 ^ x13 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = n40 & n42 ;
  assign n44 = n43 ^ n39 ;
  assign n45 = n37 & n44 ;
  assign n46 = n36 & n45 ;
  assign n47 = x4 & n46 ;
  assign n48 = ~n34 & ~n47 ;
  assign n49 = ~x0 & x2 ;
  assign n50 = ~x14 & n49 ;
  assign n51 = ~n48 & n50 ;
  assign n52 = n51 ^ x1 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n53 ^ n16 ;
  assign n55 = x0 & x6 ;
  assign n56 = ~x2 & x3 ;
  assign n57 = ~n38 & ~n56 ;
  assign n58 = ~n39 & n57 ;
  assign n59 = ~x13 & ~x14 ;
  assign n60 = ~x10 & n59 ;
  assign n61 = x2 & x9 ;
  assign n62 = x7 & n61 ;
  assign n63 = ~x4 & ~n62 ;
  assign n64 = n60 & n63 ;
  assign n65 = n58 & n64 ;
  assign n66 = ~x2 & x7 ;
  assign n67 = x3 & x4 ;
  assign n68 = x13 & n67 ;
  assign n69 = n66 & n68 ;
  assign n70 = x14 & n69 ;
  assign n71 = ~n65 & ~n70 ;
  assign n72 = n55 & ~n71 ;
  assign n73 = n38 & n49 ;
  assign n74 = n67 & n73 ;
  assign n75 = x14 ^ x6 ;
  assign n76 = n75 ^ x13 ;
  assign n77 = n76 ^ x14 ;
  assign n78 = n77 ^ n76 ;
  assign n79 = x10 ^ x7 ;
  assign n80 = n79 ^ n76 ;
  assign n81 = n80 ^ n75 ;
  assign n82 = ~n78 & n81 ;
  assign n83 = n82 ^ n79 ;
  assign n84 = x10 & ~n79 ;
  assign n85 = n84 ^ n75 ;
  assign n86 = ~n83 & n85 ;
  assign n87 = n86 ^ n84 ;
  assign n88 = n75 & n87 ;
  assign n89 = n88 ^ n82 ;
  assign n90 = n89 ^ x6 ;
  assign n91 = n90 ^ n79 ;
  assign n92 = n74 & n91 ;
  assign n93 = ~n72 & ~n92 ;
  assign n94 = ~x5 & ~n93 ;
  assign n95 = x6 & x10 ;
  assign n96 = n19 & ~n95 ;
  assign n97 = ~x0 & n68 ;
  assign n98 = n96 & n97 ;
  assign n99 = x8 & n60 ;
  assign n100 = n18 & n22 ;
  assign n101 = n99 & n100 ;
  assign n102 = n55 & n101 ;
  assign n103 = ~n98 & ~n102 ;
  assign n104 = n61 & ~n103 ;
  assign n105 = n104 ^ n94 ;
  assign n106 = ~n94 & n105 ;
  assign n107 = n106 ^ n51 ;
  assign n108 = n107 ^ n94 ;
  assign n109 = n54 & n108 ;
  assign n110 = n109 ^ n106 ;
  assign n111 = n110 ^ n94 ;
  assign n112 = n16 & ~n111 ;
  assign n113 = n112 ^ n16 ;
  assign y0 = n113 ;
endmodule
