module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 ;
  output y0 ;
  wire n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 ;
  assign n22 = ~x0 & ~x1 ;
  assign n23 = x2 & ~n22 ;
  assign n27 = x1 ^ x0 ;
  assign n37 = ~n23 & ~n27 ;
  assign n38 = x7 & n37 ;
  assign n39 = x3 & n23 ;
  assign n19 = ~x2 & ~x5 ;
  assign n20 = ~x4 & n19 ;
  assign n40 = x6 & n20 ;
  assign n41 = ~n39 & ~n40 ;
  assign n42 = ~n38 & n41 ;
  assign n21 = x9 & n20 ;
  assign n24 = n23 ^ x8 ;
  assign n25 = n24 ^ x8 ;
  assign n26 = n25 ^ n21 ;
  assign n28 = n27 ^ x10 ;
  assign n29 = ~n27 & ~n28 ;
  assign n30 = n29 ^ x8 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n26 & ~n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = ~n21 & ~n34 ;
  assign n36 = n35 ^ n21 ;
  assign n43 = n42 ^ n36 ;
  assign n44 = n42 ^ x13 ;
  assign n45 = n44 ^ n43 ;
  assign n51 = x14 & ~x15 ;
  assign n52 = ~x16 & ~n51 ;
  assign n53 = ~x11 & ~n52 ;
  assign n54 = ~x17 & ~n53 ;
  assign n55 = ~x12 & ~n54 ;
  assign n46 = ~x14 & x15 ;
  assign n47 = x16 & ~n46 ;
  assign n48 = x11 & ~n47 ;
  assign n49 = x17 & ~n48 ;
  assign n50 = x12 & ~n49 ;
  assign n56 = n55 ^ n50 ;
  assign n57 = ~x13 & n56 ;
  assign n58 = n57 ^ n50 ;
  assign n59 = ~n45 & n58 ;
  assign n60 = n59 ^ n57 ;
  assign n61 = n60 ^ n50 ;
  assign n62 = n61 ^ x13 ;
  assign n63 = ~n43 & ~n62 ;
  assign n64 = n63 ^ n36 ;
  assign y0 = n64 ;
endmodule
