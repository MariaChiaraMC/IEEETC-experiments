module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 ;
  assign n22 = x1 ^ x0 ;
  assign n23 = x2 ^ x1 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = x5 ^ x3 ;
  assign n27 = x5 ^ x1 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = ~n26 & ~n28 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = n30 ^ n26 ;
  assign n32 = n25 & ~n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ n26 ;
  assign n35 = n22 & ~n34 ;
  assign n36 = ~x4 & n35 ;
  assign n37 = ~x19 & ~x20 ;
  assign n38 = n37 ^ x18 ;
  assign n39 = n38 ^ x18 ;
  assign n40 = ~x12 & ~x13 ;
  assign n42 = ~x6 & ~x7 ;
  assign n43 = ~x8 & n42 ;
  assign n44 = ~x11 & n43 ;
  assign n63 = x10 & n44 ;
  assign n41 = ~x0 & ~x2 ;
  assign n45 = ~x10 & x11 ;
  assign n46 = x8 & n45 ;
  assign n47 = n42 & n46 ;
  assign n48 = ~n44 & ~n47 ;
  assign n49 = n41 & ~n48 ;
  assign n50 = ~x2 & x3 ;
  assign n51 = ~x1 & n50 ;
  assign n52 = x8 & x10 ;
  assign n53 = ~n43 & ~n52 ;
  assign n54 = n51 & ~n53 ;
  assign n55 = ~x11 & n54 ;
  assign n56 = ~x5 & ~n55 ;
  assign n57 = ~x11 & n52 ;
  assign n58 = ~x10 & ~n48 ;
  assign n59 = x2 & ~n58 ;
  assign n60 = ~n57 & n59 ;
  assign n61 = ~n56 & ~n60 ;
  assign n62 = ~n49 & ~n61 ;
  assign n64 = n63 ^ n62 ;
  assign n65 = n64 ^ x9 ;
  assign n73 = n65 ^ n64 ;
  assign n66 = ~x1 & n41 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = n67 ^ n64 ;
  assign n69 = n65 ^ n62 ;
  assign n70 = n69 ^ n66 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = ~n68 & ~n71 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = n74 ^ n68 ;
  assign n76 = n64 ^ x5 ;
  assign n77 = n72 ^ n68 ;
  assign n78 = n76 & ~n77 ;
  assign n79 = n78 ^ n64 ;
  assign n80 = ~n75 & ~n79 ;
  assign n81 = n80 ^ n64 ;
  assign n82 = n81 ^ n63 ;
  assign n83 = n82 ^ n64 ;
  assign n84 = n40 & n83 ;
  assign n85 = x5 & ~x9 ;
  assign n86 = ~x8 & n45 ;
  assign n87 = n85 & n86 ;
  assign n88 = x12 & ~x13 ;
  assign n89 = ~x13 & ~n42 ;
  assign n90 = ~n88 & ~n89 ;
  assign n91 = n87 & n90 ;
  assign n92 = ~x5 & ~n41 ;
  assign n93 = ~x3 & ~n92 ;
  assign n94 = ~n91 & ~n93 ;
  assign n95 = ~n84 & n94 ;
  assign n96 = ~x4 & ~n95 ;
  assign n97 = x5 ^ x0 ;
  assign n98 = n97 ^ x3 ;
  assign n99 = n98 ^ x3 ;
  assign n101 = x5 ^ x2 ;
  assign n100 = n99 ^ n98 ;
  assign n102 = n101 ^ n100 ;
  assign n103 = ~n99 & n102 ;
  assign n104 = n103 ^ n98 ;
  assign n105 = n104 ^ n99 ;
  assign n109 = n99 ^ x4 ;
  assign n110 = ~n99 & n109 ;
  assign n106 = n98 ^ x5 ;
  assign n107 = n106 ^ n99 ;
  assign n108 = ~x13 & n107 ;
  assign n111 = n110 ^ n108 ;
  assign n112 = n111 ^ n98 ;
  assign n113 = n112 ^ x5 ;
  assign n114 = n113 ^ n99 ;
  assign n115 = n114 ^ n101 ;
  assign n116 = ~x5 & ~n115 ;
  assign n117 = n116 ^ n108 ;
  assign n118 = n117 ^ n98 ;
  assign n119 = n118 ^ n99 ;
  assign n120 = n119 ^ n101 ;
  assign n121 = ~n105 & n120 ;
  assign n122 = n121 ^ n108 ;
  assign n123 = n122 ^ n103 ;
  assign n124 = n123 ^ n116 ;
  assign n125 = n124 ^ n101 ;
  assign n126 = n125 ^ x5 ;
  assign n127 = x3 & ~x5 ;
  assign n128 = n127 ^ x4 ;
  assign n129 = n128 ^ n127 ;
  assign n130 = n129 ^ n126 ;
  assign n131 = ~x3 & n40 ;
  assign n132 = ~x9 & ~n63 ;
  assign n133 = x2 & ~n132 ;
  assign n134 = n131 & n133 ;
  assign n135 = n48 & ~n57 ;
  assign n136 = n135 ^ n134 ;
  assign n137 = n134 & ~n136 ;
  assign n138 = n137 ^ n127 ;
  assign n139 = n138 ^ n134 ;
  assign n140 = n130 & n139 ;
  assign n141 = n140 ^ n137 ;
  assign n142 = n141 ^ n134 ;
  assign n143 = ~n126 & n142 ;
  assign n144 = n143 ^ n126 ;
  assign n145 = x1 & n144 ;
  assign n146 = ~x1 & ~x3 ;
  assign n147 = ~n127 & ~n146 ;
  assign n148 = x4 & ~n147 ;
  assign n149 = n86 & n146 ;
  assign n150 = n149 ^ x4 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = ~x1 & n40 ;
  assign n153 = n47 & n152 ;
  assign n154 = ~n53 & n131 ;
  assign n155 = ~x11 & n154 ;
  assign n156 = ~n153 & ~n155 ;
  assign n157 = n156 ^ n149 ;
  assign n158 = n157 ^ n149 ;
  assign n159 = ~n151 & ~n158 ;
  assign n160 = n159 ^ n149 ;
  assign n161 = x9 & n160 ;
  assign n162 = n161 ^ n149 ;
  assign n163 = x2 & n162 ;
  assign n164 = n127 & n153 ;
  assign n165 = x9 & n164 ;
  assign n166 = ~n163 & ~n165 ;
  assign n167 = ~n148 & n166 ;
  assign n168 = x0 & ~n167 ;
  assign n173 = x12 ^ x11 ;
  assign n177 = n173 ^ x12 ;
  assign n169 = x1 & x11 ;
  assign n170 = ~x8 & ~n169 ;
  assign n171 = n170 ^ x10 ;
  assign n172 = n171 ^ n170 ;
  assign n174 = n173 ^ n170 ;
  assign n175 = n174 ^ x12 ;
  assign n176 = ~n172 & n175 ;
  assign n178 = n177 ^ n176 ;
  assign n179 = n178 ^ x9 ;
  assign n180 = x13 ^ x12 ;
  assign n181 = n177 ^ x9 ;
  assign n182 = ~n180 & ~n181 ;
  assign n183 = n182 ^ n176 ;
  assign n184 = n183 ^ x12 ;
  assign n185 = n184 ^ n180 ;
  assign n186 = n185 ^ n177 ;
  assign n187 = x9 & ~n186 ;
  assign n188 = ~n179 & n187 ;
  assign n189 = ~x2 & ~n188 ;
  assign n190 = x16 & ~x17 ;
  assign n191 = ~x9 & ~n88 ;
  assign n192 = n86 & n191 ;
  assign n193 = n190 & n192 ;
  assign n194 = n42 & n193 ;
  assign n195 = ~n189 & ~n194 ;
  assign n196 = x12 ^ x2 ;
  assign n197 = n196 ^ x12 ;
  assign n198 = x15 ^ x12 ;
  assign n199 = n197 & ~n198 ;
  assign n200 = n199 ^ x12 ;
  assign n201 = x13 & ~n200 ;
  assign n202 = ~n195 & ~n201 ;
  assign n203 = ~x3 & ~n202 ;
  assign n204 = ~n51 & ~n203 ;
  assign n205 = x5 & ~n204 ;
  assign n206 = ~n168 & ~n205 ;
  assign n207 = ~n145 & n206 ;
  assign n208 = ~n96 & n207 ;
  assign n209 = n208 ^ x18 ;
  assign n210 = n39 & n209 ;
  assign n211 = n210 ^ x18 ;
  assign n212 = x14 & n211 ;
  assign n213 = ~n36 & n212 ;
  assign y0 = ~n213 ;
endmodule
