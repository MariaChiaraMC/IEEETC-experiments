module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 ;
  assign n13 = x0 & x1 ;
  assign n14 = x6 ^ x5 ;
  assign n15 = x8 & x9 ;
  assign n16 = x4 & ~x10 ;
  assign n17 = x7 & n16 ;
  assign n18 = n15 & n17 ;
  assign n19 = ~x2 & n18 ;
  assign n20 = ~x4 & ~x10 ;
  assign n21 = x2 & x3 ;
  assign n22 = ~n20 & n21 ;
  assign n23 = ~x7 & ~x8 ;
  assign n24 = ~n22 & n23 ;
  assign n25 = x9 & n24 ;
  assign n28 = n15 ^ x4 ;
  assign n32 = n28 ^ n15 ;
  assign n26 = x3 ^ x2 ;
  assign n27 = n26 ^ x2 ;
  assign n29 = n28 ^ x2 ;
  assign n30 = n29 ^ n15 ;
  assign n31 = n27 & ~n30 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = n33 ^ x7 ;
  assign n35 = n15 ^ x8 ;
  assign n36 = n32 ^ x7 ;
  assign n37 = ~n35 & n36 ;
  assign n38 = n37 ^ n31 ;
  assign n39 = n38 ^ n15 ;
  assign n40 = n39 ^ n35 ;
  assign n41 = n40 ^ n32 ;
  assign n42 = x7 & ~n41 ;
  assign n43 = n34 & n42 ;
  assign n44 = ~n25 & ~n43 ;
  assign n45 = ~x11 & ~n44 ;
  assign n46 = ~n19 & ~n45 ;
  assign n47 = n46 ^ x6 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = n48 ^ n14 ;
  assign n50 = x2 & ~x11 ;
  assign n51 = ~x3 & n50 ;
  assign n52 = n51 ^ n18 ;
  assign n53 = n51 & n52 ;
  assign n54 = n53 ^ n46 ;
  assign n55 = n54 ^ n51 ;
  assign n56 = n49 & ~n55 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n57 ^ n51 ;
  assign n59 = n14 & n58 ;
  assign n60 = n13 & n59 ;
  assign y0 = n60 ;
endmodule
