module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n10 = x7 ^ x4 ;
  assign n11 = x7 ^ x5 ;
  assign n12 = n11 ^ x5 ;
  assign n13 = x8 ^ x5 ;
  assign n14 = n12 & ~n13 ;
  assign n15 = n14 ^ x5 ;
  assign n16 = ~n10 & ~n15 ;
  assign n17 = n16 ^ x4 ;
  assign n18 = x6 & ~n17 ;
  assign n19 = x7 & x8 ;
  assign n20 = ~x6 & ~n19 ;
  assign n21 = ~x0 & ~n20 ;
  assign n22 = x4 ^ x3 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = ~x1 & x2 ;
  assign n25 = ~x8 & n24 ;
  assign n26 = ~x3 & n25 ;
  assign n27 = n26 ^ n21 ;
  assign n28 = n23 & n27 ;
  assign n29 = n28 ^ n26 ;
  assign n30 = n21 & n29 ;
  assign n31 = ~n18 & n30 ;
  assign y0 = n31 ;
endmodule
