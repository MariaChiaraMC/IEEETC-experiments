module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n9 = x6 ^ x4 ;
  assign n13 = n9 ^ x7 ;
  assign n11 = x7 ^ x5 ;
  assign n10 = n9 ^ x6 ;
  assign n12 = n11 ^ n10 ;
  assign n14 = n13 ^ n12 ;
  assign n17 = x6 ^ x2 ;
  assign n18 = n17 ^ x7 ;
  assign n19 = n18 ^ n11 ;
  assign n20 = n19 ^ n13 ;
  assign n21 = ~n13 & n20 ;
  assign n15 = n9 & ~n11 ;
  assign n24 = n21 ^ n15 ;
  assign n16 = n15 ^ n14 ;
  assign n22 = n21 ^ n13 ;
  assign n23 = ~n16 & ~n22 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = ~n14 & n25 ;
  assign n27 = n26 ^ n21 ;
  assign n28 = n27 ^ n23 ;
  assign n29 = n28 ^ n18 ;
  assign n30 = ~x3 & n29 ;
  assign n31 = ~x1 & ~n30 ;
  assign n32 = ~x0 & ~n31 ;
  assign y0 = n32 ;
endmodule
