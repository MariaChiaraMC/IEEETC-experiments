module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 ;
  assign n11 = ~x2 & ~x3 ;
  assign n12 = x6 & x7 ;
  assign n13 = x8 & n12 ;
  assign n14 = n11 & n13 ;
  assign n15 = x2 & x3 ;
  assign n16 = ~x6 & ~x8 ;
  assign n17 = ~x7 & n16 ;
  assign n18 = n15 & n17 ;
  assign n19 = ~n14 & ~n18 ;
  assign n20 = x0 & x4 ;
  assign n21 = x5 & n20 ;
  assign n22 = ~n19 & n21 ;
  assign n23 = ~x9 & n22 ;
  assign n24 = x8 & ~x9 ;
  assign n25 = ~x5 & x6 ;
  assign n26 = ~x7 & n25 ;
  assign n27 = ~x2 & x3 ;
  assign n28 = ~x0 & ~x4 ;
  assign n29 = n27 & n28 ;
  assign n30 = n26 & n29 ;
  assign n31 = n24 & n30 ;
  assign n32 = n31 ^ n23 ;
  assign n33 = ~x7 & x9 ;
  assign n34 = x6 & x8 ;
  assign n35 = x4 & n34 ;
  assign n37 = ~x2 & x5 ;
  assign n36 = x2 & ~x5 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = ~x0 & n38 ;
  assign n40 = n39 ^ n37 ;
  assign n41 = n35 & n40 ;
  assign n42 = n33 & n41 ;
  assign n43 = x0 & ~x4 ;
  assign n44 = ~x6 & ~x9 ;
  assign n45 = n36 & n44 ;
  assign n46 = n43 & n45 ;
  assign n47 = ~x8 & n46 ;
  assign n85 = ~x8 & ~x9 ;
  assign n86 = n36 & n85 ;
  assign n79 = x5 & x6 ;
  assign n49 = ~x2 & ~x8 ;
  assign n87 = ~x9 & ~n49 ;
  assign n88 = n79 & ~n87 ;
  assign n89 = ~n86 & ~n88 ;
  assign n90 = n89 ^ x9 ;
  assign n78 = x2 & ~x8 ;
  assign n91 = n89 ^ n78 ;
  assign n92 = n91 ^ n78 ;
  assign n93 = n92 ^ n90 ;
  assign n94 = x5 & ~x6 ;
  assign n95 = x2 & n94 ;
  assign n96 = n95 ^ x8 ;
  assign n97 = n95 & n96 ;
  assign n98 = n97 ^ n78 ;
  assign n99 = n98 ^ n95 ;
  assign n100 = n93 & ~n99 ;
  assign n101 = n100 ^ n97 ;
  assign n102 = n101 ^ n95 ;
  assign n103 = n90 & n102 ;
  assign n104 = n103 ^ n89 ;
  assign n105 = n43 & ~n104 ;
  assign n48 = x4 & ~x6 ;
  assign n50 = n49 ^ n48 ;
  assign n51 = ~x4 & x6 ;
  assign n52 = n51 ^ n48 ;
  assign n53 = n49 ^ x9 ;
  assign n54 = n53 ^ n48 ;
  assign n55 = ~n48 & n54 ;
  assign n56 = n55 ^ n48 ;
  assign n57 = ~n52 & ~n56 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = n58 ^ n48 ;
  assign n60 = n59 ^ n53 ;
  assign n61 = ~n50 & n60 ;
  assign n62 = n61 ^ n48 ;
  assign n63 = x5 & n62 ;
  assign n64 = x5 & ~n51 ;
  assign n65 = x2 & n24 ;
  assign n66 = ~n64 & ~n65 ;
  assign n67 = x0 & ~n66 ;
  assign n68 = x5 & ~x9 ;
  assign n69 = x5 & x8 ;
  assign n70 = ~n48 & ~n69 ;
  assign n71 = ~n68 & n70 ;
  assign n72 = n67 & ~n71 ;
  assign n73 = ~n63 & n72 ;
  assign n74 = ~x5 & ~x6 ;
  assign n75 = ~x2 & x8 ;
  assign n76 = ~n74 & ~n75 ;
  assign n77 = ~x0 & x4 ;
  assign n80 = ~n78 & ~n79 ;
  assign n81 = n77 & ~n80 ;
  assign n82 = ~n76 & n81 ;
  assign n83 = ~x9 & n82 ;
  assign n84 = ~n73 & ~n83 ;
  assign n106 = n105 ^ n84 ;
  assign n107 = n106 ^ n84 ;
  assign n117 = ~x5 & x9 ;
  assign n118 = ~n79 & ~n117 ;
  assign n114 = x2 & x8 ;
  assign n108 = ~x8 & n37 ;
  assign n115 = n114 ^ n108 ;
  assign n119 = n118 ^ n115 ;
  assign n120 = n119 ^ n115 ;
  assign n110 = x9 ^ x6 ;
  assign n109 = n108 ^ x9 ;
  assign n111 = n110 ^ n109 ;
  assign n112 = n111 ^ n110 ;
  assign n113 = n112 ^ x9 ;
  assign n116 = n115 ^ n113 ;
  assign n121 = n120 ^ n116 ;
  assign n124 = n113 ^ x9 ;
  assign n122 = n110 ^ x9 ;
  assign n123 = n122 ^ n116 ;
  assign n125 = n124 ^ n123 ;
  assign n126 = ~n121 & n125 ;
  assign n127 = n126 ^ n113 ;
  assign n128 = n127 ^ n122 ;
  assign n129 = n128 ^ n124 ;
  assign n130 = n123 ^ n120 ;
  assign n131 = n127 & ~n130 ;
  assign n132 = n131 ^ n113 ;
  assign n133 = n132 ^ n116 ;
  assign n134 = n133 ^ n120 ;
  assign n135 = n129 & ~n134 ;
  assign n136 = n135 ^ n108 ;
  assign n137 = n77 & n136 ;
  assign n138 = ~n51 & ~n75 ;
  assign n139 = n117 & ~n138 ;
  assign n140 = ~n34 & n139 ;
  assign n141 = ~x0 & n140 ;
  assign n142 = ~n137 & ~n141 ;
  assign n143 = n142 ^ n84 ;
  assign n144 = n143 ^ n84 ;
  assign n145 = ~n107 & n144 ;
  assign n146 = n145 ^ n84 ;
  assign n147 = x7 & n146 ;
  assign n148 = n147 ^ n84 ;
  assign n149 = ~n47 & n148 ;
  assign n150 = n149 ^ x3 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = x6 ^ x0 ;
  assign n160 = n152 ^ x6 ;
  assign n154 = x6 ^ x5 ;
  assign n158 = n154 ^ x7 ;
  assign n161 = n160 ^ n158 ;
  assign n162 = n161 ^ n158 ;
  assign n153 = n152 ^ x9 ;
  assign n155 = n154 ^ n153 ;
  assign n156 = n155 ^ n154 ;
  assign n157 = n156 ^ n152 ;
  assign n159 = n158 ^ n157 ;
  assign n163 = n162 ^ n159 ;
  assign n166 = n157 ^ n152 ;
  assign n164 = n154 ^ n152 ;
  assign n165 = n164 ^ n159 ;
  assign n167 = n166 ^ n165 ;
  assign n168 = ~n163 & n167 ;
  assign n169 = n168 ^ n157 ;
  assign n170 = n169 ^ n164 ;
  assign n171 = n170 ^ n166 ;
  assign n172 = n165 ^ n162 ;
  assign n173 = ~n169 & ~n172 ;
  assign n174 = n173 ^ n157 ;
  assign n175 = n174 ^ n159 ;
  assign n176 = n175 ^ n162 ;
  assign n177 = ~n171 & n176 ;
  assign n178 = n75 & n177 ;
  assign n179 = ~x4 & n178 ;
  assign n180 = ~x7 & n44 ;
  assign n181 = ~x0 & n180 ;
  assign n182 = n37 & n181 ;
  assign n183 = n12 & n77 ;
  assign n184 = x0 & ~x6 ;
  assign n185 = x7 ^ x4 ;
  assign n186 = n184 & n185 ;
  assign n187 = ~n183 & ~n186 ;
  assign n188 = ~x2 & n117 ;
  assign n189 = ~n187 & n188 ;
  assign n190 = x6 & x9 ;
  assign n191 = x5 & n190 ;
  assign n192 = ~n45 & ~n191 ;
  assign n193 = n28 & ~n192 ;
  assign n194 = ~x7 & n193 ;
  assign n195 = ~n189 & ~n194 ;
  assign n196 = ~n182 & n195 ;
  assign n197 = n196 ^ x8 ;
  assign n198 = n197 ^ n196 ;
  assign n199 = n198 ^ n179 ;
  assign n216 = ~x0 & n74 ;
  assign n217 = x4 & ~n79 ;
  assign n218 = ~n216 & ~n217 ;
  assign n203 = x5 & ~n44 ;
  assign n204 = x4 & n203 ;
  assign n200 = ~x9 & ~n51 ;
  assign n201 = ~n74 & ~n79 ;
  assign n202 = n200 & n201 ;
  assign n205 = n204 ^ n202 ;
  assign n206 = n205 ^ n202 ;
  assign n207 = ~x5 & n190 ;
  assign n208 = n207 ^ n202 ;
  assign n209 = n208 ^ n202 ;
  assign n210 = ~n206 & ~n209 ;
  assign n211 = n210 ^ n202 ;
  assign n212 = ~x0 & ~n211 ;
  assign n213 = n212 ^ n202 ;
  assign n219 = n218 ^ n213 ;
  assign n220 = n219 ^ n213 ;
  assign n214 = n213 ^ n77 ;
  assign n215 = n214 ^ n213 ;
  assign n221 = n220 ^ n215 ;
  assign n222 = n213 ^ x9 ;
  assign n223 = n222 ^ n213 ;
  assign n224 = n223 ^ n220 ;
  assign n225 = ~n220 & ~n224 ;
  assign n226 = n225 ^ n220 ;
  assign n227 = n221 & ~n226 ;
  assign n228 = n227 ^ n225 ;
  assign n229 = n228 ^ n213 ;
  assign n230 = n229 ^ n220 ;
  assign n231 = x7 & ~n230 ;
  assign n232 = n231 ^ n213 ;
  assign n233 = n232 ^ x2 ;
  assign n234 = n232 & n233 ;
  assign n235 = n234 ^ n196 ;
  assign n236 = n235 ^ n232 ;
  assign n237 = ~n199 & ~n236 ;
  assign n238 = n237 ^ n234 ;
  assign n239 = n238 ^ n232 ;
  assign n240 = ~n179 & n239 ;
  assign n241 = n240 ^ n179 ;
  assign n242 = n241 ^ n149 ;
  assign n243 = n151 & ~n242 ;
  assign n244 = n243 ^ n149 ;
  assign n245 = ~n42 & n244 ;
  assign n246 = n245 ^ x1 ;
  assign n247 = n246 ^ n245 ;
  assign n271 = ~x3 & ~x5 ;
  assign n272 = n180 & n271 ;
  assign n273 = x3 & n203 ;
  assign n274 = ~n190 & n273 ;
  assign n275 = ~n272 & ~n274 ;
  assign n248 = x3 ^ x2 ;
  assign n249 = ~x2 & n25 ;
  assign n250 = n33 & n249 ;
  assign n251 = n250 ^ n248 ;
  assign n252 = x7 & ~x9 ;
  assign n253 = n74 & n252 ;
  assign n254 = ~n191 & ~n253 ;
  assign n255 = n254 ^ x2 ;
  assign n256 = n255 ^ n254 ;
  assign n257 = x7 & x9 ;
  assign n258 = n94 & n257 ;
  assign n259 = ~n26 & ~n258 ;
  assign n260 = n259 ^ n254 ;
  assign n261 = ~n256 & n260 ;
  assign n262 = n261 ^ n254 ;
  assign n263 = n262 ^ n248 ;
  assign n264 = n251 & n263 ;
  assign n265 = n264 ^ n261 ;
  assign n266 = n265 ^ n254 ;
  assign n267 = n266 ^ n250 ;
  assign n268 = ~n248 & n267 ;
  assign n269 = n268 ^ n248 ;
  assign n270 = n269 ^ n250 ;
  assign n276 = n275 ^ n270 ;
  assign n277 = n276 ^ n270 ;
  assign n278 = n270 ^ x2 ;
  assign n279 = n278 ^ n270 ;
  assign n280 = ~n277 & ~n279 ;
  assign n281 = n280 ^ n270 ;
  assign n282 = x8 & ~n281 ;
  assign n283 = n282 ^ n270 ;
  assign n284 = n77 & ~n283 ;
  assign n285 = x8 ^ x5 ;
  assign n286 = n252 ^ x8 ;
  assign n287 = n286 ^ n252 ;
  assign n288 = n252 ^ n33 ;
  assign n289 = ~n287 & n288 ;
  assign n290 = n289 ^ n252 ;
  assign n291 = ~n285 & n290 ;
  assign n292 = ~x2 & n291 ;
  assign n293 = n78 & n252 ;
  assign n294 = ~x0 & ~n293 ;
  assign n295 = x5 & ~n294 ;
  assign n296 = ~n292 & ~n295 ;
  assign n297 = n33 & n108 ;
  assign n298 = x0 & ~n297 ;
  assign n299 = ~x3 & x6 ;
  assign n300 = ~n298 & n299 ;
  assign n301 = ~n296 & n300 ;
  assign n302 = x9 ^ x3 ;
  assign n303 = n302 ^ x9 ;
  assign n304 = n68 ^ x9 ;
  assign n305 = ~n303 & n304 ;
  assign n306 = n305 ^ x9 ;
  assign n307 = n248 & n306 ;
  assign n308 = n17 & n307 ;
  assign n309 = n308 ^ x4 ;
  assign n310 = n309 ^ n308 ;
  assign n311 = n310 ^ n301 ;
  assign n313 = x3 & ~n117 ;
  assign n312 = n190 & n271 ;
  assign n314 = n313 ^ n312 ;
  assign n315 = n314 ^ x7 ;
  assign n323 = n315 ^ n314 ;
  assign n316 = ~x6 & ~x7 ;
  assign n317 = n316 ^ n315 ;
  assign n318 = n317 ^ n314 ;
  assign n319 = n315 ^ n312 ;
  assign n320 = n319 ^ n316 ;
  assign n321 = n320 ^ n318 ;
  assign n322 = ~n318 & ~n321 ;
  assign n324 = n323 ^ n322 ;
  assign n325 = n324 ^ n318 ;
  assign n326 = n314 ^ x9 ;
  assign n327 = n322 ^ n318 ;
  assign n328 = ~n326 & ~n327 ;
  assign n329 = n328 ^ n314 ;
  assign n330 = ~n325 & n329 ;
  assign n331 = n330 ^ n314 ;
  assign n332 = n331 ^ n313 ;
  assign n333 = n332 ^ n314 ;
  assign n334 = n78 & n333 ;
  assign n335 = n12 & n68 ;
  assign n336 = n335 ^ x7 ;
  assign n337 = n336 ^ n335 ;
  assign n338 = ~x6 & x9 ;
  assign n339 = ~n94 & ~n338 ;
  assign n340 = n339 ^ n335 ;
  assign n341 = n340 ^ n335 ;
  assign n342 = ~n337 & ~n341 ;
  assign n343 = n342 ^ n335 ;
  assign n344 = ~x3 & n343 ;
  assign n345 = n344 ^ n335 ;
  assign n346 = n114 & n345 ;
  assign n347 = x5 ^ x3 ;
  assign n348 = n347 ^ n75 ;
  assign n349 = n252 ^ x3 ;
  assign n350 = n349 ^ n252 ;
  assign n351 = n316 ^ n252 ;
  assign n352 = n350 & n351 ;
  assign n353 = n352 ^ n252 ;
  assign n354 = n353 ^ n347 ;
  assign n355 = n348 & n354 ;
  assign n356 = n355 ^ n352 ;
  assign n357 = n356 ^ n252 ;
  assign n358 = n357 ^ n75 ;
  assign n359 = n347 & n358 ;
  assign n360 = n359 ^ n347 ;
  assign n361 = ~n346 & ~n360 ;
  assign n362 = ~n334 & n361 ;
  assign n363 = n362 ^ x0 ;
  assign n364 = ~n362 & ~n363 ;
  assign n365 = n364 ^ n308 ;
  assign n366 = n365 ^ n362 ;
  assign n367 = ~n311 & ~n366 ;
  assign n368 = n367 ^ n364 ;
  assign n369 = n368 ^ n362 ;
  assign n370 = ~n301 & ~n369 ;
  assign n371 = n370 ^ n301 ;
  assign n372 = ~x7 & n85 ;
  assign n373 = n95 & n372 ;
  assign n374 = ~n13 & ~n17 ;
  assign n375 = x9 & ~n374 ;
  assign n376 = n375 ^ n252 ;
  assign n377 = n376 ^ x2 ;
  assign n384 = n377 ^ n376 ;
  assign n378 = n377 ^ n16 ;
  assign n379 = n378 ^ n376 ;
  assign n380 = n377 ^ n375 ;
  assign n381 = n380 ^ n16 ;
  assign n382 = n381 ^ n379 ;
  assign n383 = ~n379 & ~n382 ;
  assign n385 = n384 ^ n383 ;
  assign n386 = n385 ^ n379 ;
  assign n387 = n376 ^ n34 ;
  assign n388 = n383 ^ n379 ;
  assign n389 = ~n387 & ~n388 ;
  assign n390 = n389 ^ n376 ;
  assign n391 = ~n386 & n390 ;
  assign n392 = n391 ^ n376 ;
  assign n393 = n392 ^ n252 ;
  assign n394 = n393 ^ n376 ;
  assign n395 = n271 & n394 ;
  assign n396 = x3 & ~x6 ;
  assign n397 = ~x5 & ~x8 ;
  assign n398 = x7 & n397 ;
  assign n399 = n33 & n69 ;
  assign n400 = ~n398 & ~n399 ;
  assign n401 = n400 ^ x5 ;
  assign n402 = n401 ^ n400 ;
  assign n403 = x8 & n257 ;
  assign n404 = n403 ^ n400 ;
  assign n405 = n404 ^ n400 ;
  assign n406 = ~n402 & n405 ;
  assign n407 = n406 ^ n400 ;
  assign n408 = ~x2 & ~n407 ;
  assign n409 = n408 ^ n400 ;
  assign n410 = n396 & ~n409 ;
  assign n411 = ~n372 & ~n403 ;
  assign n412 = n27 & n79 ;
  assign n413 = ~n411 & n412 ;
  assign n414 = ~n410 & ~n413 ;
  assign n415 = ~n395 & n414 ;
  assign n416 = ~n373 & n415 ;
  assign n417 = n416 ^ x0 ;
  assign n418 = n417 ^ n416 ;
  assign n419 = ~n291 & ~n399 ;
  assign n420 = n15 & ~n419 ;
  assign n421 = ~x2 & ~x5 ;
  assign n422 = ~x7 & n24 ;
  assign n423 = x3 & n257 ;
  assign n424 = ~x8 & n423 ;
  assign n425 = ~n422 & ~n424 ;
  assign n426 = n421 & ~n425 ;
  assign n427 = ~n420 & ~n426 ;
  assign n428 = x6 & ~n427 ;
  assign n429 = n95 & n422 ;
  assign n430 = n396 ^ n37 ;
  assign n431 = n252 ^ x9 ;
  assign n432 = ~n287 & n431 ;
  assign n433 = n432 ^ n252 ;
  assign n434 = n433 ^ n396 ;
  assign n435 = n430 & n434 ;
  assign n436 = n435 ^ n432 ;
  assign n437 = n436 ^ n252 ;
  assign n438 = n437 ^ n37 ;
  assign n439 = n396 & n438 ;
  assign n440 = n439 ^ n396 ;
  assign n441 = ~n429 & ~n440 ;
  assign n442 = ~n428 & n441 ;
  assign n443 = n442 ^ n416 ;
  assign n444 = ~n418 & n443 ;
  assign n445 = n444 ^ n416 ;
  assign n446 = ~x4 & ~n445 ;
  assign n447 = ~n371 & ~n446 ;
  assign n448 = ~n284 & n447 ;
  assign n449 = n448 ^ n245 ;
  assign n450 = n247 & n449 ;
  assign n451 = n450 ^ n245 ;
  assign n452 = n451 ^ n23 ;
  assign n453 = n32 & ~n452 ;
  assign n454 = n453 ^ n450 ;
  assign n455 = n454 ^ n245 ;
  assign n456 = n455 ^ n31 ;
  assign n457 = ~n23 & ~n456 ;
  assign n458 = n457 ^ n23 ;
  assign y0 = n458 ;
endmodule
