module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 ;
  assign n11 = ~x2 & x5 ;
  assign n12 = ~x7 & x9 ;
  assign n13 = ~x6 & n12 ;
  assign n14 = ~x1 & n13 ;
  assign n15 = ~x3 & ~x4 ;
  assign n16 = ~x0 & n15 ;
  assign n17 = n14 & n16 ;
  assign n18 = n11 & n17 ;
  assign n142 = x0 & ~x1 ;
  assign n89 = x5 & ~x7 ;
  assign n143 = x2 & ~n89 ;
  assign n144 = ~x3 & n143 ;
  assign n145 = x5 ^ x4 ;
  assign n146 = n145 ^ x5 ;
  assign n147 = n146 ^ n144 ;
  assign n148 = n12 ^ x5 ;
  assign n149 = ~n147 & n148 ;
  assign n150 = n149 ^ n12 ;
  assign n151 = n144 & n150 ;
  assign n152 = x5 ^ x2 ;
  assign n153 = x3 & ~x9 ;
  assign n154 = ~x2 & x4 ;
  assign n155 = n154 ^ x7 ;
  assign n156 = n155 ^ n154 ;
  assign n157 = n156 ^ n153 ;
  assign n19 = x4 & x5 ;
  assign n158 = n154 ^ n19 ;
  assign n159 = ~n157 & ~n158 ;
  assign n160 = n159 ^ n19 ;
  assign n161 = n153 & n160 ;
  assign n162 = n152 & n161 ;
  assign n163 = ~n151 & ~n162 ;
  assign n164 = n142 & ~n163 ;
  assign n107 = x7 & ~x9 ;
  assign n165 = ~x3 & n107 ;
  assign n166 = n11 & n165 ;
  assign n167 = ~x1 & ~x5 ;
  assign n168 = ~x2 & x3 ;
  assign n169 = n107 & n168 ;
  assign n170 = ~x3 & ~x7 ;
  assign n171 = n170 ^ x9 ;
  assign n172 = n171 ^ x9 ;
  assign n173 = n172 ^ n169 ;
  assign n174 = x2 & x9 ;
  assign n175 = x3 & x7 ;
  assign n176 = n175 ^ n174 ;
  assign n177 = n174 & ~n176 ;
  assign n178 = n177 ^ x9 ;
  assign n179 = n178 ^ n174 ;
  assign n180 = n173 & ~n179 ;
  assign n181 = n180 ^ n177 ;
  assign n182 = n181 ^ n174 ;
  assign n183 = ~n169 & n182 ;
  assign n184 = n183 ^ n169 ;
  assign n185 = n167 & n184 ;
  assign n186 = ~n166 & ~n185 ;
  assign n187 = ~x0 & x4 ;
  assign n188 = ~n186 & n187 ;
  assign n189 = ~n164 & ~n188 ;
  assign n190 = x0 & x1 ;
  assign n38 = ~x2 & ~x4 ;
  assign n191 = ~x5 & x9 ;
  assign n192 = x3 & n191 ;
  assign n193 = n38 & n192 ;
  assign n194 = ~n170 & ~n175 ;
  assign n195 = n19 & ~n194 ;
  assign n196 = n12 ^ x9 ;
  assign n197 = ~x2 & ~n196 ;
  assign n198 = n197 ^ x9 ;
  assign n199 = n195 & ~n198 ;
  assign n200 = ~n193 & ~n199 ;
  assign n201 = n190 & ~n200 ;
  assign n202 = x1 & ~x3 ;
  assign n33 = ~x5 & ~x7 ;
  assign n203 = ~x9 & n33 ;
  assign n204 = n154 & n203 ;
  assign n205 = n202 & n204 ;
  assign n206 = x6 & ~n205 ;
  assign n207 = ~n201 & n206 ;
  assign n208 = ~x0 & x1 ;
  assign n91 = ~x5 & x7 ;
  assign n92 = ~x3 & n91 ;
  assign n209 = ~x2 & n92 ;
  assign n90 = x3 & n89 ;
  assign n210 = n38 & n90 ;
  assign n211 = ~n209 & ~n210 ;
  assign n212 = n211 ^ x9 ;
  assign n213 = n212 ^ n211 ;
  assign n80 = x3 & x5 ;
  assign n214 = ~n80 & n154 ;
  assign n108 = ~x4 & ~x5 ;
  assign n217 = n214 ^ n108 ;
  assign n218 = n217 ^ n214 ;
  assign n81 = ~x3 & x4 ;
  assign n82 = ~n80 & ~n81 ;
  assign n215 = n214 ^ n82 ;
  assign n216 = n215 ^ n214 ;
  assign n219 = n218 ^ n216 ;
  assign n220 = n214 ^ x2 ;
  assign n221 = n220 ^ n214 ;
  assign n222 = n221 ^ n218 ;
  assign n223 = ~n218 & ~n222 ;
  assign n224 = n223 ^ n218 ;
  assign n225 = ~n219 & ~n224 ;
  assign n226 = n225 ^ n223 ;
  assign n227 = n226 ^ n214 ;
  assign n228 = n227 ^ n218 ;
  assign n229 = x7 & ~n228 ;
  assign n230 = n229 ^ n214 ;
  assign n231 = n230 ^ n211 ;
  assign n232 = ~n213 & ~n231 ;
  assign n233 = n232 ^ n211 ;
  assign n234 = n208 & ~n233 ;
  assign n235 = n207 & ~n234 ;
  assign n236 = n189 & n235 ;
  assign n237 = x2 & ~x4 ;
  assign n238 = n203 ^ x1 ;
  assign n239 = n238 ^ n203 ;
  assign n240 = n239 ^ x0 ;
  assign n241 = ~x9 & n89 ;
  assign n242 = n241 ^ n91 ;
  assign n243 = ~n91 & n242 ;
  assign n244 = n243 ^ n203 ;
  assign n245 = n244 ^ n91 ;
  assign n246 = ~n240 & n245 ;
  assign n247 = n246 ^ n243 ;
  assign n248 = n247 ^ n91 ;
  assign n249 = ~x0 & ~n248 ;
  assign n250 = n249 ^ x0 ;
  assign n251 = n250 ^ n89 ;
  assign n252 = n251 ^ n250 ;
  assign n253 = ~x1 & x9 ;
  assign n254 = n253 ^ n250 ;
  assign n255 = n254 ^ n250 ;
  assign n256 = n252 & n255 ;
  assign n257 = n256 ^ n250 ;
  assign n258 = x3 & ~n257 ;
  assign n259 = n258 ^ n250 ;
  assign n260 = n237 & ~n259 ;
  assign n261 = n91 ^ n89 ;
  assign n262 = x9 & n261 ;
  assign n263 = n262 ^ n89 ;
  assign n264 = n168 & n263 ;
  assign n265 = n170 & n191 ;
  assign n266 = ~n264 & ~n265 ;
  assign n267 = x4 & n208 ;
  assign n268 = ~n266 & n267 ;
  assign n269 = x1 & x2 ;
  assign n270 = n81 & n269 ;
  assign n271 = x9 ^ x7 ;
  assign n272 = x9 ^ x5 ;
  assign n273 = n272 ^ x5 ;
  assign n274 = x5 ^ x0 ;
  assign n275 = ~n273 & ~n274 ;
  assign n276 = n275 ^ x5 ;
  assign n277 = n271 & n276 ;
  assign n278 = n270 & n277 ;
  assign n279 = ~x6 & ~n278 ;
  assign n280 = ~n268 & n279 ;
  assign n281 = x4 ^ x2 ;
  assign n57 = x5 & ~x9 ;
  assign n282 = n57 ^ x4 ;
  assign n283 = n282 ^ n57 ;
  assign n284 = n191 ^ n57 ;
  assign n285 = n283 & n284 ;
  assign n286 = n285 ^ n57 ;
  assign n287 = n281 & n286 ;
  assign n288 = n175 & n287 ;
  assign n289 = n81 & n152 ;
  assign n290 = n263 & n289 ;
  assign n291 = ~n288 & ~n290 ;
  assign n292 = n142 & ~n291 ;
  assign n28 = ~x2 & ~x9 ;
  assign n293 = ~n91 & ~n167 ;
  assign n294 = n28 & ~n293 ;
  assign n295 = ~x7 & n284 ;
  assign n296 = n295 ^ n57 ;
  assign n297 = n269 & n296 ;
  assign n298 = ~n294 & ~n297 ;
  assign n299 = x0 & n15 ;
  assign n300 = ~n298 & n299 ;
  assign n301 = ~n292 & ~n300 ;
  assign n302 = n280 & n301 ;
  assign n303 = ~n260 & n302 ;
  assign n304 = ~n236 & ~n303 ;
  assign n305 = ~n19 & ~n38 ;
  assign n306 = n165 & ~n305 ;
  assign n307 = n142 & n306 ;
  assign n308 = ~n11 & n307 ;
  assign n309 = ~n304 & ~n308 ;
  assign n20 = x6 & x9 ;
  assign n21 = n19 & n20 ;
  assign n22 = ~x5 & ~x6 ;
  assign n23 = x9 & n22 ;
  assign n24 = ~n21 & ~n23 ;
  assign n25 = ~x7 & ~n24 ;
  assign n26 = ~x2 & n25 ;
  assign n27 = ~x4 & x9 ;
  assign n29 = ~x6 & ~x9 ;
  assign n30 = ~n28 & n29 ;
  assign n31 = ~n27 & ~n30 ;
  assign n34 = n33 ^ n31 ;
  assign n43 = n34 ^ n31 ;
  assign n32 = n31 ^ n22 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = n36 ^ n31 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n39 ^ n35 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = ~n37 & ~n41 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = n44 ^ n37 ;
  assign n46 = n31 ^ n29 ;
  assign n47 = n42 ^ n37 ;
  assign n48 = n46 & ~n47 ;
  assign n49 = n48 ^ n31 ;
  assign n50 = ~n45 & n49 ;
  assign n51 = n50 ^ n31 ;
  assign n52 = n51 ^ n33 ;
  assign n53 = n52 ^ n31 ;
  assign n54 = ~n26 & ~n53 ;
  assign n55 = x0 & ~n54 ;
  assign n56 = ~x2 & x6 ;
  assign n58 = x7 & n57 ;
  assign n59 = n56 & n58 ;
  assign n62 = n59 ^ n13 ;
  assign n63 = n62 ^ n59 ;
  assign n60 = n59 ^ x5 ;
  assign n61 = n60 ^ n59 ;
  assign n64 = n63 ^ n61 ;
  assign n65 = n59 ^ x2 ;
  assign n66 = n65 ^ n59 ;
  assign n67 = n66 ^ n63 ;
  assign n68 = n63 & n67 ;
  assign n69 = n68 ^ n63 ;
  assign n70 = ~n64 & n69 ;
  assign n71 = n70 ^ n68 ;
  assign n72 = n71 ^ n59 ;
  assign n73 = n72 ^ n63 ;
  assign n74 = ~x4 & n73 ;
  assign n75 = n74 ^ n59 ;
  assign n76 = ~n55 & ~n75 ;
  assign n77 = x3 & ~n76 ;
  assign n78 = n77 ^ x0 ;
  assign n79 = n78 ^ n77 ;
  assign n83 = n13 & ~n82 ;
  assign n84 = x3 & x4 ;
  assign n85 = ~x2 & ~n84 ;
  assign n86 = n83 & n85 ;
  assign n87 = n86 ^ x6 ;
  assign n88 = x9 ^ x4 ;
  assign n93 = ~n90 & ~n92 ;
  assign n94 = n93 ^ x9 ;
  assign n95 = n94 ^ n93 ;
  assign n96 = n95 ^ n88 ;
  assign n97 = n33 ^ x3 ;
  assign n98 = ~x3 & n97 ;
  assign n99 = n98 ^ n93 ;
  assign n100 = n99 ^ x3 ;
  assign n101 = n96 & n100 ;
  assign n102 = n101 ^ n98 ;
  assign n103 = n102 ^ x3 ;
  assign n104 = ~n88 & ~n103 ;
  assign n105 = n104 ^ x2 ;
  assign n106 = n105 ^ n104 ;
  assign n113 = x4 & n89 ;
  assign n114 = ~x9 & n113 ;
  assign n109 = n107 & n108 ;
  assign n110 = x4 & x9 ;
  assign n111 = ~x5 & n110 ;
  assign n112 = ~n109 & ~n111 ;
  assign n115 = n114 ^ n112 ;
  assign n116 = n115 ^ n112 ;
  assign n117 = x5 & x7 ;
  assign n118 = n27 & n117 ;
  assign n119 = n118 ^ n112 ;
  assign n120 = n119 ^ n112 ;
  assign n121 = ~n116 & ~n120 ;
  assign n122 = n121 ^ n112 ;
  assign n123 = ~x3 & n122 ;
  assign n124 = n123 ^ n112 ;
  assign n125 = n124 ^ n104 ;
  assign n126 = ~n106 & ~n125 ;
  assign n127 = n126 ^ n104 ;
  assign n128 = n127 ^ n86 ;
  assign n129 = ~n87 & ~n128 ;
  assign n130 = n129 ^ n126 ;
  assign n131 = n130 ^ n104 ;
  assign n132 = n131 ^ x6 ;
  assign n133 = ~n86 & n132 ;
  assign n134 = n133 ^ n86 ;
  assign n135 = n134 ^ n86 ;
  assign n136 = n135 ^ n77 ;
  assign n137 = n136 ^ n77 ;
  assign n138 = n79 & ~n137 ;
  assign n139 = n138 ^ n77 ;
  assign n140 = x1 & n139 ;
  assign n141 = n140 ^ n77 ;
  assign n310 = n309 ^ n141 ;
  assign n311 = n310 ^ n309 ;
  assign n312 = n15 & n203 ;
  assign n313 = n84 & n107 ;
  assign n314 = ~n90 & ~n313 ;
  assign n315 = ~n19 & ~n314 ;
  assign n316 = ~n312 & ~n315 ;
  assign n317 = x6 & ~n316 ;
  assign n318 = ~x3 & ~x6 ;
  assign n319 = n89 & n318 ;
  assign n320 = ~x9 & n319 ;
  assign n321 = x2 & ~n320 ;
  assign n322 = ~n317 & n321 ;
  assign n323 = ~x0 & ~n322 ;
  assign n325 = ~x4 & n29 ;
  assign n326 = ~n21 & ~n325 ;
  assign n327 = x7 & n202 ;
  assign n328 = ~n326 & n327 ;
  assign n329 = n88 ^ x4 ;
  assign n330 = x4 ^ x1 ;
  assign n331 = n329 & ~n330 ;
  assign n332 = n331 ^ x4 ;
  assign n333 = n319 & n332 ;
  assign n334 = ~n328 & ~n333 ;
  assign n324 = x2 ^ x1 ;
  assign n335 = n334 ^ n324 ;
  assign n337 = n165 ^ x4 ;
  assign n338 = n337 ^ n165 ;
  assign n339 = n338 ^ x1 ;
  assign n340 = n12 ^ x3 ;
  assign n341 = n12 & n340 ;
  assign n342 = n341 ^ n165 ;
  assign n343 = n342 ^ n12 ;
  assign n344 = n339 & n343 ;
  assign n345 = n344 ^ n341 ;
  assign n346 = n345 ^ n12 ;
  assign n347 = x1 & n346 ;
  assign n348 = n347 ^ x1 ;
  assign n349 = ~n11 & ~n348 ;
  assign n350 = n349 ^ n334 ;
  assign n336 = n335 ^ x2 ;
  assign n351 = n350 ^ n336 ;
  assign n352 = n349 ^ n336 ;
  assign n353 = n352 ^ n335 ;
  assign n354 = n351 & n353 ;
  assign n355 = n354 ^ n349 ;
  assign n356 = ~x4 & ~x6 ;
  assign n357 = n107 ^ x3 ;
  assign n358 = n356 & ~n357 ;
  assign n359 = n349 & n358 ;
  assign n360 = n359 ^ n335 ;
  assign n361 = n355 & n360 ;
  assign n362 = n361 ^ n359 ;
  assign n363 = n335 & n362 ;
  assign n364 = n363 ^ n354 ;
  assign n365 = n364 ^ n334 ;
  assign n366 = n365 ^ n349 ;
  assign n367 = n323 & ~n366 ;
  assign n368 = n367 ^ n309 ;
  assign n369 = n368 ^ n309 ;
  assign n370 = ~n311 & ~n369 ;
  assign n371 = n370 ^ n309 ;
  assign n372 = x8 & n371 ;
  assign n373 = n372 ^ n309 ;
  assign n374 = ~n18 & n373 ;
  assign y0 = ~n374 ;
endmodule
