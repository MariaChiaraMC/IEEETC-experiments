module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 ;
  assign n9 = x2 ^ x1 ;
  assign n10 = n9 ^ x1 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = n12 ^ x0 ;
  assign n14 = ~n11 & n13 ;
  assign n15 = n14 ^ n10 ;
  assign n16 = n15 ^ n11 ;
  assign n23 = x5 ^ x4 ;
  assign n24 = n23 ^ x6 ;
  assign n21 = x4 ^ x2 ;
  assign n22 = n21 ^ x6 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = x6 ^ x4 ;
  assign n28 = n27 ^ n22 ;
  assign n29 = n28 ^ n22 ;
  assign n30 = n29 ^ x4 ;
  assign n31 = n30 ^ x7 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = ~n22 & ~n32 ;
  assign n34 = n33 ^ x4 ;
  assign n35 = n34 ^ n26 ;
  assign n36 = n30 ^ n22 ;
  assign n37 = n36 ^ n26 ;
  assign n38 = x4 & n37 ;
  assign n39 = n38 ^ n22 ;
  assign n40 = ~n35 & ~n39 ;
  assign n41 = ~n26 & n40 ;
  assign n42 = n41 ^ n33 ;
  assign n43 = n42 ^ n38 ;
  assign n44 = n43 ^ n40 ;
  assign n45 = n44 ^ n11 ;
  assign n46 = ~n11 & n45 ;
  assign n17 = x4 & ~x5 ;
  assign n18 = n10 ^ x3 ;
  assign n19 = n18 ^ n11 ;
  assign n20 = ~n17 & ~n19 ;
  assign n47 = n46 ^ n20 ;
  assign n48 = n47 ^ n10 ;
  assign n49 = n48 ^ x3 ;
  assign n50 = n49 ^ n11 ;
  assign n51 = n50 ^ x0 ;
  assign n52 = ~x3 & ~n51 ;
  assign n53 = n52 ^ n20 ;
  assign n54 = n53 ^ n10 ;
  assign n55 = n54 ^ n11 ;
  assign n56 = n55 ^ x0 ;
  assign n57 = n16 & n56 ;
  assign n58 = n57 ^ n20 ;
  assign n59 = n58 ^ n14 ;
  assign n60 = n59 ^ n52 ;
  assign n61 = n60 ^ x0 ;
  assign n62 = n61 ^ x0 ;
  assign y0 = n62 ;
endmodule
