module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 ;
  assign n16 = x2 & x3 ;
  assign n17 = ~x9 & ~n16 ;
  assign n18 = ~x2 & ~x3 ;
  assign n19 = x10 & x12 ;
  assign n20 = x14 & n19 ;
  assign n21 = ~n18 & n20 ;
  assign n22 = n17 & n21 ;
  assign n23 = x11 & n22 ;
  assign n24 = ~x4 & ~x6 ;
  assign n25 = n18 & n24 ;
  assign n26 = ~x1 & n25 ;
  assign n27 = x9 & ~n26 ;
  assign n28 = ~x10 & ~x11 ;
  assign n29 = ~x12 & n28 ;
  assign n31 = ~x1 & ~x9 ;
  assign n32 = ~x4 & x7 ;
  assign n33 = x6 & n32 ;
  assign n34 = ~n31 & ~n33 ;
  assign n30 = ~x1 & ~x3 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n34 ^ x5 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = n37 ^ n29 ;
  assign n39 = n38 ^ n28 ;
  assign n40 = ~n35 & ~n39 ;
  assign n41 = n40 ^ n34 ;
  assign n42 = n29 & ~n41 ;
  assign n43 = n42 ^ n29 ;
  assign n44 = n43 ^ n27 ;
  assign n45 = ~x7 & n24 ;
  assign n46 = x1 & ~n45 ;
  assign n47 = ~x5 & ~n46 ;
  assign n48 = ~n17 & ~n47 ;
  assign n49 = n48 ^ x0 ;
  assign n50 = n49 ^ n48 ;
  assign n53 = ~x3 & ~x5 ;
  assign n51 = x5 & ~x7 ;
  assign n52 = ~x6 & ~n51 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = ~x2 & ~n54 ;
  assign n56 = n54 ^ n52 ;
  assign n57 = ~x1 & ~x7 ;
  assign n58 = x3 & ~n57 ;
  assign n59 = x4 & ~n58 ;
  assign n60 = n59 ^ n55 ;
  assign n61 = n56 & n60 ;
  assign n62 = n61 ^ n59 ;
  assign n63 = n55 & n62 ;
  assign n64 = n63 ^ n53 ;
  assign n65 = n64 ^ n48 ;
  assign n66 = n50 & n65 ;
  assign n67 = n66 ^ n48 ;
  assign n68 = n67 ^ n27 ;
  assign n69 = ~n44 & ~n68 ;
  assign n70 = n69 ^ n66 ;
  assign n71 = n70 ^ n48 ;
  assign n72 = n71 ^ n43 ;
  assign n73 = ~n27 & n72 ;
  assign n74 = n73 ^ n27 ;
  assign n75 = ~n23 & n74 ;
  assign n76 = ~x13 & ~n75 ;
  assign y0 = n76 ;
endmodule
