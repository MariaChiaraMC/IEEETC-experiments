module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 ;
  assign n15 = ~x2 & ~x8 ;
  assign n16 = x12 & ~x13 ;
  assign n17 = ~x11 & n16 ;
  assign n18 = ~x10 & n17 ;
  assign n19 = n15 & n18 ;
  assign n20 = x2 & ~x3 ;
  assign n21 = x0 & x13 ;
  assign n22 = n20 & ~n21 ;
  assign n23 = ~x12 & n22 ;
  assign n24 = ~x4 & x5 ;
  assign n25 = ~x6 & ~x7 ;
  assign n26 = ~x10 & ~n25 ;
  assign n27 = n24 & n26 ;
  assign n28 = n23 & n27 ;
  assign n29 = x2 & ~x12 ;
  assign n32 = x12 ^ x4 ;
  assign n30 = x12 ^ x7 ;
  assign n31 = n30 ^ x12 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = x12 ^ x5 ;
  assign n35 = n34 ^ x12 ;
  assign n36 = n35 ^ n31 ;
  assign n37 = n31 & ~n36 ;
  assign n38 = n37 ^ n31 ;
  assign n39 = n33 & n38 ;
  assign n40 = n39 ^ n37 ;
  assign n41 = n40 ^ x12 ;
  assign n42 = n41 ^ n31 ;
  assign n43 = ~x6 & ~n42 ;
  assign n44 = n43 ^ n37 ;
  assign n45 = n44 ^ n31 ;
  assign n46 = n45 ^ x12 ;
  assign n47 = n46 ^ x12 ;
  assign n48 = ~n29 & ~n47 ;
  assign n49 = x10 & x13 ;
  assign n50 = ~n48 & n49 ;
  assign n51 = ~x6 & x7 ;
  assign n52 = x5 & n51 ;
  assign n53 = x12 & ~n52 ;
  assign n54 = x11 & ~n53 ;
  assign n55 = ~n50 & n54 ;
  assign n56 = ~n28 & ~n55 ;
  assign n57 = x12 ^ x0 ;
  assign n58 = x12 ^ x10 ;
  assign n59 = n58 ^ n57 ;
  assign n60 = n57 & n59 ;
  assign n61 = n60 ^ x12 ;
  assign n62 = n61 ^ n57 ;
  assign n63 = x11 ^ x0 ;
  assign n69 = n63 ^ x13 ;
  assign n64 = n63 ^ x0 ;
  assign n65 = n64 ^ x12 ;
  assign n66 = n65 ^ n57 ;
  assign n67 = ~x12 & n66 ;
  assign n68 = n67 ^ n64 ;
  assign n70 = n69 ^ n68 ;
  assign n71 = n64 ^ x1 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = ~x1 & ~n72 ;
  assign n74 = n73 ^ x12 ;
  assign n75 = n70 & ~n74 ;
  assign n76 = n75 ^ n64 ;
  assign n77 = n76 ^ n57 ;
  assign n78 = n77 ^ n58 ;
  assign n79 = ~n62 & ~n78 ;
  assign n80 = n79 ^ n67 ;
  assign n81 = n80 ^ n75 ;
  assign n82 = n81 ^ x12 ;
  assign n83 = n82 ^ x10 ;
  assign n84 = n56 & n83 ;
  assign n85 = x8 & ~n84 ;
  assign n86 = x11 & x13 ;
  assign n87 = ~x6 & x8 ;
  assign n88 = ~n86 & ~n87 ;
  assign n89 = ~n29 & ~n88 ;
  assign n90 = x4 & n49 ;
  assign n91 = ~x12 & n90 ;
  assign n92 = ~x8 & n91 ;
  assign n93 = ~x3 & ~x12 ;
  assign n94 = ~x10 & x13 ;
  assign n95 = ~n93 & n94 ;
  assign n96 = n15 & ~n95 ;
  assign n97 = ~n92 & ~n96 ;
  assign n98 = n97 ^ x11 ;
  assign n99 = n98 ^ n97 ;
  assign n100 = n97 ^ x10 ;
  assign n101 = n99 & n100 ;
  assign n102 = n101 ^ n97 ;
  assign n103 = ~n89 & ~n102 ;
  assign n104 = ~n85 & ~n103 ;
  assign n105 = n104 ^ x9 ;
  assign n106 = n105 ^ n104 ;
  assign n107 = x10 & x11 ;
  assign n108 = n93 & n107 ;
  assign n109 = x3 & x6 ;
  assign n110 = x1 & n109 ;
  assign n111 = ~x4 & n110 ;
  assign n112 = n18 & ~n111 ;
  assign n113 = ~n108 & ~n112 ;
  assign n114 = ~x8 & ~n113 ;
  assign n115 = x8 & n20 ;
  assign n116 = ~n107 & ~n115 ;
  assign n117 = ~x12 & n51 ;
  assign n118 = ~x11 & ~n117 ;
  assign n119 = ~n116 & ~n118 ;
  assign n128 = ~x5 & n51 ;
  assign n120 = ~x0 & ~x11 ;
  assign n121 = ~x0 & x1 ;
  assign n122 = n15 & n121 ;
  assign n123 = n109 & n122 ;
  assign n124 = n16 & n123 ;
  assign n125 = ~n120 & ~n124 ;
  assign n129 = n128 ^ n125 ;
  assign n130 = n129 ^ n125 ;
  assign n126 = n125 ^ x13 ;
  assign n127 = n126 ^ n125 ;
  assign n131 = n130 ^ n127 ;
  assign n132 = n125 ^ x12 ;
  assign n133 = n132 ^ n125 ;
  assign n134 = n133 ^ n130 ;
  assign n135 = n130 & n134 ;
  assign n136 = n135 ^ n130 ;
  assign n137 = n131 & n136 ;
  assign n138 = n137 ^ n135 ;
  assign n139 = n138 ^ n125 ;
  assign n140 = n139 ^ n130 ;
  assign n141 = ~x10 & ~n140 ;
  assign n142 = n141 ^ n125 ;
  assign n143 = n119 & ~n142 ;
  assign n144 = ~x4 & n143 ;
  assign n145 = ~n114 & ~n144 ;
  assign n146 = n145 ^ n104 ;
  assign n147 = n106 & n146 ;
  assign n148 = n147 ^ n104 ;
  assign n149 = ~n19 & n148 ;
  assign y0 = ~n149 ;
endmodule
