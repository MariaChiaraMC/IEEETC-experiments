module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 ;
  assign n17 = ~x14 & ~x15 ;
  assign n18 = ~x12 & ~x13 ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = x5 & ~x7 ;
  assign n21 = n20 ^ x4 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = ~x8 & ~x9 ;
  assign n24 = x11 ^ x10 ;
  assign n25 = n23 & n24 ;
  assign n26 = x7 & ~n25 ;
  assign n27 = ~x10 & ~x11 ;
  assign n28 = x9 ^ x8 ;
  assign n29 = n27 & n28 ;
  assign n30 = n26 & ~n29 ;
  assign n31 = n30 ^ n21 ;
  assign n32 = n31 ^ n22 ;
  assign n33 = ~n22 & n32 ;
  assign n34 = n33 ^ n21 ;
  assign n35 = n34 ^ n22 ;
  assign n36 = n20 ^ x5 ;
  assign n37 = x6 & ~n36 ;
  assign n38 = n37 ^ n21 ;
  assign n39 = ~n35 & n38 ;
  assign n40 = n39 ^ n21 ;
  assign n41 = n40 ^ n21 ;
  assign n42 = ~n19 & n41 ;
  assign n43 = ~x10 & x11 ;
  assign n44 = ~x13 & ~x15 ;
  assign n45 = ~n43 & ~n44 ;
  assign n46 = x14 ^ x12 ;
  assign n48 = x14 ^ x13 ;
  assign n47 = x15 ^ x14 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = n49 ^ n46 ;
  assign n51 = x10 & ~x11 ;
  assign n52 = n51 ^ x15 ;
  assign n53 = ~x15 & ~n52 ;
  assign n54 = n53 ^ n48 ;
  assign n55 = n54 ^ x15 ;
  assign n56 = ~n50 & ~n55 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n57 ^ x15 ;
  assign n59 = n46 & ~n58 ;
  assign n60 = x5 & x6 ;
  assign n61 = x4 & n60 ;
  assign n62 = n28 & n61 ;
  assign n63 = n59 & n62 ;
  assign n64 = ~n45 & n63 ;
  assign n65 = ~n42 & ~n64 ;
  assign n66 = ~x1 & ~x2 ;
  assign n67 = ~x0 & n66 ;
  assign n68 = ~x3 & n67 ;
  assign n69 = ~n65 & n68 ;
  assign y0 = n69 ;
endmodule
