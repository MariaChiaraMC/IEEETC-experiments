module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 ;
  assign n94 = x19 ^ x18 ;
  assign n95 = ~x19 & x20 ;
  assign n96 = n94 & n95 ;
  assign n97 = n96 ^ n94 ;
  assign n98 = ~x17 & n97 ;
  assign n22 = ~x5 & x9 ;
  assign n27 = x12 & x13 ;
  assign n28 = x14 & n27 ;
  assign n29 = ~x16 & ~n28 ;
  assign n23 = ~x12 & ~x13 ;
  assign n24 = x14 & ~n23 ;
  assign n25 = x4 & ~n24 ;
  assign n26 = x2 & n25 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n30 ^ n26 ;
  assign n32 = ~x2 & x4 ;
  assign n33 = x10 & n32 ;
  assign n34 = n33 ^ n26 ;
  assign n35 = n34 ^ n26 ;
  assign n36 = n31 & n35 ;
  assign n37 = n36 ^ n26 ;
  assign n38 = x1 & n37 ;
  assign n39 = n38 ^ n26 ;
  assign n40 = n22 & n39 ;
  assign n41 = n40 ^ x0 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = n40 ^ x2 ;
  assign n44 = n43 ^ n41 ;
  assign n45 = n44 ^ x1 ;
  assign n63 = n45 ^ n41 ;
  assign n64 = n63 ^ n40 ;
  assign n46 = x3 & x7 ;
  assign n47 = x3 & x4 ;
  assign n48 = n29 & n47 ;
  assign n49 = ~x5 & n48 ;
  assign n50 = ~n46 & ~n49 ;
  assign n51 = ~x8 & ~n50 ;
  assign n52 = ~x5 & n25 ;
  assign n53 = ~x8 & ~n52 ;
  assign n54 = ~x6 & n53 ;
  assign n55 = x0 & ~n54 ;
  assign n56 = ~x3 & n55 ;
  assign n57 = ~n51 & ~n56 ;
  assign n58 = n57 ^ n45 ;
  assign n59 = n58 ^ x1 ;
  assign n60 = n59 ^ n58 ;
  assign n61 = n60 ^ n40 ;
  assign n62 = n61 ^ n42 ;
  assign n65 = n64 ^ n62 ;
  assign n66 = ~n42 & n65 ;
  assign n67 = n66 ^ n60 ;
  assign n68 = n67 ^ n64 ;
  assign n84 = n58 ^ n45 ;
  assign n69 = ~n27 & n47 ;
  assign n70 = x13 & x15 ;
  assign n71 = x7 ^ x6 ;
  assign n72 = x3 & n71 ;
  assign n73 = n72 ^ x6 ;
  assign n74 = ~n70 & n73 ;
  assign n75 = ~n25 & ~n74 ;
  assign n76 = ~n69 & n75 ;
  assign n77 = ~x15 & x16 ;
  assign n78 = x5 & ~n77 ;
  assign n79 = ~n76 & n78 ;
  assign n80 = n79 ^ n58 ;
  assign n81 = n64 ^ n60 ;
  assign n82 = ~n80 & ~n81 ;
  assign n83 = n82 ^ n66 ;
  assign n85 = n84 ^ n83 ;
  assign n86 = n85 ^ n80 ;
  assign n87 = n86 ^ n60 ;
  assign n88 = ~n64 & n87 ;
  assign n89 = n88 ^ n42 ;
  assign n90 = ~n68 & ~n89 ;
  assign n91 = n90 ^ n42 ;
  assign n92 = n91 ^ x0 ;
  assign n93 = n92 ^ n42 ;
  assign n99 = n98 ^ n93 ;
  assign n100 = ~x11 & ~n99 ;
  assign n101 = n100 ^ n93 ;
  assign y0 = ~n101 ;
endmodule
