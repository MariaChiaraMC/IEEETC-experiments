module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 ;
  assign n9 = x3 ^ x2 ;
  assign n7 = x3 ^ x1 ;
  assign n16 = n9 ^ n7 ;
  assign n8 = n7 ^ x3 ;
  assign n10 = n9 ^ n8 ;
  assign n11 = n10 ^ n7 ;
  assign n12 = n8 ^ x4 ;
  assign n13 = n12 ^ n8 ;
  assign n14 = n13 ^ n11 ;
  assign n15 = n11 & n14 ;
  assign n17 = n16 ^ n15 ;
  assign n18 = n17 ^ n11 ;
  assign n19 = n7 ^ x5 ;
  assign n20 = n15 ^ n11 ;
  assign n21 = ~n19 & n20 ;
  assign n22 = n21 ^ n7 ;
  assign n23 = n18 & n22 ;
  assign n24 = n23 ^ n7 ;
  assign n25 = n24 ^ x1 ;
  assign n26 = n25 ^ n7 ;
  assign n27 = ~x0 & n26 ;
  assign y0 = n27 ;
endmodule
