module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n9 = ~x1 & ~x3 ;
  assign n10 = ~x0 & n9 ;
  assign n11 = x6 ^ x4 ;
  assign n12 = n11 ^ x7 ;
  assign n13 = x5 ^ x2 ;
  assign n14 = n13 ^ x6 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = x7 ^ x5 ;
  assign n17 = n16 ^ x7 ;
  assign n18 = x7 ^ x6 ;
  assign n19 = n18 ^ x7 ;
  assign n20 = ~n17 & n19 ;
  assign n21 = n20 ^ x7 ;
  assign n22 = n21 ^ n12 ;
  assign n23 = ~n15 & n22 ;
  assign n24 = n23 ^ n20 ;
  assign n25 = n24 ^ x7 ;
  assign n26 = n25 ^ n14 ;
  assign n27 = ~n12 & ~n26 ;
  assign n28 = n27 ^ n12 ;
  assign n29 = n10 & ~n28 ;
  assign y0 = n29 ;
endmodule
