module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 ;
  assign n17 = x14 & ~x15 ;
  assign n18 = ~x14 & x15 ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = x12 & ~x13 ;
  assign n21 = ~x12 & x13 ;
  assign n22 = ~n20 & ~n21 ;
  assign n23 = n19 & n22 ;
  assign n43 = ~x4 & ~x5 ;
  assign n24 = x5 & ~x10 ;
  assign n25 = x8 & ~x9 ;
  assign n26 = n24 & n25 ;
  assign n27 = ~x11 & n26 ;
  assign n28 = x6 ^ x4 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = x10 & ~x11 ;
  assign n31 = x11 & n24 ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = ~x8 & ~x9 ;
  assign n34 = ~n32 & n33 ;
  assign n35 = n34 ^ x5 ;
  assign n36 = x6 & ~n35 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = n29 & ~n37 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n39 ^ n34 ;
  assign n41 = n40 ^ x6 ;
  assign n42 = ~n27 & ~n41 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = n44 ^ x7 ;
  assign n56 = n45 ^ n44 ;
  assign n46 = x7 & ~x10 ;
  assign n47 = ~x8 & ~x11 ;
  assign n48 = n46 & n47 ;
  assign n49 = x9 & n48 ;
  assign n50 = n49 ^ n45 ;
  assign n51 = n50 ^ n44 ;
  assign n52 = n45 ^ n42 ;
  assign n53 = n52 ^ n49 ;
  assign n54 = n53 ^ n51 ;
  assign n55 = ~n51 & n54 ;
  assign n57 = n56 ^ n55 ;
  assign n58 = n57 ^ n51 ;
  assign n59 = x4 & x5 ;
  assign n60 = n59 ^ n44 ;
  assign n61 = n55 ^ n51 ;
  assign n62 = n60 & ~n61 ;
  assign n63 = n62 ^ n44 ;
  assign n64 = ~n58 & n63 ;
  assign n65 = n64 ^ n44 ;
  assign n66 = n65 ^ n43 ;
  assign n67 = n66 ^ n44 ;
  assign n68 = ~n23 & ~n67 ;
  assign n94 = x7 & n43 ;
  assign n95 = n30 & n94 ;
  assign n71 = x13 ^ x12 ;
  assign n72 = n71 ^ x14 ;
  assign n73 = n72 ^ x15 ;
  assign n74 = x15 ^ x13 ;
  assign n75 = x14 ^ x13 ;
  assign n76 = n74 & n75 ;
  assign n77 = n76 ^ x13 ;
  assign n78 = n73 & n77 ;
  assign n79 = n31 & n78 ;
  assign n69 = n43 ^ x7 ;
  assign n70 = n69 ^ n43 ;
  assign n80 = n79 ^ n70 ;
  assign n81 = n80 ^ n79 ;
  assign n82 = n81 ^ n69 ;
  assign n83 = n82 ^ n81 ;
  assign n84 = n25 & ~n83 ;
  assign n85 = n84 ^ n79 ;
  assign n86 = n79 ^ n30 ;
  assign n87 = n82 & ~n86 ;
  assign n88 = n87 ^ n81 ;
  assign n89 = n88 ^ n82 ;
  assign n90 = ~n85 & ~n89 ;
  assign n91 = ~n81 & n90 ;
  assign n92 = n91 ^ n84 ;
  assign n93 = n92 ^ x7 ;
  assign n96 = n95 ^ n93 ;
  assign n97 = n96 ^ n95 ;
  assign n98 = x10 ^ x7 ;
  assign n99 = ~n17 & ~n20 ;
  assign n100 = n99 ^ x10 ;
  assign n101 = n100 ^ n99 ;
  assign n102 = n101 ^ n98 ;
  assign n103 = ~x5 & ~n25 ;
  assign n104 = n103 ^ n23 ;
  assign n105 = ~n103 & n104 ;
  assign n106 = n105 ^ n99 ;
  assign n107 = n106 ^ n103 ;
  assign n108 = ~n102 & n107 ;
  assign n109 = n108 ^ n105 ;
  assign n110 = n109 ^ n103 ;
  assign n111 = n98 & ~n110 ;
  assign n112 = ~x11 & n111 ;
  assign n113 = n112 ^ n95 ;
  assign n114 = n113 ^ n95 ;
  assign n115 = n97 & ~n114 ;
  assign n116 = n115 ^ n95 ;
  assign n117 = x6 & ~n116 ;
  assign n118 = n117 ^ n95 ;
  assign n119 = ~n68 & ~n118 ;
  assign y0 = ~n119 ;
endmodule
