module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 ;
  assign n16 = ~x1 & ~x3 ;
  assign n17 = ~x0 & n16 ;
  assign n18 = x12 & x13 ;
  assign n19 = ~x2 & ~n18 ;
  assign n20 = ~x5 & ~x6 ;
  assign n21 = ~x8 & n20 ;
  assign n22 = n19 & n21 ;
  assign n23 = n17 & n22 ;
  assign n24 = ~x7 & ~x9 ;
  assign n25 = ~x4 & ~x10 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = ~x12 & ~x13 ;
  assign n28 = ~x14 & n27 ;
  assign n29 = n28 ^ x11 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = n28 ^ n27 ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = n32 ^ n28 ;
  assign n34 = n33 ^ n24 ;
  assign n35 = n26 & n34 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ n28 ;
  assign n38 = n37 ^ n25 ;
  assign n39 = n24 & n38 ;
  assign n40 = n39 ^ n24 ;
  assign n41 = n23 & n40 ;
  assign y0 = n41 ;
endmodule
