module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 ;
  assign n9 = x1 & x5 ;
  assign n10 = x3 & x7 ;
  assign n11 = ~x2 & ~n10 ;
  assign n12 = ~x6 & n11 ;
  assign n13 = ~n9 & n12 ;
  assign n15 = x2 & x3 ;
  assign n14 = ~x1 & ~x5 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = n14 ^ x0 ;
  assign n18 = x6 & x7 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n19 ^ n14 ;
  assign n21 = ~n14 & n20 ;
  assign n22 = n21 ^ n14 ;
  assign n23 = ~n17 & ~n22 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n24 ^ n14 ;
  assign n26 = n25 ^ n19 ;
  assign n27 = ~n16 & n26 ;
  assign n28 = n27 ^ n14 ;
  assign n29 = ~n13 & ~n28 ;
  assign n30 = x6 & n9 ;
  assign n31 = ~x0 & ~n30 ;
  assign n32 = x4 & ~n31 ;
  assign n33 = n29 & n32 ;
  assign n34 = x0 & n9 ;
  assign n35 = ~x3 & ~n18 ;
  assign n36 = n34 & ~n35 ;
  assign n37 = x2 & n36 ;
  assign n38 = ~n33 & ~n37 ;
  assign y0 = ~n38 ;
endmodule
