module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 ;
  assign n9 = ~x0 & ~x1 ;
  assign n10 = ~x2 & ~x3 ;
  assign n11 = n9 & n10 ;
  assign n12 = x5 ^ x4 ;
  assign n13 = n12 ^ x6 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = x5 & ~x7 ;
  assign n17 = n16 ^ x4 ;
  assign n18 = ~x4 & ~n17 ;
  assign n19 = n18 ^ n12 ;
  assign n20 = n19 ^ x4 ;
  assign n21 = ~n15 & n20 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = n22 ^ x4 ;
  assign n24 = n11 & ~n23 ;
  assign n25 = n24 ^ n11 ;
  assign y0 = n25 ;
endmodule
