module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 ;
  assign n16 = x7 & ~x9 ;
  assign n17 = x0 & ~x10 ;
  assign n18 = ~x4 & ~x5 ;
  assign n19 = n17 & n18 ;
  assign n20 = ~x13 & ~x14 ;
  assign n21 = ~x1 & x6 ;
  assign n22 = n20 & n21 ;
  assign n23 = n19 & n22 ;
  assign n24 = n16 & n23 ;
  assign n25 = ~x2 & ~x8 ;
  assign n26 = n24 & n25 ;
  assign n27 = ~x3 & ~n26 ;
  assign n28 = ~x11 & ~n27 ;
  assign n29 = ~x12 & n28 ;
  assign n30 = ~x0 & x9 ;
  assign n31 = x1 & n30 ;
  assign n32 = ~x5 & ~x13 ;
  assign n33 = x4 & ~x8 ;
  assign n34 = ~n32 & n33 ;
  assign n35 = n31 & n34 ;
  assign n36 = n35 ^ n20 ;
  assign n37 = x6 & ~x10 ;
  assign n38 = ~x5 & ~n37 ;
  assign n39 = n38 ^ x7 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = x6 & x10 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = ~n40 & ~n42 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = n44 ^ n35 ;
  assign n46 = ~n36 & n45 ;
  assign n47 = n46 ^ n43 ;
  assign n48 = n47 ^ n38 ;
  assign n49 = n48 ^ n20 ;
  assign n50 = n35 & ~n49 ;
  assign n51 = n50 ^ n35 ;
  assign n52 = ~n24 & ~n51 ;
  assign n53 = x2 & ~n52 ;
  assign n54 = x8 & n23 ;
  assign n55 = x9 ^ x7 ;
  assign n56 = n54 & n55 ;
  assign n57 = x3 & ~n56 ;
  assign n58 = ~n53 & n57 ;
  assign n59 = n29 & ~n58 ;
  assign y0 = n59 ;
endmodule
