module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 ;
  assign n17 = ~x2 & ~x3 ;
  assign n18 = ~x0 & n17 ;
  assign n19 = ~x1 & n18 ;
  assign n20 = ~x4 & ~x5 ;
  assign n21 = x4 & x5 ;
  assign n22 = ~n20 & ~n21 ;
  assign n23 = ~x7 & ~n22 ;
  assign n24 = ~x14 & ~x15 ;
  assign n25 = ~x12 & ~x13 ;
  assign n26 = ~n24 & ~n25 ;
  assign n27 = x8 ^ x5 ;
  assign n28 = n27 ^ x9 ;
  assign n29 = x8 ^ x6 ;
  assign n30 = n29 ^ x9 ;
  assign n32 = n30 ^ x8 ;
  assign n33 = n32 ^ n30 ;
  assign n31 = n30 ^ x4 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n30 ^ x9 ;
  assign n36 = n35 ^ n30 ;
  assign n37 = n36 ^ n33 ;
  assign n38 = n33 & ~n37 ;
  assign n39 = n38 ^ n33 ;
  assign n40 = ~n34 & n39 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n41 ^ n30 ;
  assign n43 = n42 ^ n33 ;
  assign n44 = n28 & ~n43 ;
  assign n45 = n44 ^ x5 ;
  assign n46 = ~x10 & n45 ;
  assign n47 = ~x11 & n46 ;
  assign n48 = x6 ^ x4 ;
  assign n49 = n48 ^ x7 ;
  assign n50 = x5 & ~x8 ;
  assign n51 = ~x9 & n50 ;
  assign n52 = x11 ^ x10 ;
  assign n53 = n51 & n52 ;
  assign n54 = n53 ^ x5 ;
  assign n55 = x6 & ~n54 ;
  assign n56 = n55 ^ n53 ;
  assign n57 = ~n49 & ~n56 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = n58 ^ n53 ;
  assign n60 = n59 ^ x6 ;
  assign n61 = x7 & ~n60 ;
  assign n62 = ~n47 & n61 ;
  assign n63 = ~n26 & ~n62 ;
  assign n64 = ~n23 & n63 ;
  assign n65 = x6 & ~x8 ;
  assign n66 = n20 & n65 ;
  assign n67 = x9 & n66 ;
  assign n68 = n67 ^ x7 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = n69 ^ n64 ;
  assign n71 = x14 ^ x12 ;
  assign n73 = x14 ^ x13 ;
  assign n72 = x15 ^ x14 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = n74 ^ n71 ;
  assign n76 = x10 & ~x11 ;
  assign n77 = n76 ^ x15 ;
  assign n78 = ~x15 & ~n77 ;
  assign n79 = n78 ^ n73 ;
  assign n80 = n79 ^ x15 ;
  assign n81 = ~n75 & ~n80 ;
  assign n82 = n81 ^ n78 ;
  assign n83 = n82 ^ x15 ;
  assign n84 = n71 & ~n83 ;
  assign n85 = ~x10 & x11 ;
  assign n86 = ~x13 & ~x15 ;
  assign n87 = ~n85 & ~n86 ;
  assign n88 = x5 & x6 ;
  assign n89 = ~n87 & n88 ;
  assign n90 = n89 ^ n84 ;
  assign n91 = n84 & n90 ;
  assign n92 = n91 ^ n67 ;
  assign n93 = n92 ^ n84 ;
  assign n94 = n70 & n93 ;
  assign n95 = n94 ^ n91 ;
  assign n96 = n95 ^ n84 ;
  assign n97 = ~n64 & n96 ;
  assign n98 = n97 ^ n64 ;
  assign n99 = n19 & n98 ;
  assign y0 = n99 ;
endmodule
