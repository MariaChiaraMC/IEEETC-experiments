module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n13 = x4 & ~x8 ;
  assign n14 = ~x7 & n13 ;
  assign n15 = x2 & x3 ;
  assign n16 = x9 & ~n15 ;
  assign n17 = n14 & n16 ;
  assign n18 = ~x3 & ~x10 ;
  assign n19 = ~x2 & ~n18 ;
  assign n20 = x7 & ~n19 ;
  assign n21 = x8 ^ x4 ;
  assign n22 = x9 ^ x3 ;
  assign n23 = x8 ^ x3 ;
  assign n24 = n23 ^ x3 ;
  assign n25 = n22 & n24 ;
  assign n26 = n25 ^ x3 ;
  assign n27 = n21 & n26 ;
  assign n28 = n20 & n27 ;
  assign n29 = ~n17 & ~n28 ;
  assign n30 = x0 & x5 ;
  assign n31 = ~x11 & n30 ;
  assign n32 = ~x6 & n31 ;
  assign n33 = x1 & n32 ;
  assign n34 = ~n29 & n33 ;
  assign y0 = n34 ;
endmodule
