module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
  assign n8 = ~x4 & ~x5 ;
  assign n9 = ~x3 & n8 ;
  assign n10 = x2 & ~n9 ;
  assign n11 = ~x0 & x1 ;
  assign n12 = ~n10 & n11 ;
  assign n13 = x2 ^ x0 ;
  assign n14 = ~x1 & n13 ;
  assign n15 = n14 ^ x3 ;
  assign n16 = ~x5 & ~x6 ;
  assign n17 = n16 ^ x4 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = x6 ^ x5 ;
  assign n20 = x5 ^ x0 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = n21 ^ x0 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = ~n18 & ~n23 ;
  assign n25 = n24 ^ n16 ;
  assign n26 = n25 ^ n14 ;
  assign n27 = n15 & n26 ;
  assign n28 = n27 ^ n24 ;
  assign n29 = n28 ^ n16 ;
  assign n30 = n29 ^ x3 ;
  assign n31 = n14 & n30 ;
  assign n32 = n31 ^ n14 ;
  assign n33 = ~n12 & ~n32 ;
  assign y0 = ~n33 ;
endmodule
