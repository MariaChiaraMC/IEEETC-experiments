module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n13 = x0 & ~x8 ;
  assign n16 = ~x4 & x5 ;
  assign n17 = ~x2 & n16 ;
  assign n14 = x7 & ~x11 ;
  assign n15 = x6 & n14 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n19 ^ n13 ;
  assign n21 = x3 ^ x1 ;
  assign n22 = ~x3 & n21 ;
  assign n23 = n22 ^ n15 ;
  assign n24 = n23 ^ x3 ;
  assign n25 = n20 & n24 ;
  assign n26 = n25 ^ n22 ;
  assign n27 = n26 ^ x3 ;
  assign n28 = n13 & ~n27 ;
  assign n29 = n28 ^ n13 ;
  assign y0 = n29 ;
endmodule
