module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n17 = ~x3 & ~x6 ;
  assign n18 = ~x12 & ~x15 ;
  assign n19 = n17 & n18 ;
  assign n20 = x5 & x7 ;
  assign n21 = ~x14 & n20 ;
  assign n22 = n19 & n21 ;
  assign n23 = ~x4 & ~x13 ;
  assign n24 = ~x8 & n23 ;
  assign n25 = ~x9 & ~x11 ;
  assign n26 = ~x10 & n25 ;
  assign n27 = n24 & n26 ;
  assign n28 = n22 & n27 ;
  assign n29 = x0 & ~n28 ;
  assign n30 = x1 & n29 ;
  assign y0 = ~n30 ;
endmodule
