module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 ;
  assign n9 = x5 ^ x2 ;
  assign n11 = n9 ^ x5 ;
  assign n12 = n11 ^ n9 ;
  assign n13 = n9 ^ x0 ;
  assign n14 = ~n12 & n13 ;
  assign n15 = n14 ^ n9 ;
  assign n16 = x1 & ~x6 ;
  assign n17 = ~x1 & x6 ;
  assign n18 = ~n16 & ~n17 ;
  assign n19 = n9 & n18 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = n15 & n20 ;
  assign n8 = x6 ^ x1 ;
  assign n10 = ~n8 & n9 ;
  assign n22 = n21 ^ n10 ;
  assign n23 = x3 & n22 ;
  assign n24 = n23 ^ x3 ;
  assign n25 = n24 ^ x3 ;
  assign n26 = x3 ^ x0 ;
  assign n27 = x4 ^ x1 ;
  assign n28 = ~n26 & ~n27 ;
  assign n29 = x0 & ~x3 ;
  assign n30 = ~n16 & ~n29 ;
  assign n31 = x5 & ~n30 ;
  assign n32 = ~x2 & ~n8 ;
  assign n33 = n31 & ~n32 ;
  assign n34 = x5 & x6 ;
  assign n35 = x3 & ~n34 ;
  assign n36 = ~x2 & ~x5 ;
  assign n37 = x6 & n36 ;
  assign n38 = ~n35 & ~n37 ;
  assign n39 = ~n33 & n38 ;
  assign n40 = n39 ^ x4 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = ~x6 & n36 ;
  assign n43 = n42 ^ n34 ;
  assign n44 = ~x3 & n43 ;
  assign n45 = n44 ^ n34 ;
  assign n46 = n45 ^ n39 ;
  assign n47 = ~n41 & ~n46 ;
  assign n48 = n47 ^ n39 ;
  assign n49 = ~n28 & n48 ;
  assign n50 = ~n25 & n49 ;
  assign y0 = n50 ;
endmodule
