module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 ;
  assign n8 = ~x3 & ~x5 ;
  assign n9 = x3 & x5 ;
  assign n10 = ~n8 & ~n9 ;
  assign n11 = x2 ^ x0 ;
  assign n12 = ~x5 & ~x6 ;
  assign n13 = n12 ^ x2 ;
  assign n14 = n11 & ~n13 ;
  assign n15 = n14 ^ x2 ;
  assign n16 = n10 & ~n15 ;
  assign n17 = ~x1 & n16 ;
  assign n20 = x6 ^ x4 ;
  assign n34 = n20 ^ x6 ;
  assign n18 = ~x0 & ~x2 ;
  assign n19 = n18 ^ x6 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n22 ^ x6 ;
  assign n24 = x5 ^ x3 ;
  assign n25 = x5 ^ x2 ;
  assign n26 = n25 ^ x2 ;
  assign n27 = n11 & ~n26 ;
  assign n28 = n27 ^ x2 ;
  assign n29 = ~n24 & ~n28 ;
  assign n30 = x1 & n29 ;
  assign n31 = n30 ^ n21 ;
  assign n32 = n31 ^ n21 ;
  assign n33 = ~n23 & ~n32 ;
  assign n35 = n34 ^ n33 ;
  assign n36 = x0 & x2 ;
  assign n37 = x1 & ~n10 ;
  assign n38 = n36 & ~n37 ;
  assign n39 = ~x1 & x5 ;
  assign n40 = ~x3 & n39 ;
  assign n41 = x6 & ~n40 ;
  assign n42 = ~n38 & ~n41 ;
  assign n43 = n42 ^ n20 ;
  assign n44 = n34 & ~n43 ;
  assign n45 = n44 ^ n42 ;
  assign n46 = n35 & n45 ;
  assign n47 = n46 ^ n33 ;
  assign n48 = n47 ^ n20 ;
  assign n49 = n48 ^ x4 ;
  assign n50 = n49 ^ x6 ;
  assign n51 = ~n17 & n50 ;
  assign y0 = n51 ;
endmodule
