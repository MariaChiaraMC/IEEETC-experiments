module top( x0 , x1 , x2 , x3 , x4 , y0 );
  input x0 , x1 , x2 , x3 , x4 ;
  output y0 ;
  wire n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n6 = x1 ^ x0 ;
  assign n14 = x2 ^ x1 ;
  assign n15 = n14 ^ x1 ;
  assign n16 = ~n14 & n15 ;
  assign n7 = x3 ^ x2 ;
  assign n8 = n7 ^ x4 ;
  assign n9 = n8 ^ n7 ;
  assign n10 = n7 ^ x2 ;
  assign n11 = n10 ^ x1 ;
  assign n12 = n9 & ~n11 ;
  assign n19 = n16 ^ n12 ;
  assign n13 = n12 ^ n6 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = ~n13 & ~n17 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = ~n6 & n20 ;
  assign n22 = n21 ^ n12 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = n23 ^ n18 ;
  assign y0 = n24 ;
endmodule
