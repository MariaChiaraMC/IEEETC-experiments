module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ;
  assign n8 = ~x0 & ~x1 ;
  assign n9 = x2 & n8 ;
  assign n10 = ~x5 & ~n9 ;
  assign n11 = x4 & ~n10 ;
  assign n12 = ~x3 & ~n11 ;
  assign n14 = ~x4 & ~x5 ;
  assign n13 = x1 ^ x0 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = ~x1 & ~n15 ;
  assign n17 = n16 ^ x1 ;
  assign n18 = n16 ^ x2 ;
  assign n19 = n14 & ~n18 ;
  assign n20 = n19 ^ n14 ;
  assign n21 = n20 ^ n13 ;
  assign n22 = ~n17 & ~n21 ;
  assign n23 = n22 ^ n13 ;
  assign n24 = ~n12 & ~n23 ;
  assign n25 = x0 & x6 ;
  assign n26 = x3 & ~n25 ;
  assign n27 = ~n8 & ~n26 ;
  assign n28 = ~x2 & n27 ;
  assign n29 = ~n24 & ~n28 ;
  assign y0 = ~n29 ;
endmodule
