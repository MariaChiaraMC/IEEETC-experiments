// Benchmark "./inc.pla" written by ABC on Thu Apr 23 10:59:53 2020

module \./inc.pla  ( 
    x0, x1, x2, x3, x4, x5, x6,
    z8  );
  input  x0, x1, x2, x3, x4, x5, x6;
  output z8;
  assign z8 = ~x2 | ~x3;
endmodule


