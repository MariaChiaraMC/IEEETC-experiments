module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n10 = x1 ^ x0 ;
  assign n11 = ~x3 & ~x4 ;
  assign n12 = ~x2 & ~x8 ;
  assign n13 = ~x5 & ~x6 ;
  assign n14 = ~x7 & n13 ;
  assign n15 = n12 & n14 ;
  assign n16 = n11 & n15 ;
  assign n17 = n16 ^ x1 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = x2 & x8 ;
  assign n20 = x3 & x4 ;
  assign n21 = x5 & x6 ;
  assign n22 = n20 & n21 ;
  assign n23 = n19 & n22 ;
  assign n24 = x7 & n23 ;
  assign n25 = n24 ^ n16 ;
  assign n26 = ~n18 & n25 ;
  assign n27 = n26 ^ n16 ;
  assign n28 = ~n10 & ~n27 ;
  assign y0 = ~n28 ;
endmodule
