module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 ;
  assign n17 = x11 & ~x15 ;
  assign n18 = ~x6 & ~x11 ;
  assign n19 = ~x0 & ~x13 ;
  assign n20 = n18 & n19 ;
  assign n21 = ~x14 & n20 ;
  assign n22 = ~x7 & ~x9 ;
  assign n23 = ~x8 & n22 ;
  assign n24 = n23 ^ x10 ;
  assign n25 = n23 ^ x1 ;
  assign n26 = n25 ^ x1 ;
  assign n27 = ~x4 & ~x5 ;
  assign n28 = ~x3 & n27 ;
  assign n29 = ~x2 & n28 ;
  assign n30 = n29 ^ x1 ;
  assign n31 = n26 & n30 ;
  assign n32 = n31 ^ x1 ;
  assign n33 = n24 & ~n32 ;
  assign n34 = n21 & n33 ;
  assign n35 = x12 & n34 ;
  assign n36 = ~n17 & ~n35 ;
  assign y0 = ~n36 ;
endmodule
