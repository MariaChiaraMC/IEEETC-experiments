// Benchmark "./sqr6.pla" written by ABC on Thu Apr 23 11:00:04 2020

module \./sqr6.pla  ( 
    x0, x1, x2, x3, x4, x5,
    z8  );
  input  x0, x1, x2, x3, x4, x5;
  output z8;
  assign z8 = 1'b1;
endmodule


