module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 ;
  assign n11 = ~x1 & ~x7 ;
  assign n12 = ~x9 & n11 ;
  assign n13 = x3 & ~n12 ;
  assign n14 = x1 & x7 ;
  assign n15 = ~x9 & n14 ;
  assign n16 = x7 & x9 ;
  assign n17 = ~x3 & ~n16 ;
  assign n18 = ~x1 & ~n17 ;
  assign n19 = ~n15 & ~n18 ;
  assign n20 = x0 & x8 ;
  assign n21 = x5 & ~x6 ;
  assign n22 = n20 & n21 ;
  assign n23 = x2 & n22 ;
  assign n24 = ~n19 & n23 ;
  assign n25 = ~n13 & n24 ;
  assign n26 = ~x0 & ~x8 ;
  assign n27 = x3 ^ x2 ;
  assign n29 = x5 & ~x7 ;
  assign n28 = x6 ^ x1 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = n27 & ~n30 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = x6 ^ x3 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = ~n28 & ~n34 ;
  assign n36 = n35 ^ n28 ;
  assign n37 = n36 ^ n29 ;
  assign n38 = n32 & ~n37 ;
  assign n39 = n26 & n38 ;
  assign n40 = ~x5 & ~x7 ;
  assign n41 = ~x0 & ~x6 ;
  assign n42 = n40 & n41 ;
  assign n44 = ~x3 & x8 ;
  assign n43 = x3 & ~x8 ;
  assign n45 = n44 ^ n43 ;
  assign n46 = ~x1 & n45 ;
  assign n47 = n46 ^ n44 ;
  assign n48 = n42 & n47 ;
  assign n49 = ~x2 & n48 ;
  assign n50 = x2 & x3 ;
  assign n51 = x0 & x1 ;
  assign n52 = ~x6 & ~x8 ;
  assign n53 = ~x7 & n52 ;
  assign n54 = n51 & n53 ;
  assign n55 = x8 ^ x0 ;
  assign n56 = x7 ^ x1 ;
  assign n57 = n56 ^ x8 ;
  assign n58 = ~n55 & ~n57 ;
  assign n59 = x6 & n58 ;
  assign n60 = ~n54 & ~n59 ;
  assign n61 = n50 & ~n60 ;
  assign n62 = x8 & n41 ;
  assign n63 = x2 & ~n62 ;
  assign n64 = x7 & ~n43 ;
  assign n65 = ~x1 & ~x6 ;
  assign n66 = ~x3 & ~n65 ;
  assign n67 = ~x0 & ~n66 ;
  assign n68 = n64 & ~n67 ;
  assign n69 = ~n63 & n68 ;
  assign n70 = ~x2 & n44 ;
  assign n71 = ~n51 & ~n70 ;
  assign n72 = n71 ^ x8 ;
  assign n73 = n72 ^ n71 ;
  assign n74 = x1 & x3 ;
  assign n75 = x0 & ~n74 ;
  assign n76 = n75 ^ n71 ;
  assign n77 = n76 ^ n71 ;
  assign n78 = n73 & ~n77 ;
  assign n79 = n78 ^ n71 ;
  assign n80 = x6 & n79 ;
  assign n81 = n80 ^ n71 ;
  assign n82 = n69 & n81 ;
  assign n83 = ~n61 & ~n82 ;
  assign n84 = n83 ^ x7 ;
  assign n85 = n84 ^ n83 ;
  assign n86 = x8 ^ x2 ;
  assign n87 = ~x0 & x1 ;
  assign n88 = n87 ^ x8 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = n89 ^ n86 ;
  assign n91 = x3 ^ x0 ;
  assign n92 = ~x3 & n91 ;
  assign n93 = n92 ^ n87 ;
  assign n94 = n93 ^ x3 ;
  assign n95 = n90 & ~n94 ;
  assign n96 = n95 ^ n92 ;
  assign n97 = n96 ^ x3 ;
  assign n98 = ~n86 & ~n97 ;
  assign n99 = x6 & n98 ;
  assign n100 = x8 ^ x3 ;
  assign n101 = x6 ^ x2 ;
  assign n102 = n101 ^ n55 ;
  assign n103 = n102 ^ n100 ;
  assign n104 = n101 ^ x6 ;
  assign n105 = n101 ^ x8 ;
  assign n106 = n105 ^ n104 ;
  assign n107 = n104 & n106 ;
  assign n108 = n107 ^ n101 ;
  assign n109 = n108 ^ n104 ;
  assign n110 = ~n103 & ~n109 ;
  assign n111 = n110 ^ n107 ;
  assign n112 = n111 ^ n104 ;
  assign n113 = n100 & n112 ;
  assign n114 = ~x1 & n113 ;
  assign n115 = ~n99 & ~n114 ;
  assign n116 = n115 ^ n83 ;
  assign n117 = n116 ^ n83 ;
  assign n118 = n85 & ~n117 ;
  assign n119 = n118 ^ n83 ;
  assign n120 = ~x5 & ~n119 ;
  assign n121 = n120 ^ n83 ;
  assign n122 = ~n49 & n121 ;
  assign n123 = n122 ^ x9 ;
  assign n124 = n123 ^ n122 ;
  assign n125 = n124 ^ n39 ;
  assign n126 = x5 & ~n43 ;
  assign n127 = ~n50 & n126 ;
  assign n128 = n53 ^ x2 ;
  assign n129 = n128 ^ n53 ;
  assign n130 = x7 & ~x8 ;
  assign n131 = x0 & x6 ;
  assign n132 = ~x3 & n131 ;
  assign n133 = n130 & n132 ;
  assign n134 = ~x0 & x3 ;
  assign n135 = ~x7 & n134 ;
  assign n136 = ~x6 & n135 ;
  assign n137 = ~n133 & ~n136 ;
  assign n138 = n137 ^ n53 ;
  assign n139 = ~n129 & ~n138 ;
  assign n140 = n139 ^ n53 ;
  assign n141 = n127 & n140 ;
  assign n142 = ~x1 & ~n141 ;
  assign n143 = ~x0 & ~x2 ;
  assign n144 = x6 & x7 ;
  assign n145 = n143 & n144 ;
  assign n146 = ~x2 & x6 ;
  assign n147 = ~x5 & x6 ;
  assign n148 = ~x2 & x5 ;
  assign n149 = ~x7 & n148 ;
  assign n150 = ~n147 & ~n149 ;
  assign n151 = x0 & ~n150 ;
  assign n152 = ~n146 & n151 ;
  assign n153 = ~n145 & ~n152 ;
  assign n154 = n44 & ~n153 ;
  assign n164 = n131 ^ x6 ;
  assign n165 = ~x5 & ~n164 ;
  assign n166 = n165 ^ x6 ;
  assign n155 = x7 ^ x6 ;
  assign n156 = x7 ^ x3 ;
  assign n157 = n156 ^ x3 ;
  assign n158 = ~n91 & ~n157 ;
  assign n159 = n158 ^ x3 ;
  assign n160 = n155 & n159 ;
  assign n161 = n148 & n160 ;
  assign n167 = n166 ^ n161 ;
  assign n168 = n167 ^ n161 ;
  assign n162 = n161 ^ n50 ;
  assign n163 = n162 ^ n161 ;
  assign n169 = n168 ^ n163 ;
  assign n170 = n161 ^ x7 ;
  assign n171 = n170 ^ n161 ;
  assign n172 = n171 ^ n168 ;
  assign n173 = ~n168 & ~n172 ;
  assign n174 = n173 ^ n168 ;
  assign n175 = ~n169 & ~n174 ;
  assign n176 = n175 ^ n173 ;
  assign n177 = n176 ^ n161 ;
  assign n178 = n177 ^ n168 ;
  assign n179 = ~x8 & ~n178 ;
  assign n180 = n179 ^ n161 ;
  assign n181 = ~n154 & ~n180 ;
  assign n182 = x1 & n181 ;
  assign n183 = n182 ^ n142 ;
  assign n184 = ~n142 & n183 ;
  assign n185 = n184 ^ n122 ;
  assign n186 = n185 ^ n142 ;
  assign n187 = n125 & n186 ;
  assign n188 = n187 ^ n184 ;
  assign n189 = n188 ^ n142 ;
  assign n190 = ~n39 & ~n189 ;
  assign n191 = n190 ^ n39 ;
  assign n192 = n191 ^ x4 ;
  assign n193 = n192 ^ n191 ;
  assign n214 = ~x3 & ~x5 ;
  assign n234 = x7 & n214 ;
  assign n235 = x3 & x5 ;
  assign n236 = x9 & n235 ;
  assign n237 = ~n234 & ~n236 ;
  assign n238 = ~n16 & n62 ;
  assign n239 = ~n237 & n238 ;
  assign n256 = ~x8 & x9 ;
  assign n265 = n42 & n256 ;
  assign n266 = ~x3 & n265 ;
  assign n267 = ~x7 & ~n43 ;
  assign n268 = ~n214 & n267 ;
  assign n269 = x6 & ~n235 ;
  assign n270 = n268 & n269 ;
  assign n271 = ~n131 & ~n270 ;
  assign n254 = x5 & x8 ;
  assign n255 = x7 & n254 ;
  assign n272 = ~x5 & x7 ;
  assign n273 = n43 & n272 ;
  assign n274 = x0 & ~n273 ;
  assign n275 = ~n255 & n274 ;
  assign n276 = n275 ^ x9 ;
  assign n277 = n276 ^ n275 ;
  assign n278 = n275 ^ x8 ;
  assign n279 = n277 & ~n278 ;
  assign n280 = n279 ^ n275 ;
  assign n281 = ~n271 & ~n280 ;
  assign n282 = ~n266 & ~n281 ;
  assign n215 = x5 & x6 ;
  assign n243 = ~x7 & n215 ;
  assign n244 = ~n42 & ~n243 ;
  assign n240 = x6 ^ x0 ;
  assign n241 = n155 & n240 ;
  assign n242 = n241 ^ x0 ;
  assign n245 = n244 ^ n242 ;
  assign n246 = n245 ^ n244 ;
  assign n247 = n244 ^ x5 ;
  assign n248 = n247 ^ n244 ;
  assign n249 = ~n246 & n248 ;
  assign n250 = n249 ^ n244 ;
  assign n251 = x9 & ~n250 ;
  assign n252 = n251 ^ n244 ;
  assign n253 = n43 & ~n252 ;
  assign n257 = n40 & n256 ;
  assign n258 = ~n255 & ~n257 ;
  assign n259 = n132 & ~n258 ;
  assign n222 = ~x6 & x7 ;
  assign n260 = x8 & n214 ;
  assign n261 = n222 & n260 ;
  assign n262 = ~x9 & n261 ;
  assign n263 = ~n259 & ~n262 ;
  assign n264 = ~n253 & n263 ;
  assign n283 = n282 ^ n264 ;
  assign n284 = n283 ^ n264 ;
  assign n285 = ~x7 & n214 ;
  assign n286 = x9 & ~n285 ;
  assign n287 = n286 ^ n264 ;
  assign n288 = n287 ^ n264 ;
  assign n289 = ~n284 & ~n288 ;
  assign n290 = n289 ^ n264 ;
  assign n291 = x1 & ~n290 ;
  assign n292 = n291 ^ n264 ;
  assign n293 = ~n239 & n292 ;
  assign n194 = n134 & n147 ;
  assign n195 = n14 & n194 ;
  assign n196 = x9 & ~n195 ;
  assign n211 = x6 & x8 ;
  assign n212 = n29 & n134 ;
  assign n213 = n211 & n212 ;
  assign n216 = n20 & ~n215 ;
  assign n217 = ~n214 & n216 ;
  assign n218 = n217 ^ x3 ;
  assign n219 = x6 & ~x7 ;
  assign n220 = n219 ^ n217 ;
  assign n221 = n220 ^ n219 ;
  assign n223 = n26 & n222 ;
  assign n224 = n223 ^ n219 ;
  assign n225 = ~n221 & ~n224 ;
  assign n226 = n225 ^ n219 ;
  assign n227 = ~n218 & n226 ;
  assign n228 = n227 ^ x3 ;
  assign n229 = ~n213 & n228 ;
  assign n197 = x5 ^ x3 ;
  assign n198 = x5 ^ x0 ;
  assign n199 = n198 ^ x7 ;
  assign n200 = n199 ^ x6 ;
  assign n201 = n200 ^ n197 ;
  assign n202 = n155 ^ x0 ;
  assign n203 = x0 & ~n202 ;
  assign n204 = n203 ^ x6 ;
  assign n205 = n204 ^ x0 ;
  assign n206 = ~n201 & n205 ;
  assign n207 = n206 ^ n203 ;
  assign n208 = n207 ^ x0 ;
  assign n209 = ~n197 & n208 ;
  assign n210 = ~x8 & n209 ;
  assign n230 = n229 ^ n210 ;
  assign n231 = x1 & ~n230 ;
  assign n232 = n231 ^ n229 ;
  assign n233 = n196 & n232 ;
  assign n294 = n293 ^ n233 ;
  assign n295 = n294 ^ n293 ;
  assign n296 = n51 & n222 ;
  assign n297 = n11 & n211 ;
  assign n298 = ~n296 & ~n297 ;
  assign n299 = x5 & ~n298 ;
  assign n300 = n211 ^ x5 ;
  assign n301 = n300 ^ n211 ;
  assign n302 = n211 ^ n52 ;
  assign n303 = n302 ^ n211 ;
  assign n304 = ~n301 & n303 ;
  assign n305 = n304 ^ n211 ;
  assign n306 = ~x7 & n305 ;
  assign n307 = n306 ^ n211 ;
  assign n308 = n87 & n307 ;
  assign n309 = n26 & ~n144 ;
  assign n310 = ~x1 & n309 ;
  assign n311 = x6 ^ x5 ;
  assign n312 = n310 & n311 ;
  assign n313 = ~n308 & ~n312 ;
  assign n314 = ~n299 & n313 ;
  assign n315 = ~x3 & ~n314 ;
  assign n323 = x5 & ~n51 ;
  assign n324 = ~n52 & ~n323 ;
  assign n325 = x7 & ~n324 ;
  assign n316 = x0 & x3 ;
  assign n320 = ~n87 & ~n316 ;
  assign n321 = n320 ^ n211 ;
  assign n317 = n40 & n316 ;
  assign n318 = ~n52 & n317 ;
  assign n319 = n318 ^ n211 ;
  assign n322 = n321 ^ n319 ;
  assign n326 = n325 ^ n322 ;
  assign n327 = n326 ^ n322 ;
  assign n328 = n322 ^ n319 ;
  assign n329 = n328 ^ n211 ;
  assign n330 = n327 & ~n329 ;
  assign n331 = n330 ^ n319 ;
  assign n332 = ~x5 & n51 ;
  assign n333 = ~n319 & n332 ;
  assign n334 = n333 ^ n211 ;
  assign n335 = ~n331 & ~n334 ;
  assign n336 = n335 ^ n333 ;
  assign n337 = ~n211 & n336 ;
  assign n338 = n337 ^ n330 ;
  assign n339 = n338 ^ n318 ;
  assign n340 = n339 ^ n319 ;
  assign n341 = ~n315 & n340 ;
  assign n342 = ~x9 & n341 ;
  assign n343 = n342 ^ n293 ;
  assign n344 = n343 ^ n293 ;
  assign n345 = ~n295 & ~n344 ;
  assign n346 = n345 ^ n293 ;
  assign n347 = x2 & ~n346 ;
  assign n348 = n347 ^ n293 ;
  assign n349 = n348 ^ n191 ;
  assign n350 = n193 & ~n349 ;
  assign n351 = n350 ^ n191 ;
  assign n352 = ~n25 & ~n351 ;
  assign y0 = ~n352 ;
endmodule
