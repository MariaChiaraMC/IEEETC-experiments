module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;
  assign n11 = ~x1 & ~x2 ;
  assign n12 = ~x6 & ~x7 ;
  assign n13 = x4 & x5 ;
  assign n14 = n12 & n13 ;
  assign n15 = n11 & n14 ;
  assign n16 = x7 ^ x6 ;
  assign n17 = x2 & ~x5 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = x4 ^ x1 ;
  assign n20 = x7 ^ x4 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = n18 & ~n23 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = n26 ^ n17 ;
  assign n28 = n16 & ~n27 ;
  assign n29 = n28 ^ n16 ;
  assign n30 = ~n15 & ~n29 ;
  assign n9 = ~x2 & x6 ;
  assign n10 = x7 & n9 ;
  assign n31 = n30 ^ n10 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = x5 ^ x4 ;
  assign n34 = ~x5 & ~n33 ;
  assign n35 = x1 & n34 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = n37 ^ n30 ;
  assign n39 = n32 & ~n38 ;
  assign n40 = n39 ^ n30 ;
  assign n41 = x3 & ~n40 ;
  assign n42 = n41 ^ n30 ;
  assign n43 = ~x0 & ~n42 ;
  assign y0 = n43 ;
endmodule
