module top( x0 , x1 , x2 , x3 , y0 );
  input x0 , x1 , x2 , x3 ;
  output y0 ;
  wire n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n6 = x2 ^ x1 ;
  assign n11 = n6 ^ x2 ;
  assign n5 = x2 ^ x0 ;
  assign n7 = n6 ^ n5 ;
  assign n8 = n7 ^ x3 ;
  assign n9 = n8 ^ n7 ;
  assign n10 = n9 ^ x2 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = n7 ^ n6 ;
  assign n14 = n13 ^ x2 ;
  assign n15 = n14 ^ x2 ;
  assign n16 = ~n9 & ~n15 ;
  assign n17 = n16 ^ n9 ;
  assign n18 = ~n14 & ~n17 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = n12 & n19 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = n21 ^ x2 ;
  assign n23 = n22 ^ x0 ;
  assign n24 = n23 ^ n11 ;
  assign y0 = n24 ;
endmodule
