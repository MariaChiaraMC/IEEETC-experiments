module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 ;
  assign n8 = x4 ^ x3 ;
  assign n9 = n8 ^ x5 ;
  assign n10 = ~x2 & x4 ;
  assign n11 = ~x1 & ~n10 ;
  assign n12 = x0 & ~n11 ;
  assign n13 = n12 ^ x4 ;
  assign n14 = n13 ^ x4 ;
  assign n15 = x5 ^ x4 ;
  assign n16 = n15 ^ x4 ;
  assign n17 = ~n14 & ~n16 ;
  assign n18 = n17 ^ x4 ;
  assign n19 = ~x2 & ~x4 ;
  assign n20 = n19 ^ n9 ;
  assign n21 = ~n18 & ~n20 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = ~n9 & n22 ;
  assign n24 = n23 ^ x4 ;
  assign n25 = n24 ^ n9 ;
  assign n26 = x6 & n25 ;
  assign y0 = n26 ;
endmodule
