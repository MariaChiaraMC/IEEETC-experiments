module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 ;
  assign n15 = ~x4 & x6 ;
  assign n13 = ~x1 & ~x3 ;
  assign n9 = x5 & x7 ;
  assign n10 = x5 & x6 ;
  assign n11 = ~n9 & ~n10 ;
  assign n12 = x3 & ~n11 ;
  assign n14 = n13 ^ n12 ;
  assign n16 = n15 ^ n14 ;
  assign n24 = n16 ^ n14 ;
  assign n17 = ~x5 & ~x6 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = n18 ^ n14 ;
  assign n20 = n16 ^ n12 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n19 & ~n22 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ n19 ;
  assign n27 = n14 ^ n9 ;
  assign n28 = n23 ^ n19 ;
  assign n29 = ~n27 & n28 ;
  assign n30 = n29 ^ n14 ;
  assign n31 = ~n26 & n30 ;
  assign n32 = n31 ^ n14 ;
  assign n33 = n32 ^ n13 ;
  assign n34 = n33 ^ n14 ;
  assign n35 = ~x2 & n34 ;
  assign n36 = ~x4 & ~x6 ;
  assign n37 = x2 & n36 ;
  assign n38 = ~x2 & ~x3 ;
  assign n39 = ~x1 & ~x5 ;
  assign n40 = n38 & n39 ;
  assign n41 = x4 & n40 ;
  assign n42 = ~n37 & ~n41 ;
  assign n43 = ~x7 & ~n42 ;
  assign n44 = x2 & ~x3 ;
  assign n45 = ~x1 & ~n44 ;
  assign n46 = x4 & ~n45 ;
  assign n47 = ~n11 & n46 ;
  assign n48 = ~n43 & ~n47 ;
  assign n49 = x3 ^ x1 ;
  assign n57 = x6 & n49 ;
  assign n50 = n49 ^ x2 ;
  assign n51 = n50 ^ x3 ;
  assign n52 = n51 ^ x3 ;
  assign n53 = n52 ^ x4 ;
  assign n54 = n51 ^ x4 ;
  assign n55 = n54 ^ n49 ;
  assign n56 = n53 & n55 ;
  assign n58 = n57 ^ n56 ;
  assign n59 = n58 ^ n51 ;
  assign n60 = n57 ^ n51 ;
  assign n61 = n51 ^ x5 ;
  assign n62 = n61 ^ n56 ;
  assign n63 = n62 ^ n53 ;
  assign n64 = n60 & n63 ;
  assign n65 = n64 ^ n49 ;
  assign n66 = n59 & n65 ;
  assign n67 = n66 ^ n57 ;
  assign n68 = n67 ^ n64 ;
  assign n69 = n68 ^ x1 ;
  assign n70 = n48 & ~n69 ;
  assign n71 = ~n35 & n70 ;
  assign n72 = ~x0 & ~n71 ;
  assign y0 = n72 ;
endmodule
