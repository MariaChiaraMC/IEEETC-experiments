module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 ;
  assign n19 = ~x3 & ~x4 ;
  assign n17 = ~x2 & x6 ;
  assign n20 = n19 ^ n17 ;
  assign n16 = ~x1 & ~x2 ;
  assign n18 = n17 ^ n16 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n21 ^ x5 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n23 ^ n17 ;
  assign n25 = x1 & x2 ;
  assign n26 = x3 & ~n25 ;
  assign n27 = n26 ^ n22 ;
  assign n28 = ~x5 & ~n27 ;
  assign n29 = n20 ^ n17 ;
  assign n30 = n23 & n29 ;
  assign n31 = n30 ^ n24 ;
  assign n32 = n28 & ~n31 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = ~n24 & n33 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n35 ^ n19 ;
  assign n37 = ~x10 & n36 ;
  assign n38 = x3 & x6 ;
  assign n39 = x5 & ~n38 ;
  assign n40 = n25 & n39 ;
  assign n41 = n40 ^ x4 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = ~x5 & n38 ;
  assign n44 = x5 & ~x6 ;
  assign n45 = x1 & ~n44 ;
  assign n46 = n45 ^ x3 ;
  assign n47 = n45 ^ x10 ;
  assign n48 = n47 ^ x10 ;
  assign n49 = ~x13 & ~x14 ;
  assign n50 = ~x12 & n49 ;
  assign n51 = ~x8 & ~x11 ;
  assign n52 = x10 ^ x9 ;
  assign n53 = x9 ^ x7 ;
  assign n54 = ~n52 & n53 ;
  assign n55 = n54 ^ x9 ;
  assign n56 = n51 & n55 ;
  assign n57 = n50 & n56 ;
  assign n58 = x6 & ~n57 ;
  assign n59 = x2 & ~n58 ;
  assign n60 = n59 ^ x10 ;
  assign n61 = n48 & n60 ;
  assign n62 = n61 ^ x10 ;
  assign n63 = ~n46 & ~n62 ;
  assign n64 = n63 ^ x3 ;
  assign n65 = ~n43 & ~n64 ;
  assign n66 = n65 ^ n40 ;
  assign n67 = n42 & ~n66 ;
  assign n68 = n67 ^ n40 ;
  assign n69 = ~n37 & ~n68 ;
  assign n70 = ~x0 & ~n69 ;
  assign y0 = n70 ;
endmodule
