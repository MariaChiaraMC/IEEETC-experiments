module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
  assign n13 = ~x0 & ~x3 ;
  assign n14 = ~x2 & n13 ;
  assign n15 = ~x1 & n14 ;
  assign n16 = ~x4 & n15 ;
  assign n17 = x5 & ~x6 ;
  assign n18 = ~x5 & x6 ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = ~x8 & ~x9 ;
  assign n21 = n18 & n20 ;
  assign n22 = x11 ^ x10 ;
  assign n23 = n21 & n22 ;
  assign n24 = ~n19 & ~n23 ;
  assign n25 = n23 ^ x7 ;
  assign n26 = ~x10 & ~x11 ;
  assign n27 = ~n17 & ~n26 ;
  assign n28 = x9 ^ x8 ;
  assign n29 = ~n27 & n28 ;
  assign n30 = n29 ^ n24 ;
  assign n31 = ~n25 & n30 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = n24 & n32 ;
  assign n34 = n33 ^ n23 ;
  assign n35 = n16 & n34 ;
  assign y0 = n35 ;
endmodule
