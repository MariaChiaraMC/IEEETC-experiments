module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 ;
  output y0 ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 ;
  assign n20 = ~x3 & ~x15 ;
  assign n22 = n20 ^ x18 ;
  assign n32 = n22 ^ n20 ;
  assign n21 = n20 ^ x7 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n24 ^ n20 ;
  assign n26 = x16 ^ x6 ;
  assign n27 = ~x8 & ~n26 ;
  assign n28 = n27 ^ n23 ;
  assign n29 = n28 ^ n23 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = n25 & n30 ;
  assign n33 = n32 ^ n31 ;
  assign n34 = n33 ^ n25 ;
  assign n35 = ~x2 & ~x10 ;
  assign n36 = x15 & n35 ;
  assign n37 = ~x9 & n36 ;
  assign n38 = n37 ^ n23 ;
  assign n39 = n38 ^ n23 ;
  assign n40 = n39 ^ n32 ;
  assign n41 = n40 ^ n25 ;
  assign n42 = ~x4 & ~n41 ;
  assign n43 = n42 ^ n29 ;
  assign n44 = n39 ^ n20 ;
  assign n45 = n44 ^ n29 ;
  assign n46 = n32 & n45 ;
  assign n47 = n46 ^ n32 ;
  assign n48 = n43 & n47 ;
  assign n49 = n48 ^ n39 ;
  assign n50 = n49 ^ n29 ;
  assign n51 = n34 & ~n50 ;
  assign n52 = n51 ^ n46 ;
  assign n53 = n52 ^ n48 ;
  assign n54 = n53 ^ x18 ;
  assign n55 = n54 ^ n32 ;
  assign n56 = x17 & n55 ;
  assign n82 = x16 & ~x17 ;
  assign n77 = ~n26 & n35 ;
  assign n78 = n77 ^ x16 ;
  assign n79 = x17 & n78 ;
  assign n80 = n79 ^ x16 ;
  assign n81 = x8 & n80 ;
  assign n83 = n82 ^ n81 ;
  assign n84 = n83 ^ x7 ;
  assign n94 = n84 ^ n83 ;
  assign n85 = x6 & ~x9 ;
  assign n86 = ~x8 & ~n85 ;
  assign n87 = n35 & ~n86 ;
  assign n88 = n87 ^ n84 ;
  assign n89 = n88 ^ n83 ;
  assign n90 = n84 ^ n81 ;
  assign n91 = n90 ^ n87 ;
  assign n92 = n91 ^ n89 ;
  assign n93 = ~n89 & ~n92 ;
  assign n95 = n94 ^ n93 ;
  assign n96 = n95 ^ n89 ;
  assign n97 = n83 ^ x6 ;
  assign n98 = n93 ^ n89 ;
  assign n99 = ~n97 & ~n98 ;
  assign n100 = n99 ^ n83 ;
  assign n101 = n96 & n100 ;
  assign n102 = n101 ^ n83 ;
  assign n103 = n102 ^ n82 ;
  assign n104 = n103 ^ n83 ;
  assign n57 = x13 ^ x11 ;
  assign n58 = ~x12 & x13 ;
  assign n59 = n57 & n58 ;
  assign n60 = n59 ^ n57 ;
  assign n61 = x1 & n60 ;
  assign n62 = n61 ^ x16 ;
  assign n63 = n62 ^ n61 ;
  assign n64 = n63 ^ x17 ;
  assign n65 = x4 & x7 ;
  assign n66 = ~x6 & x8 ;
  assign n67 = n65 & n66 ;
  assign n68 = n67 ^ x3 ;
  assign n69 = ~x3 & n68 ;
  assign n70 = n69 ^ n61 ;
  assign n71 = n70 ^ x3 ;
  assign n72 = ~n64 & n71 ;
  assign n73 = n72 ^ n69 ;
  assign n74 = n73 ^ x3 ;
  assign n75 = ~x17 & ~n74 ;
  assign n76 = n75 ^ x17 ;
  assign n105 = n104 ^ n76 ;
  assign n106 = ~x15 & ~n105 ;
  assign n107 = n106 ^ n104 ;
  assign n108 = ~x18 & n107 ;
  assign n109 = ~n56 & ~n108 ;
  assign n110 = ~x14 & ~n109 ;
  assign n111 = ~x9 & n65 ;
  assign n112 = ~x14 & ~n111 ;
  assign n113 = x8 & ~n26 ;
  assign n114 = n113 ^ x18 ;
  assign n115 = n114 ^ x17 ;
  assign n116 = x14 ^ x7 ;
  assign n117 = x18 & n116 ;
  assign n118 = n117 ^ x7 ;
  assign n119 = n115 & ~n118 ;
  assign n120 = n119 ^ n117 ;
  assign n121 = n120 ^ x7 ;
  assign n122 = n121 ^ x18 ;
  assign n123 = x17 & ~n122 ;
  assign n124 = ~n112 & n123 ;
  assign n125 = ~x18 & n82 ;
  assign n126 = n125 ^ n116 ;
  assign n127 = x4 & n85 ;
  assign n128 = ~x8 & n127 ;
  assign n129 = n128 ^ n66 ;
  assign n130 = x14 & n129 ;
  assign n131 = n130 ^ n128 ;
  assign n132 = ~n126 & n131 ;
  assign n133 = n132 ^ n130 ;
  assign n134 = n133 ^ n128 ;
  assign n135 = n134 ^ x14 ;
  assign n136 = n125 & n135 ;
  assign n137 = ~n124 & ~n136 ;
  assign n138 = ~x15 & ~n137 ;
  assign n139 = ~n110 & ~n138 ;
  assign n140 = ~x0 & ~n139 ;
  assign y0 = n140 ;
endmodule
