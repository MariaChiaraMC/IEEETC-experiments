module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 ;
  assign n9 = x1 & ~x5 ;
  assign n11 = x4 & ~x6 ;
  assign n10 = x6 & ~x7 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = n12 ^ n11 ;
  assign n14 = n11 ^ x4 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = n13 & ~n15 ;
  assign n17 = n16 ^ n11 ;
  assign n18 = x3 & n17 ;
  assign n19 = n18 ^ n11 ;
  assign n20 = n9 & n19 ;
  assign n21 = n20 ^ x2 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n22 ^ x0 ;
  assign n24 = ~x1 & x7 ;
  assign n25 = x6 & n24 ;
  assign n26 = ~x3 & x4 ;
  assign n27 = x3 & ~x4 ;
  assign n28 = ~x5 & n27 ;
  assign n29 = ~n26 & ~n28 ;
  assign n30 = n25 & ~n29 ;
  assign n31 = x3 & n11 ;
  assign n32 = x7 & n31 ;
  assign n33 = n9 & n32 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = ~n30 & n34 ;
  assign n36 = n35 ^ n20 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = n23 & n37 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n39 ^ n30 ;
  assign n41 = x0 & ~n40 ;
  assign n42 = n41 ^ x0 ;
  assign n43 = x2 & x3 ;
  assign n44 = n11 & n24 ;
  assign n45 = n43 & n44 ;
  assign n67 = ~x2 & x3 ;
  assign n63 = ~x6 & ~x7 ;
  assign n75 = x6 ^ x1 ;
  assign n76 = n75 ^ x7 ;
  assign n77 = n63 & ~n76 ;
  assign n78 = n77 ^ n76 ;
  assign n79 = x4 & ~n78 ;
  assign n61 = ~x4 & ~x6 ;
  assign n80 = ~x1 & n61 ;
  assign n81 = x7 & n80 ;
  assign n82 = ~n79 & ~n81 ;
  assign n83 = n67 & ~n82 ;
  assign n84 = ~x6 & x7 ;
  assign n85 = x2 & ~x3 ;
  assign n86 = n84 & n85 ;
  assign n87 = ~x4 & x6 ;
  assign n88 = ~x2 & ~n87 ;
  assign n89 = ~x7 & ~n27 ;
  assign n90 = ~x1 & ~n11 ;
  assign n91 = n89 & n90 ;
  assign n92 = ~n88 & n91 ;
  assign n93 = ~n86 & ~n92 ;
  assign n94 = ~n83 & n93 ;
  assign n46 = x3 ^ x2 ;
  assign n47 = n46 ^ x4 ;
  assign n48 = x4 ^ x3 ;
  assign n49 = n48 ^ x4 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = x6 ^ x4 ;
  assign n52 = n51 ^ x1 ;
  assign n53 = x1 & n52 ;
  assign n54 = n53 ^ x4 ;
  assign n55 = n54 ^ x1 ;
  assign n56 = ~n50 & n55 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n57 ^ x1 ;
  assign n59 = n47 & n58 ;
  assign n60 = x7 & n59 ;
  assign n62 = x2 & ~n61 ;
  assign n64 = n63 ^ n62 ;
  assign n65 = n62 ^ n27 ;
  assign n66 = n65 ^ n27 ;
  assign n68 = n67 ^ n27 ;
  assign n69 = ~n66 & ~n68 ;
  assign n70 = n69 ^ n27 ;
  assign n71 = n64 & n70 ;
  assign n72 = n71 ^ n63 ;
  assign n73 = ~x1 & n72 ;
  assign n74 = ~n60 & ~n73 ;
  assign n95 = n94 ^ n74 ;
  assign n96 = ~x0 & n95 ;
  assign n97 = n96 ^ n94 ;
  assign n98 = ~n45 & n97 ;
  assign n99 = n98 ^ x5 ;
  assign n100 = n99 ^ n98 ;
  assign n101 = x2 & ~x7 ;
  assign n102 = ~n31 & ~n87 ;
  assign n103 = n102 ^ n61 ;
  assign n104 = x1 & ~n103 ;
  assign n105 = n104 ^ n61 ;
  assign n106 = n101 & n105 ;
  assign n107 = ~x1 & x6 ;
  assign n108 = ~n26 & ~n43 ;
  assign n109 = ~n89 & n108 ;
  assign n110 = n107 & n109 ;
  assign n111 = ~n106 & ~n110 ;
  assign n112 = ~x0 & ~n111 ;
  assign n113 = ~x2 & ~x3 ;
  assign n114 = n44 & n113 ;
  assign n115 = ~n112 & ~n114 ;
  assign n116 = n115 ^ n98 ;
  assign n117 = ~n100 & n116 ;
  assign n118 = n117 ^ n98 ;
  assign n119 = ~n42 & n118 ;
  assign y0 = ~n119 ;
endmodule
