module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 ;
  assign n10 = ~x2 & ~x3 ;
  assign n11 = ~x5 & ~x7 ;
  assign n12 = n11 ^ x6 ;
  assign n13 = n12 ^ x0 ;
  assign n22 = n13 ^ n12 ;
  assign n14 = ~x7 & x8 ;
  assign n15 = ~x5 & n14 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = n16 ^ n12 ;
  assign n18 = n13 ^ n11 ;
  assign n19 = n18 ^ n15 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n17 & ~n20 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n23 ^ n17 ;
  assign n25 = n12 ^ x5 ;
  assign n26 = n21 ^ n17 ;
  assign n27 = ~n25 & n26 ;
  assign n28 = n27 ^ n12 ;
  assign n29 = ~n24 & n28 ;
  assign n30 = n29 ^ n12 ;
  assign n31 = n30 ^ x6 ;
  assign n32 = n31 ^ n12 ;
  assign n33 = x4 & n32 ;
  assign n52 = x5 & ~x8 ;
  assign n53 = ~x4 & n11 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = x0 & ~n54 ;
  assign n34 = ~x5 & ~x8 ;
  assign n35 = ~x4 & ~n34 ;
  assign n37 = n35 ^ x7 ;
  assign n36 = n35 ^ x0 ;
  assign n38 = n37 ^ n36 ;
  assign n39 = n38 ^ x8 ;
  assign n40 = ~x4 & ~x5 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n37 ^ n35 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = ~n41 & ~n43 ;
  assign n45 = n44 ^ n37 ;
  assign n46 = n45 ^ n41 ;
  assign n47 = n39 & ~n46 ;
  assign n48 = n47 ^ n44 ;
  assign n49 = n48 ^ n41 ;
  assign n50 = x8 & ~n49 ;
  assign n51 = n50 ^ n35 ;
  assign n56 = n55 ^ n51 ;
  assign n57 = n56 ^ n51 ;
  assign n58 = x7 & x8 ;
  assign n59 = ~x4 & x5 ;
  assign n60 = n58 & n59 ;
  assign n61 = n60 ^ n51 ;
  assign n62 = n61 ^ n51 ;
  assign n63 = ~n57 & ~n62 ;
  assign n64 = n63 ^ n51 ;
  assign n65 = x6 & ~n64 ;
  assign n66 = n65 ^ n51 ;
  assign n67 = ~n33 & ~n66 ;
  assign n68 = n10 & ~n67 ;
  assign n69 = n68 ^ x0 ;
  assign n70 = n69 ^ x1 ;
  assign n192 = n70 ^ n69 ;
  assign n71 = x3 ^ x2 ;
  assign n72 = x5 & ~x6 ;
  assign n73 = n58 & n72 ;
  assign n74 = ~n15 & ~n73 ;
  assign n75 = n74 ^ n71 ;
  assign n76 = n75 ^ x3 ;
  assign n77 = n76 ^ n75 ;
  assign n78 = x7 & ~x8 ;
  assign n79 = x6 & n78 ;
  assign n80 = ~x7 & ~x8 ;
  assign n81 = ~x3 & ~x6 ;
  assign n82 = n80 & n81 ;
  assign n83 = ~n79 & ~n82 ;
  assign n84 = x5 & x7 ;
  assign n85 = ~x3 & n84 ;
  assign n86 = ~n15 & ~n85 ;
  assign n87 = x6 & ~n86 ;
  assign n88 = n83 & ~n87 ;
  assign n89 = n88 ^ n75 ;
  assign n90 = n89 ^ n71 ;
  assign n91 = n77 & ~n90 ;
  assign n92 = n91 ^ n88 ;
  assign n93 = ~x6 & x8 ;
  assign n94 = ~x7 & n93 ;
  assign n95 = n88 & ~n94 ;
  assign n96 = n95 ^ n71 ;
  assign n97 = n92 & ~n96 ;
  assign n98 = n97 ^ n95 ;
  assign n99 = ~n71 & n98 ;
  assign n100 = n99 ^ n91 ;
  assign n101 = n100 ^ x2 ;
  assign n102 = n101 ^ n88 ;
  assign n103 = x4 & n102 ;
  assign n104 = x3 & ~x5 ;
  assign n105 = ~n79 & ~n94 ;
  assign n106 = n104 & ~n105 ;
  assign n107 = ~n103 & ~n106 ;
  assign n108 = ~x2 & x3 ;
  assign n109 = ~x5 & x6 ;
  assign n110 = ~x4 & n109 ;
  assign n111 = ~n73 & ~n110 ;
  assign n112 = n108 & ~n111 ;
  assign n113 = n93 ^ n78 ;
  assign n114 = n113 ^ n93 ;
  assign n115 = n93 ^ x5 ;
  assign n116 = n115 ^ n93 ;
  assign n117 = n114 & ~n116 ;
  assign n118 = n117 ^ n93 ;
  assign n119 = ~x4 & n118 ;
  assign n120 = n119 ^ n93 ;
  assign n121 = x3 & n120 ;
  assign n122 = ~n112 & ~n121 ;
  assign n123 = n52 ^ x5 ;
  assign n124 = n123 ^ n52 ;
  assign n125 = x6 & ~x7 ;
  assign n126 = n125 ^ n52 ;
  assign n127 = n126 ^ n52 ;
  assign n128 = ~n124 & ~n127 ;
  assign n129 = n128 ^ n52 ;
  assign n130 = x3 & n129 ;
  assign n131 = n130 ^ n52 ;
  assign n132 = x4 & n131 ;
  assign n133 = n14 & n59 ;
  assign n134 = ~x5 & n58 ;
  assign n135 = ~x6 & n134 ;
  assign n136 = ~n133 & ~n135 ;
  assign n137 = n83 & n136 ;
  assign n138 = ~n132 & n137 ;
  assign n139 = n138 ^ x2 ;
  assign n140 = n139 ^ n138 ;
  assign n141 = x4 & n72 ;
  assign n142 = x8 & n141 ;
  assign n143 = n142 ^ n138 ;
  assign n144 = ~n140 & ~n143 ;
  assign n145 = n144 ^ n138 ;
  assign n146 = n122 & n145 ;
  assign n147 = ~x1 & ~n146 ;
  assign n151 = ~x2 & n109 ;
  assign n152 = x2 & ~x6 ;
  assign n153 = ~n104 & n152 ;
  assign n154 = ~x7 & n108 ;
  assign n155 = ~n153 & ~n154 ;
  assign n156 = ~n151 & n155 ;
  assign n157 = ~x8 & ~n11 ;
  assign n158 = ~n156 & n157 ;
  assign n148 = x2 & ~x3 ;
  assign n149 = n148 ^ x4 ;
  assign n150 = n149 ^ n135 ;
  assign n159 = n158 ^ n150 ;
  assign n160 = n159 ^ n149 ;
  assign n161 = n150 ^ n148 ;
  assign n162 = n161 ^ n150 ;
  assign n163 = n162 ^ n160 ;
  assign n164 = ~n160 & ~n163 ;
  assign n165 = n164 ^ n158 ;
  assign n166 = n165 ^ n160 ;
  assign n167 = n158 ^ x7 ;
  assign n168 = n167 ^ n149 ;
  assign n169 = ~x7 & n168 ;
  assign n170 = n169 ^ x7 ;
  assign n171 = n170 ^ n158 ;
  assign n172 = n72 ^ x7 ;
  assign n173 = n167 & ~n172 ;
  assign n174 = n173 ^ n72 ;
  assign n175 = n174 ^ n149 ;
  assign n176 = n171 & n175 ;
  assign n177 = n176 ^ n149 ;
  assign n178 = n166 & n177 ;
  assign n179 = n178 ^ n164 ;
  assign n180 = n179 ^ n176 ;
  assign n181 = n180 ^ n160 ;
  assign n182 = n181 ^ x4 ;
  assign n183 = n182 ^ n158 ;
  assign n184 = ~n147 & n183 ;
  assign n185 = n107 & n184 ;
  assign n186 = n185 ^ n70 ;
  assign n187 = n186 ^ n69 ;
  assign n188 = n70 ^ n68 ;
  assign n189 = n188 ^ n185 ;
  assign n190 = n189 ^ n187 ;
  assign n191 = ~n187 & n190 ;
  assign n193 = n192 ^ n191 ;
  assign n194 = n193 ^ n187 ;
  assign n195 = ~n10 & n93 ;
  assign n196 = n84 & ~n195 ;
  assign n197 = x6 & ~n80 ;
  assign n198 = n197 ^ x8 ;
  assign n199 = n198 ^ n197 ;
  assign n200 = n197 ^ x2 ;
  assign n201 = n200 ^ n197 ;
  assign n202 = ~n199 & n201 ;
  assign n203 = n202 ^ n197 ;
  assign n204 = n11 & n203 ;
  assign n205 = n204 ^ n197 ;
  assign n206 = x3 & n205 ;
  assign n207 = n134 ^ x3 ;
  assign n208 = n207 ^ n134 ;
  assign n209 = n134 ^ n34 ;
  assign n210 = ~n208 & n209 ;
  assign n211 = n210 ^ n134 ;
  assign n212 = ~x2 & n211 ;
  assign n213 = ~n206 & ~n212 ;
  assign n214 = ~n196 & n213 ;
  assign n215 = ~x4 & ~n214 ;
  assign n216 = ~x6 & n15 ;
  assign n217 = ~x2 & n216 ;
  assign n218 = ~n141 & ~n151 ;
  assign n219 = n218 ^ x3 ;
  assign n220 = n219 ^ n218 ;
  assign n221 = x4 & n34 ;
  assign n222 = x2 & n72 ;
  assign n223 = ~n221 & ~n222 ;
  assign n224 = n223 ^ n218 ;
  assign n225 = n220 & n224 ;
  assign n226 = n225 ^ n218 ;
  assign n227 = x7 & ~n226 ;
  assign n228 = ~n217 & ~n227 ;
  assign n229 = ~n215 & n228 ;
  assign n230 = n81 ^ n80 ;
  assign n231 = x4 & ~n148 ;
  assign n232 = n231 ^ x6 ;
  assign n233 = n232 ^ n231 ;
  assign n234 = n231 ^ x2 ;
  assign n235 = ~n233 & ~n234 ;
  assign n236 = n235 ^ n231 ;
  assign n237 = n236 ^ n81 ;
  assign n238 = ~n230 & ~n237 ;
  assign n239 = n238 ^ n235 ;
  assign n240 = n239 ^ n231 ;
  assign n241 = n240 ^ n80 ;
  assign n242 = ~n81 & n241 ;
  assign n243 = n242 ^ n81 ;
  assign n244 = n229 & n243 ;
  assign n245 = n244 ^ n69 ;
  assign n246 = n191 ^ n187 ;
  assign n247 = ~n245 & ~n246 ;
  assign n248 = n247 ^ n69 ;
  assign n249 = n194 & ~n248 ;
  assign n250 = n249 ^ n69 ;
  assign n251 = n250 ^ x0 ;
  assign n252 = n251 ^ n69 ;
  assign y0 = ~n252 ;
endmodule
