module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 ;
  assign n11 = x2 & x6 ;
  assign n13 = x7 & x8 ;
  assign n12 = x5 ^ x3 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n11 & ~n14 ;
  assign n16 = n15 ^ n11 ;
  assign n17 = x9 ^ x3 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = ~n12 & n18 ;
  assign n20 = n19 ^ n12 ;
  assign n21 = n20 ^ n13 ;
  assign n22 = n16 & ~n21 ;
  assign n25 = ~x6 & ~x7 ;
  assign n26 = ~x8 & x9 ;
  assign n27 = n25 & n26 ;
  assign n28 = ~x2 & x5 ;
  assign n29 = n27 & n28 ;
  assign n32 = n29 ^ x2 ;
  assign n33 = n32 ^ n29 ;
  assign n23 = ~x8 & ~x9 ;
  assign n24 = x6 & n23 ;
  assign n30 = n29 ^ n24 ;
  assign n31 = n30 ^ n29 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = x5 & x7 ;
  assign n36 = n35 ^ n29 ;
  assign n37 = n36 ^ n29 ;
  assign n38 = n37 ^ n31 ;
  assign n39 = n31 & n38 ;
  assign n40 = n39 ^ n31 ;
  assign n41 = ~n34 & n40 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = n42 ^ n29 ;
  assign n44 = n43 ^ n31 ;
  assign n45 = ~x3 & n44 ;
  assign n46 = n45 ^ n29 ;
  assign n47 = ~n22 & ~n46 ;
  assign n48 = ~x4 & ~n47 ;
  assign n49 = x7 & n26 ;
  assign n50 = x2 & ~x6 ;
  assign n51 = n49 & n50 ;
  assign n52 = x4 & ~x5 ;
  assign n53 = x3 & n52 ;
  assign n54 = n51 & n53 ;
  assign n55 = ~n48 & ~n54 ;
  assign n56 = ~x0 & ~n55 ;
  assign n57 = x2 & x5 ;
  assign n58 = ~x3 & x4 ;
  assign n59 = ~x7 & x9 ;
  assign n60 = x0 & ~x6 ;
  assign n61 = n59 & n60 ;
  assign n62 = n58 & n61 ;
  assign n63 = n57 & n62 ;
  assign n64 = ~x8 & n63 ;
  assign n65 = n64 ^ n56 ;
  assign n66 = ~x5 & n23 ;
  assign n67 = ~x4 & n66 ;
  assign n68 = ~x6 & x7 ;
  assign n69 = ~x0 & ~x3 ;
  assign n70 = n68 & n69 ;
  assign n71 = n67 & n70 ;
  assign n72 = x5 & x6 ;
  assign n73 = ~x4 & n72 ;
  assign n74 = ~x6 & x9 ;
  assign n75 = n52 & n74 ;
  assign n76 = ~n73 & ~n75 ;
  assign n77 = x3 & ~x7 ;
  assign n78 = x8 & n77 ;
  assign n79 = x0 & n78 ;
  assign n80 = ~n76 & n79 ;
  assign n81 = ~n71 & ~n80 ;
  assign n177 = x8 & x9 ;
  assign n176 = ~x5 & n26 ;
  assign n178 = n177 ^ n176 ;
  assign n179 = ~x4 & n178 ;
  assign n180 = n179 ^ n177 ;
  assign n181 = n60 & n180 ;
  assign n182 = x5 & x8 ;
  assign n183 = x6 & ~n182 ;
  assign n184 = n183 ^ n66 ;
  assign n185 = n183 ^ x4 ;
  assign n186 = n185 ^ x4 ;
  assign n87 = x4 & x5 ;
  assign n187 = x4 & n177 ;
  assign n188 = ~n87 & ~n187 ;
  assign n189 = n188 ^ x4 ;
  assign n190 = n186 & ~n189 ;
  assign n191 = n190 ^ x4 ;
  assign n192 = n184 & n191 ;
  assign n193 = n192 ^ n66 ;
  assign n194 = n193 ^ x0 ;
  assign n195 = n194 ^ n193 ;
  assign n196 = x9 & n73 ;
  assign n197 = n196 ^ n193 ;
  assign n198 = n195 & n197 ;
  assign n199 = n198 ^ n193 ;
  assign n200 = ~n181 & ~n199 ;
  assign n201 = n77 & ~n200 ;
  assign n202 = x4 & x7 ;
  assign n203 = n66 & n202 ;
  assign n204 = n69 & n203 ;
  assign n205 = ~n201 & ~n204 ;
  assign n82 = x6 & x7 ;
  assign n83 = ~n25 & ~n82 ;
  assign n84 = x4 & ~x6 ;
  assign n85 = ~x5 & ~n84 ;
  assign n86 = ~n83 & n85 ;
  assign n88 = x0 & ~n87 ;
  assign n89 = ~x8 & ~n88 ;
  assign n90 = ~n86 & n89 ;
  assign n91 = ~x4 & ~x7 ;
  assign n92 = ~x3 & ~n91 ;
  assign n93 = ~n68 & ~n92 ;
  assign n94 = x5 & ~n93 ;
  assign n95 = x6 & ~x7 ;
  assign n96 = x3 & n95 ;
  assign n97 = ~n53 & ~n96 ;
  assign n98 = x6 & ~x9 ;
  assign n99 = ~x4 & ~n98 ;
  assign n100 = ~n25 & ~n99 ;
  assign n101 = n97 & ~n100 ;
  assign n102 = ~n94 & n101 ;
  assign n103 = n90 & n102 ;
  assign n104 = ~n74 & n103 ;
  assign n122 = ~x5 & x8 ;
  assign n123 = x3 & ~x4 ;
  assign n124 = n122 & n123 ;
  assign n125 = ~x7 & ~x8 ;
  assign n126 = x5 & n125 ;
  assign n127 = ~x3 & n126 ;
  assign n128 = ~n124 & ~n127 ;
  assign n105 = x4 ^ x3 ;
  assign n106 = ~x7 & n66 ;
  assign n107 = x5 & ~x9 ;
  assign n108 = n13 & n107 ;
  assign n109 = ~n106 & ~n108 ;
  assign n110 = n109 ^ x4 ;
  assign n111 = n110 ^ n109 ;
  assign n112 = n111 ^ n105 ;
  assign n113 = ~n49 & ~n107 ;
  assign n114 = n113 ^ n35 ;
  assign n115 = ~n113 & n114 ;
  assign n116 = n115 ^ n109 ;
  assign n117 = n116 ^ n113 ;
  assign n118 = ~n112 & n117 ;
  assign n119 = n118 ^ n115 ;
  assign n120 = n119 ^ n113 ;
  assign n121 = n105 & ~n120 ;
  assign n129 = n128 ^ n121 ;
  assign n130 = n129 ^ n121 ;
  assign n131 = n121 ^ x9 ;
  assign n132 = n131 ^ n121 ;
  assign n133 = ~n130 & n132 ;
  assign n134 = n133 ^ n121 ;
  assign n135 = ~x6 & n134 ;
  assign n136 = n135 ^ n121 ;
  assign n137 = n136 ^ x0 ;
  assign n138 = n137 ^ n136 ;
  assign n139 = n138 ^ n104 ;
  assign n140 = x7 & n98 ;
  assign n141 = n140 ^ x6 ;
  assign n142 = n141 ^ n140 ;
  assign n143 = n140 ^ n59 ;
  assign n144 = n143 ^ n140 ;
  assign n145 = n142 & n144 ;
  assign n146 = n145 ^ n140 ;
  assign n147 = ~x5 & n146 ;
  assign n148 = n147 ^ n140 ;
  assign n151 = n148 ^ x6 ;
  assign n152 = n151 ^ n148 ;
  assign n149 = n148 ^ x8 ;
  assign n150 = n149 ^ n148 ;
  assign n153 = n152 ^ n150 ;
  assign n154 = ~x5 & x9 ;
  assign n155 = ~n35 & ~n154 ;
  assign n156 = n155 ^ n148 ;
  assign n157 = n156 ^ n148 ;
  assign n158 = n157 ^ n152 ;
  assign n159 = ~n152 & n158 ;
  assign n160 = n159 ^ n152 ;
  assign n161 = ~n153 & ~n160 ;
  assign n162 = n161 ^ n159 ;
  assign n163 = n162 ^ n148 ;
  assign n164 = n163 ^ n152 ;
  assign n165 = x4 & ~n164 ;
  assign n166 = n165 ^ n148 ;
  assign n167 = n166 ^ x3 ;
  assign n168 = n166 & ~n167 ;
  assign n169 = n168 ^ n136 ;
  assign n170 = n169 ^ n166 ;
  assign n171 = n139 & n170 ;
  assign n172 = n171 ^ n168 ;
  assign n173 = n172 ^ n166 ;
  assign n174 = ~n104 & n173 ;
  assign n175 = n174 ^ n104 ;
  assign n206 = n205 ^ n175 ;
  assign n207 = n206 ^ n175 ;
  assign n208 = x0 & ~x3 ;
  assign n209 = ~n83 & n122 ;
  assign n210 = ~x4 & ~n209 ;
  assign n211 = ~x8 & ~n25 ;
  assign n212 = x5 & ~n82 ;
  assign n213 = ~n211 & ~n212 ;
  assign n214 = ~x9 & n213 ;
  assign n215 = n210 & n214 ;
  assign n216 = n49 & n73 ;
  assign n217 = ~n215 & ~n216 ;
  assign n218 = ~x6 & n182 ;
  assign n219 = ~x5 & x6 ;
  assign n220 = ~x8 & n219 ;
  assign n221 = ~n218 & ~n220 ;
  assign n222 = x9 & ~n221 ;
  assign n223 = x7 ^ x4 ;
  assign n224 = n222 & ~n223 ;
  assign n225 = n217 & ~n224 ;
  assign n226 = n208 & ~n225 ;
  assign n227 = ~x0 & ~x8 ;
  assign n228 = x5 & ~n227 ;
  assign n229 = ~n26 & ~n228 ;
  assign n230 = x0 & ~n23 ;
  assign n231 = x3 & x7 ;
  assign n232 = n84 & n231 ;
  assign n233 = ~n230 & n232 ;
  assign n234 = ~n229 & n233 ;
  assign n235 = ~n226 & ~n234 ;
  assign n236 = n235 ^ n175 ;
  assign n237 = n236 ^ n175 ;
  assign n238 = n207 & n237 ;
  assign n239 = n238 ^ n175 ;
  assign n240 = x2 & ~n239 ;
  assign n241 = n240 ^ n175 ;
  assign n242 = n81 & ~n241 ;
  assign n243 = n242 ^ x1 ;
  assign n244 = n243 ^ n242 ;
  assign n245 = ~x2 & ~x3 ;
  assign n246 = ~x5 & ~x6 ;
  assign n247 = ~x0 & ~n246 ;
  assign n248 = n83 & ~n247 ;
  assign n249 = n248 ^ x0 ;
  assign n250 = n249 ^ n248 ;
  assign n251 = n248 ^ n82 ;
  assign n252 = n251 ^ n248 ;
  assign n253 = ~n250 & n252 ;
  assign n254 = n253 ^ n248 ;
  assign n255 = x9 & n254 ;
  assign n256 = n255 ^ n248 ;
  assign n257 = x8 & n256 ;
  assign n258 = ~x6 & n106 ;
  assign n259 = ~n257 & ~n258 ;
  assign n260 = n245 & ~n259 ;
  assign n261 = n29 & ~n208 ;
  assign n285 = ~x7 & ~x9 ;
  assign n286 = x3 & n26 ;
  assign n287 = ~n285 & ~n286 ;
  assign n288 = x6 & ~n77 ;
  assign n289 = ~n287 & n288 ;
  assign n290 = ~n27 & ~n289 ;
  assign n291 = ~x0 & ~n290 ;
  assign n292 = n177 & n208 ;
  assign n293 = n95 & n292 ;
  assign n294 = ~n291 & ~n293 ;
  assign n262 = n13 ^ x0 ;
  assign n263 = n262 ^ x3 ;
  assign n270 = n263 ^ n262 ;
  assign n264 = n263 ^ n77 ;
  assign n265 = n264 ^ n262 ;
  assign n266 = n263 ^ n13 ;
  assign n267 = n266 ^ n77 ;
  assign n268 = n267 ^ n265 ;
  assign n269 = ~n265 & ~n268 ;
  assign n271 = n270 ^ n269 ;
  assign n272 = n271 ^ n265 ;
  assign n273 = n262 ^ x8 ;
  assign n274 = n269 ^ n265 ;
  assign n275 = n273 & ~n274 ;
  assign n276 = n275 ^ n262 ;
  assign n277 = ~n272 & n276 ;
  assign n278 = n277 ^ n262 ;
  assign n279 = n278 ^ x0 ;
  assign n280 = n279 ^ n262 ;
  assign n281 = ~x9 & n280 ;
  assign n282 = n59 & n227 ;
  assign n283 = x6 & ~n282 ;
  assign n284 = ~n281 & n283 ;
  assign n295 = n294 ^ n284 ;
  assign n296 = n295 ^ n294 ;
  assign n297 = x9 ^ x7 ;
  assign n298 = n227 & ~n297 ;
  assign n299 = ~n231 & n298 ;
  assign n300 = ~x6 & ~n299 ;
  assign n301 = x7 & n292 ;
  assign n302 = n300 & ~n301 ;
  assign n303 = n302 ^ n294 ;
  assign n304 = n303 ^ n294 ;
  assign n305 = ~n296 & ~n304 ;
  assign n306 = n305 ^ n294 ;
  assign n307 = x5 & ~n306 ;
  assign n308 = n307 ^ n294 ;
  assign n309 = x2 & ~n308 ;
  assign n310 = ~n261 & ~n309 ;
  assign n311 = ~n260 & n310 ;
  assign n312 = ~x4 & ~n311 ;
  assign n313 = n50 & n59 ;
  assign n314 = ~x3 & n140 ;
  assign n315 = ~n313 & ~n314 ;
  assign n316 = n122 & ~n315 ;
  assign n317 = ~x6 & n177 ;
  assign n318 = n23 & n219 ;
  assign n319 = ~n317 & ~n318 ;
  assign n320 = n231 & ~n319 ;
  assign n321 = x6 & x8 ;
  assign n322 = ~x2 & ~n321 ;
  assign n323 = n107 & ~n245 ;
  assign n324 = ~n322 & n323 ;
  assign n325 = ~x3 & ~x5 ;
  assign n326 = n27 & n325 ;
  assign n327 = ~n324 & ~n326 ;
  assign n328 = ~n320 & n327 ;
  assign n329 = ~x3 & ~x8 ;
  assign n330 = n68 & n329 ;
  assign n331 = ~n78 & ~n330 ;
  assign n332 = n107 & ~n331 ;
  assign n333 = x2 & ~n332 ;
  assign n334 = ~n328 & ~n333 ;
  assign n335 = n28 & ~n82 ;
  assign n336 = n286 & n335 ;
  assign n337 = ~x0 & ~n336 ;
  assign n338 = ~n334 & n337 ;
  assign n339 = ~n316 & n338 ;
  assign n340 = x4 & ~n339 ;
  assign n341 = n340 ^ x0 ;
  assign n342 = x3 & x5 ;
  assign n343 = x9 ^ x8 ;
  assign n344 = x8 ^ x7 ;
  assign n345 = n344 ^ n343 ;
  assign n346 = n11 ^ x9 ;
  assign n347 = n346 ^ n11 ;
  assign n348 = ~x2 & ~x6 ;
  assign n349 = n348 ^ n11 ;
  assign n350 = n347 & n349 ;
  assign n351 = n350 ^ n11 ;
  assign n352 = n351 ^ n343 ;
  assign n353 = n345 & ~n352 ;
  assign n354 = n353 ^ n350 ;
  assign n355 = n354 ^ n11 ;
  assign n356 = n355 ^ n344 ;
  assign n357 = ~n343 & ~n356 ;
  assign n358 = n357 ^ n343 ;
  assign n359 = n342 & ~n358 ;
  assign n360 = n359 ^ n340 ;
  assign n361 = n360 ^ n359 ;
  assign n362 = n361 ^ n341 ;
  assign n363 = x6 ^ x2 ;
  assign n364 = n363 ^ n343 ;
  assign n370 = n364 ^ x9 ;
  assign n371 = n370 ^ n364 ;
  assign n365 = n343 ^ x5 ;
  assign n366 = n365 ^ n364 ;
  assign n367 = n366 ^ n343 ;
  assign n368 = n367 ^ x2 ;
  assign n369 = n368 ^ n364 ;
  assign n372 = n371 ^ n369 ;
  assign n375 = n368 ^ x2 ;
  assign n373 = n343 ^ x2 ;
  assign n374 = n373 ^ n369 ;
  assign n376 = n375 ^ n374 ;
  assign n377 = ~n372 & n376 ;
  assign n378 = n377 ^ n368 ;
  assign n379 = n378 ^ n373 ;
  assign n380 = n379 ^ n375 ;
  assign n381 = n374 ^ n371 ;
  assign n382 = n378 & n381 ;
  assign n383 = n382 ^ n368 ;
  assign n384 = n383 ^ n369 ;
  assign n385 = n384 ^ n371 ;
  assign n386 = ~n380 & ~n385 ;
  assign n387 = n231 & n386 ;
  assign n388 = x8 & ~x9 ;
  assign n389 = n95 & n388 ;
  assign n390 = ~n51 & ~n389 ;
  assign n391 = n325 & ~n390 ;
  assign n392 = ~n387 & ~n391 ;
  assign n393 = x7 ^ x6 ;
  assign n394 = n388 ^ n13 ;
  assign n395 = n394 ^ n13 ;
  assign n396 = n13 ^ x7 ;
  assign n397 = n396 ^ n13 ;
  assign n398 = ~n395 & ~n397 ;
  assign n399 = n398 ^ n13 ;
  assign n400 = ~x6 & n399 ;
  assign n401 = n400 ^ n13 ;
  assign n402 = ~x3 & n401 ;
  assign n403 = n402 ^ n393 ;
  assign n404 = n26 ^ x6 ;
  assign n405 = n404 ^ n26 ;
  assign n406 = n388 ^ n26 ;
  assign n407 = ~n405 & n406 ;
  assign n408 = n407 ^ n26 ;
  assign n409 = n408 ^ n393 ;
  assign n410 = ~n403 & n409 ;
  assign n411 = n410 ^ n407 ;
  assign n412 = n411 ^ n26 ;
  assign n413 = n412 ^ n402 ;
  assign n414 = n393 & ~n413 ;
  assign n415 = n414 ^ n393 ;
  assign n416 = n415 ^ n402 ;
  assign n417 = n57 & n416 ;
  assign n418 = n218 & n285 ;
  assign n419 = n82 & n176 ;
  assign n420 = ~n418 & ~n419 ;
  assign n421 = n245 & ~n420 ;
  assign n422 = ~n24 & ~n317 ;
  assign n423 = n28 & ~n422 ;
  assign n424 = n77 & n423 ;
  assign n425 = ~n421 & ~n424 ;
  assign n426 = ~n417 & n425 ;
  assign n427 = n426 ^ n392 ;
  assign n428 = n392 & n427 ;
  assign n429 = n428 ^ n359 ;
  assign n430 = n429 ^ n392 ;
  assign n431 = ~n362 & n430 ;
  assign n432 = n431 ^ n428 ;
  assign n433 = n432 ^ n392 ;
  assign n434 = ~n341 & n433 ;
  assign n435 = n434 ^ n340 ;
  assign n436 = ~n312 & ~n435 ;
  assign n437 = n436 ^ n242 ;
  assign n438 = ~n244 & n437 ;
  assign n439 = n438 ^ n242 ;
  assign n440 = n439 ^ n56 ;
  assign n441 = n65 & ~n440 ;
  assign n442 = n441 ^ n438 ;
  assign n443 = n442 ^ n242 ;
  assign n444 = n443 ^ n64 ;
  assign n445 = ~n56 & ~n444 ;
  assign n446 = n445 ^ n56 ;
  assign y0 = n446 ;
endmodule
