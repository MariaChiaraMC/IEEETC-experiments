module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 ;
  assign n18 = ~x11 & ~x13 ;
  assign n24 = x15 & x16 ;
  assign n25 = x14 & n24 ;
  assign n19 = ~x15 & ~x16 ;
  assign n20 = x1 & x3 ;
  assign n21 = n19 & n20 ;
  assign n22 = ~x4 & x6 ;
  assign n23 = n21 & n22 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = n25 ^ x14 ;
  assign n29 = n28 ^ n25 ;
  assign n30 = n27 & ~n29 ;
  assign n31 = n30 ^ n25 ;
  assign n32 = ~x12 & n31 ;
  assign n33 = n32 ^ n25 ;
  assign n34 = n18 & n33 ;
  assign n35 = n25 ^ x13 ;
  assign n36 = ~x12 & ~x14 ;
  assign n37 = ~n24 & n36 ;
  assign n38 = n37 ^ x11 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = n37 ^ x12 ;
  assign n41 = ~n39 & n40 ;
  assign n42 = n41 ^ n37 ;
  assign n43 = n42 ^ n25 ;
  assign n44 = ~n35 & ~n43 ;
  assign n45 = n44 ^ n41 ;
  assign n46 = n45 ^ n37 ;
  assign n47 = n46 ^ x13 ;
  assign n48 = ~n25 & n47 ;
  assign n49 = n48 ^ n25 ;
  assign n50 = ~n34 & n49 ;
  assign n51 = ~x0 & ~n50 ;
  assign y0 = n51 ;
endmodule
