module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n10 = x7 ^ x3 ;
  assign n11 = n10 ^ x6 ;
  assign n13 = x4 & x8 ;
  assign n12 = ~x4 & ~x8 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = ~x3 & n14 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = ~n11 & ~n16 ;
  assign n18 = n17 ^ n15 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = n19 ^ x3 ;
  assign n21 = ~x6 & n20 ;
  assign n22 = x2 & ~n21 ;
  assign n23 = x3 & n14 ;
  assign n24 = n23 ^ n13 ;
  assign n25 = n11 & n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n26 ^ n13 ;
  assign n28 = n27 ^ x3 ;
  assign n29 = x6 & n28 ;
  assign n30 = ~n22 & ~n29 ;
  assign y0 = ~n30 ;
endmodule
