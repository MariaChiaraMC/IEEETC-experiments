module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 ;
  assign n9 = x4 & x7 ;
  assign n10 = ~x0 & n9 ;
  assign n11 = x6 ^ x3 ;
  assign n12 = n11 ^ x6 ;
  assign n13 = x6 ^ x2 ;
  assign n14 = ~n12 & n13 ;
  assign n15 = n14 ^ x6 ;
  assign n16 = x1 & ~x6 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = ~n15 & n17 ;
  assign n19 = n18 ^ n16 ;
  assign n20 = x5 & n19 ;
  assign n21 = n20 ^ x5 ;
  assign n22 = n10 & n21 ;
  assign y0 = n22 ;
endmodule
