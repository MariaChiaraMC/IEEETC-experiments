module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 ;
  assign n11 = x4 ^ x3 ;
  assign n12 = x5 ^ x4 ;
  assign n13 = ~n11 & n12 ;
  assign n14 = x0 & n13 ;
  assign n15 = ~x1 & n14 ;
  assign n7 = ~x4 & x5 ;
  assign n8 = ~x3 & n7 ;
  assign n9 = ~x0 & x1 ;
  assign n10 = n8 & n9 ;
  assign n16 = n15 ^ n10 ;
  assign n17 = n16 ^ n10 ;
  assign n18 = x4 & ~x5 ;
  assign n19 = n9 & n18 ;
  assign n20 = n19 ^ n10 ;
  assign n21 = n20 ^ n10 ;
  assign n22 = ~n17 & ~n21 ;
  assign n23 = n22 ^ n10 ;
  assign n24 = x2 & ~n23 ;
  assign n25 = n24 ^ n10 ;
  assign y0 = n25 ;
endmodule
