module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 ;
  assign n7 = ~x0 & ~x1 ;
  assign n8 = x5 ^ x4 ;
  assign n9 = n8 ^ x3 ;
  assign n10 = n8 ^ x5 ;
  assign n11 = x5 ^ x2 ;
  assign n12 = ~x5 & ~n11 ;
  assign n13 = n12 ^ x5 ;
  assign n14 = n10 & ~n13 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n15 ^ x5 ;
  assign n17 = n16 ^ x2 ;
  assign n18 = n9 & ~n17 ;
  assign n19 = n18 ^ n8 ;
  assign n20 = n7 & ~n19 ;
  assign y0 = n20 ;
endmodule
