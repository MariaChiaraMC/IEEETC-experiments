module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 ;
  assign n17 = x4 ^ x3 ;
  assign n18 = ~x9 & ~x10 ;
  assign n19 = ~x8 & n18 ;
  assign n20 = ~x7 & ~n19 ;
  assign n21 = ~x11 & ~x12 ;
  assign n22 = ~x14 & ~x15 ;
  assign n23 = ~x8 & n22 ;
  assign n24 = n23 ^ x13 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = x15 ^ x14 ;
  assign n27 = x9 & x10 ;
  assign n28 = n27 ^ x15 ;
  assign n29 = x14 ^ x8 ;
  assign n30 = n29 ^ x15 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = ~n27 & ~n31 ;
  assign n33 = n32 ^ n27 ;
  assign n34 = n28 & ~n33 ;
  assign n35 = n34 ^ n32 ;
  assign n36 = n35 ^ n27 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = ~n26 & ~n37 ;
  assign n39 = n38 ^ n30 ;
  assign n40 = n39 ^ n23 ;
  assign n41 = ~n25 & n40 ;
  assign n42 = n41 ^ n23 ;
  assign n43 = n21 & n42 ;
  assign n44 = n20 & ~n43 ;
  assign n45 = x1 & ~x2 ;
  assign n46 = x6 & n45 ;
  assign n47 = ~n44 & n46 ;
  assign n48 = ~x0 & n47 ;
  assign n49 = n48 ^ x5 ;
  assign n50 = n49 ^ n48 ;
  assign n51 = x0 & ~x1 ;
  assign n52 = n51 ^ n48 ;
  assign n53 = n50 & n52 ;
  assign n54 = n53 ^ n48 ;
  assign n55 = n54 ^ x4 ;
  assign n56 = n17 & ~n55 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = n57 ^ n48 ;
  assign n59 = n58 ^ x3 ;
  assign n60 = ~x4 & ~n59 ;
  assign n61 = n60 ^ x4 ;
  assign y0 = ~n61 ;
endmodule
