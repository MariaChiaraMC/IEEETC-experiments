module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 ;
  assign n11 = ~x2 & ~x3 ;
  assign n12 = x1 & n11 ;
  assign n13 = x5 & ~n12 ;
  assign n14 = x3 ^ x2 ;
  assign n15 = x3 ^ x1 ;
  assign n16 = n15 ^ x3 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = x7 ^ x6 ;
  assign n19 = x3 & n18 ;
  assign n20 = n19 ^ x7 ;
  assign n21 = n17 & n20 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ x7 ;
  assign n24 = n23 ^ x3 ;
  assign n25 = n14 & n24 ;
  assign n26 = n25 ^ x2 ;
  assign n27 = n13 & ~n26 ;
  assign n28 = x2 & ~x5 ;
  assign n29 = x3 & ~x7 ;
  assign n30 = n28 & n29 ;
  assign n31 = ~x7 & ~x8 ;
  assign n32 = ~x7 & ~x9 ;
  assign n33 = n11 & ~n32 ;
  assign n34 = ~n31 & n33 ;
  assign n35 = ~n30 & ~n34 ;
  assign n36 = ~x1 & x6 ;
  assign n37 = ~n35 & n36 ;
  assign n42 = x2 & x5 ;
  assign n38 = x6 & ~n31 ;
  assign n39 = ~x2 & ~x5 ;
  assign n40 = x1 & n39 ;
  assign n41 = ~n38 & n40 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = n43 ^ x3 ;
  assign n52 = n44 ^ n43 ;
  assign n45 = n44 ^ n41 ;
  assign n46 = n45 ^ n44 ;
  assign n47 = n46 ^ n43 ;
  assign n48 = n45 ^ x6 ;
  assign n49 = n48 ^ n45 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = n47 & n50 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n53 ^ n47 ;
  assign n55 = x7 & x8 ;
  assign n56 = n55 ^ n43 ;
  assign n57 = n51 ^ n47 ;
  assign n58 = n56 & n57 ;
  assign n59 = n58 ^ n43 ;
  assign n60 = ~n54 & n59 ;
  assign n61 = n60 ^ n43 ;
  assign n62 = n61 ^ n42 ;
  assign n63 = n62 ^ n43 ;
  assign n64 = ~x0 & n63 ;
  assign n65 = ~n37 & ~n64 ;
  assign n66 = ~n27 & n65 ;
  assign n67 = x4 & ~n66 ;
  assign n68 = x1 & x2 ;
  assign n69 = x6 & n28 ;
  assign n70 = ~n68 & ~n69 ;
  assign n71 = x5 & ~x6 ;
  assign n72 = x1 & n71 ;
  assign n73 = ~n31 & n72 ;
  assign n74 = n70 & ~n73 ;
  assign n75 = x3 & ~n74 ;
  assign n76 = x7 & x9 ;
  assign n77 = x1 & x3 ;
  assign n78 = ~n76 & n77 ;
  assign n79 = x2 & ~x6 ;
  assign n80 = ~n55 & n79 ;
  assign n81 = n78 & n80 ;
  assign n82 = x3 & ~x5 ;
  assign n83 = x8 ^ x1 ;
  assign n84 = n83 ^ x1 ;
  assign n85 = x6 ^ x1 ;
  assign n86 = n85 ^ x1 ;
  assign n87 = n84 & ~n86 ;
  assign n88 = n87 ^ x1 ;
  assign n89 = ~x2 & n88 ;
  assign n90 = n89 ^ x1 ;
  assign n91 = n82 & n90 ;
  assign n92 = ~x1 & ~x5 ;
  assign n93 = n92 ^ n14 ;
  assign n94 = x6 ^ x2 ;
  assign n95 = n94 ^ x6 ;
  assign n96 = n18 & ~n95 ;
  assign n97 = n96 ^ x6 ;
  assign n98 = n97 ^ n14 ;
  assign n99 = n93 & ~n98 ;
  assign n100 = n99 ^ n96 ;
  assign n101 = n100 ^ x6 ;
  assign n102 = n101 ^ n92 ;
  assign n103 = n14 & ~n102 ;
  assign n104 = n103 ^ n14 ;
  assign n105 = ~n91 & ~n104 ;
  assign n106 = ~n81 & n105 ;
  assign n107 = n29 ^ x5 ;
  assign n108 = n107 ^ x1 ;
  assign n115 = n108 ^ n107 ;
  assign n110 = x3 & ~x6 ;
  assign n109 = n108 ^ n29 ;
  assign n111 = n110 ^ n109 ;
  assign n112 = n110 ^ n108 ;
  assign n113 = n112 ^ n107 ;
  assign n114 = ~n111 & n113 ;
  assign n116 = n115 ^ n114 ;
  assign n117 = ~x6 & ~x7 ;
  assign n118 = ~x3 & ~n117 ;
  assign n119 = n118 ^ n108 ;
  assign n120 = ~n115 & ~n119 ;
  assign n121 = n120 ^ n118 ;
  assign n122 = ~n116 & n121 ;
  assign n123 = n122 ^ n114 ;
  assign n124 = n123 ^ n108 ;
  assign n125 = n124 ^ x5 ;
  assign n126 = n125 ^ n107 ;
  assign n127 = ~x2 & ~n126 ;
  assign n128 = x5 ^ x1 ;
  assign n129 = x6 & n55 ;
  assign n130 = n129 ^ x5 ;
  assign n131 = n128 & n130 ;
  assign n132 = n131 ^ x5 ;
  assign n133 = x3 & x5 ;
  assign n134 = n133 ^ x2 ;
  assign n135 = n132 & n134 ;
  assign n136 = n135 ^ n133 ;
  assign n137 = x2 & n136 ;
  assign n138 = n137 ^ x2 ;
  assign n139 = n82 ^ x9 ;
  assign n140 = n139 ^ n82 ;
  assign n141 = ~x6 & n31 ;
  assign n142 = ~x1 & x3 ;
  assign n143 = n141 & n142 ;
  assign n144 = ~n28 & ~n143 ;
  assign n145 = n144 ^ n82 ;
  assign n146 = ~n140 & ~n145 ;
  assign n147 = n146 ^ n82 ;
  assign n148 = n82 & ~n117 ;
  assign n149 = n148 ^ n138 ;
  assign n150 = n147 & ~n149 ;
  assign n151 = n150 ^ n148 ;
  assign n152 = ~n138 & n151 ;
  assign n153 = n152 ^ n138 ;
  assign n154 = ~n127 & ~n153 ;
  assign n155 = n106 & n154 ;
  assign n156 = ~x4 & ~n155 ;
  assign n157 = ~n75 & ~n156 ;
  assign n158 = n157 ^ x0 ;
  assign n159 = n158 ^ n157 ;
  assign n160 = ~x3 & ~n141 ;
  assign n161 = ~n110 & ~n160 ;
  assign n162 = n39 & ~n161 ;
  assign n163 = ~x6 & ~n55 ;
  assign n164 = n42 & ~n163 ;
  assign n165 = n142 & n164 ;
  assign n166 = ~x4 & ~n165 ;
  assign n167 = n106 & n166 ;
  assign n168 = ~n162 & n167 ;
  assign n169 = n141 ^ x5 ;
  assign n170 = n169 ^ x2 ;
  assign n171 = ~x1 & ~x9 ;
  assign n172 = n171 ^ n77 ;
  assign n173 = x5 & n172 ;
  assign n174 = n173 ^ n77 ;
  assign n175 = n170 & n174 ;
  assign n176 = n175 ^ n173 ;
  assign n177 = n176 ^ n77 ;
  assign n178 = n177 ^ x5 ;
  assign n179 = ~x2 & n178 ;
  assign n180 = n179 ^ x4 ;
  assign n181 = x7 & n68 ;
  assign n182 = ~n69 & ~n181 ;
  assign n183 = x9 & n129 ;
  assign n184 = n183 ^ x5 ;
  assign n185 = n182 & ~n184 ;
  assign n186 = n185 ^ x3 ;
  assign n187 = n186 ^ n185 ;
  assign n188 = n79 & n92 ;
  assign n189 = n188 ^ n185 ;
  assign n190 = n187 & ~n189 ;
  assign n191 = n190 ^ n185 ;
  assign n192 = n191 ^ n179 ;
  assign n193 = ~n180 & ~n192 ;
  assign n194 = n193 ^ n190 ;
  assign n195 = n194 ^ n185 ;
  assign n196 = n195 ^ x4 ;
  assign n197 = ~n179 & n196 ;
  assign n198 = n197 ^ n179 ;
  assign n199 = ~n168 & n198 ;
  assign n200 = x6 & ~n55 ;
  assign n201 = ~x3 & n92 ;
  assign n202 = n200 & n201 ;
  assign n203 = x1 & ~n71 ;
  assign n204 = n11 & ~n203 ;
  assign n205 = ~n202 & ~n204 ;
  assign n206 = ~n199 & n205 ;
  assign n207 = n206 ^ n157 ;
  assign n208 = n159 & n207 ;
  assign n209 = n208 ^ n157 ;
  assign n210 = ~n67 & n209 ;
  assign y0 = ~n210 ;
endmodule
