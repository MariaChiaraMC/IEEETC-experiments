module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 ;
  assign n9 = ~x2 & x3 ;
  assign n10 = x4 & ~x6 ;
  assign n11 = ~x0 & ~x5 ;
  assign n12 = x7 & n11 ;
  assign n13 = n10 & n12 ;
  assign n14 = n9 & n13 ;
  assign n52 = x4 ^ x3 ;
  assign n53 = n52 ^ x6 ;
  assign n37 = x0 & ~x7 ;
  assign n54 = n53 ^ n37 ;
  assign n55 = x6 ^ x4 ;
  assign n56 = n55 ^ x6 ;
  assign n57 = x6 ^ x2 ;
  assign n58 = n56 & ~n57 ;
  assign n59 = n58 ^ x6 ;
  assign n60 = n59 ^ n53 ;
  assign n61 = ~n54 & ~n60 ;
  assign n62 = n61 ^ n58 ;
  assign n63 = n62 ^ x6 ;
  assign n64 = n63 ^ n37 ;
  assign n65 = ~n53 & n64 ;
  assign n66 = n65 ^ n53 ;
  assign n67 = x5 & n66 ;
  assign n68 = x2 & ~x3 ;
  assign n69 = n10 & n37 ;
  assign n70 = ~x0 & x6 ;
  assign n71 = x4 & n70 ;
  assign n72 = ~n69 & ~n71 ;
  assign n73 = n68 & ~n72 ;
  assign n74 = x7 & ~n73 ;
  assign n15 = x2 & x3 ;
  assign n75 = ~x0 & ~x4 ;
  assign n76 = ~n10 & ~n75 ;
  assign n77 = n15 & ~n76 ;
  assign n78 = n77 ^ n73 ;
  assign n79 = x4 & x6 ;
  assign n80 = ~x2 & ~x3 ;
  assign n81 = x6 ^ x0 ;
  assign n82 = n80 & n81 ;
  assign n83 = ~n79 & n82 ;
  assign n84 = n83 ^ n74 ;
  assign n85 = n78 & n84 ;
  assign n86 = n85 ^ n83 ;
  assign n87 = n74 & n86 ;
  assign n88 = n87 ^ n73 ;
  assign n89 = n67 & ~n88 ;
  assign n90 = ~n9 & ~n68 ;
  assign n91 = ~x4 & ~x7 ;
  assign n32 = ~x2 & x6 ;
  assign n92 = x0 & ~n32 ;
  assign n93 = n91 & ~n92 ;
  assign n94 = ~n90 & n93 ;
  assign n95 = n69 & n90 ;
  assign n96 = ~x5 & ~n95 ;
  assign n97 = x4 ^ x0 ;
  assign n21 = ~x6 & x7 ;
  assign n98 = n97 ^ n21 ;
  assign n99 = x2 ^ x0 ;
  assign n100 = n99 ^ x2 ;
  assign n101 = n15 ^ x2 ;
  assign n102 = n100 & ~n101 ;
  assign n103 = n102 ^ x2 ;
  assign n104 = n103 ^ n97 ;
  assign n105 = n98 & ~n104 ;
  assign n106 = n105 ^ n102 ;
  assign n107 = n106 ^ x2 ;
  assign n108 = n107 ^ n21 ;
  assign n109 = n97 & ~n108 ;
  assign n110 = n109 ^ n97 ;
  assign n111 = n96 & ~n110 ;
  assign n112 = ~n94 & n111 ;
  assign n113 = ~n89 & ~n112 ;
  assign n16 = x5 ^ x0 ;
  assign n22 = n21 ^ x0 ;
  assign n23 = ~x0 & n22 ;
  assign n17 = x3 & x6 ;
  assign n18 = ~x2 & n17 ;
  assign n19 = x7 & n18 ;
  assign n26 = n23 ^ n19 ;
  assign n20 = n19 ^ n16 ;
  assign n24 = n23 ^ x0 ;
  assign n25 = ~n20 & ~n24 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = ~n16 & n27 ;
  assign n29 = n28 ^ n23 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = ~n15 & n30 ;
  assign n33 = ~x3 & ~x5 ;
  assign n34 = ~x0 & ~x7 ;
  assign n35 = n33 & n34 ;
  assign n36 = n32 & n35 ;
  assign n39 = x3 & x5 ;
  assign n40 = ~n33 & ~n39 ;
  assign n38 = ~x2 & ~x6 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = ~x3 & ~x6 ;
  assign n44 = x2 & ~n43 ;
  assign n45 = n44 ^ n38 ;
  assign n46 = n42 & n45 ;
  assign n47 = n46 ^ n38 ;
  assign n48 = n37 & n47 ;
  assign n49 = ~n36 & ~n48 ;
  assign n50 = ~n31 & n49 ;
  assign n51 = ~x4 & ~n50 ;
  assign n114 = n113 ^ n51 ;
  assign n115 = n114 ^ n113 ;
  assign n116 = ~n33 & ~n79 ;
  assign n117 = ~n12 & ~n116 ;
  assign n118 = n90 ^ x4 ;
  assign n119 = n118 ^ n90 ;
  assign n120 = n90 ^ x2 ;
  assign n121 = n120 ^ n90 ;
  assign n122 = n119 & ~n121 ;
  assign n123 = n122 ^ n90 ;
  assign n124 = ~x6 & ~n123 ;
  assign n125 = n124 ^ n90 ;
  assign n126 = n117 & ~n125 ;
  assign n127 = n39 ^ x7 ;
  assign n128 = n127 ^ n39 ;
  assign n129 = ~x0 & x5 ;
  assign n130 = ~x0 & ~x6 ;
  assign n131 = ~n39 & ~n130 ;
  assign n132 = ~n129 & ~n131 ;
  assign n133 = n132 ^ n39 ;
  assign n134 = ~n128 & ~n133 ;
  assign n135 = n134 ^ n39 ;
  assign n136 = n126 & ~n135 ;
  assign n137 = n136 ^ n113 ;
  assign n138 = n137 ^ n113 ;
  assign n139 = ~n115 & ~n138 ;
  assign n140 = n139 ^ n113 ;
  assign n141 = x1 & ~n140 ;
  assign n142 = n141 ^ n113 ;
  assign n143 = ~n14 & ~n142 ;
  assign y0 = ~n143 ;
endmodule
