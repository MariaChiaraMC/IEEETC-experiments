module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 ;
  assign n16 = x7 & ~x9 ;
  assign n17 = x6 & n16 ;
  assign n18 = x3 & ~x4 ;
  assign n19 = n17 & n18 ;
  assign n20 = x2 & ~x10 ;
  assign n21 = n19 & n20 ;
  assign n22 = x2 & x5 ;
  assign n23 = ~x3 & ~x4 ;
  assign n24 = ~x1 & x2 ;
  assign n25 = ~x10 & ~n24 ;
  assign n26 = n23 & n25 ;
  assign n27 = n17 & n26 ;
  assign n28 = ~n22 & ~n27 ;
  assign n29 = ~n21 & n28 ;
  assign n30 = x13 & x14 ;
  assign n31 = ~x0 & x2 ;
  assign n32 = ~x1 & n31 ;
  assign n33 = ~x6 & x9 ;
  assign n34 = ~x3 & x4 ;
  assign n35 = x10 & n34 ;
  assign n36 = n33 & n35 ;
  assign n37 = n32 & n36 ;
  assign n38 = n37 ^ x5 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = n37 ^ x0 ;
  assign n41 = ~n39 & n40 ;
  assign n42 = n41 ^ n37 ;
  assign n43 = ~n30 & n42 ;
  assign n44 = ~n29 & n43 ;
  assign n45 = ~x13 & ~x14 ;
  assign n46 = n31 & n45 ;
  assign n49 = x1 & x4 ;
  assign n50 = x9 & n49 ;
  assign n47 = ~x1 & ~x4 ;
  assign n48 = n17 & n47 ;
  assign n51 = n50 ^ n48 ;
  assign n52 = n51 ^ x5 ;
  assign n61 = n52 ^ n51 ;
  assign n53 = x6 & x10 ;
  assign n54 = ~x7 & ~n53 ;
  assign n55 = n54 ^ n52 ;
  assign n56 = n55 ^ n51 ;
  assign n57 = n52 ^ n48 ;
  assign n58 = n57 ^ n54 ;
  assign n59 = n58 ^ n56 ;
  assign n60 = ~n56 & ~n59 ;
  assign n62 = n61 ^ n60 ;
  assign n63 = n62 ^ n56 ;
  assign n64 = x7 & x10 ;
  assign n65 = x6 & ~n64 ;
  assign n66 = n65 ^ n51 ;
  assign n67 = n60 ^ n56 ;
  assign n68 = n66 & ~n67 ;
  assign n69 = n68 ^ n51 ;
  assign n70 = ~n63 & n69 ;
  assign n71 = n70 ^ n51 ;
  assign n72 = n71 ^ n50 ;
  assign n73 = n72 ^ n51 ;
  assign n74 = n46 & n73 ;
  assign n75 = x3 & n74 ;
  assign n76 = ~n44 & ~n75 ;
  assign n77 = ~x8 & ~n76 ;
  assign n98 = ~x1 & x7 ;
  assign n99 = n31 & n98 ;
  assign n100 = ~x9 & x10 ;
  assign n101 = x3 & x4 ;
  assign n102 = n100 & n101 ;
  assign n103 = n99 & n102 ;
  assign n105 = n103 ^ x5 ;
  assign n114 = n105 ^ n103 ;
  assign n78 = ~x0 & ~x1 ;
  assign n79 = ~x2 & n78 ;
  assign n80 = ~x7 & x10 ;
  assign n81 = n79 & n80 ;
  assign n82 = ~x3 & ~x10 ;
  assign n83 = x0 & x1 ;
  assign n84 = n83 ^ n82 ;
  assign n85 = n22 ^ x7 ;
  assign n86 = n85 ^ n22 ;
  assign n87 = n22 ^ x5 ;
  assign n88 = ~n86 & ~n87 ;
  assign n89 = n88 ^ n22 ;
  assign n90 = n89 ^ n82 ;
  assign n91 = n84 & n90 ;
  assign n92 = n91 ^ n88 ;
  assign n93 = n92 ^ n22 ;
  assign n94 = n93 ^ n83 ;
  assign n95 = n82 & n94 ;
  assign n96 = n95 ^ n82 ;
  assign n97 = ~n81 & ~n96 ;
  assign n104 = n103 ^ n97 ;
  assign n106 = n105 ^ n104 ;
  assign n107 = n106 ^ n105 ;
  assign n108 = n107 ^ n103 ;
  assign n109 = ~x4 & x9 ;
  assign n110 = n109 ^ n106 ;
  assign n111 = n110 ^ n106 ;
  assign n112 = n111 ^ n108 ;
  assign n113 = ~n108 & ~n112 ;
  assign n115 = n114 ^ n113 ;
  assign n116 = n115 ^ n108 ;
  assign n117 = n103 ^ x3 ;
  assign n118 = n113 ^ n108 ;
  assign n119 = n117 & ~n118 ;
  assign n120 = n119 ^ n103 ;
  assign n121 = ~n116 & ~n120 ;
  assign n122 = n121 ^ n103 ;
  assign n123 = n122 ^ x5 ;
  assign n124 = n123 ^ n103 ;
  assign n125 = x8 & n124 ;
  assign n126 = ~x8 & ~x9 ;
  assign n127 = ~x10 & n126 ;
  assign n128 = x5 & ~x7 ;
  assign n129 = n34 & n128 ;
  assign n130 = n127 & n129 ;
  assign n131 = n32 & n130 ;
  assign n132 = ~n125 & ~n131 ;
  assign n136 = n132 ^ x8 ;
  assign n137 = n136 ^ n132 ;
  assign n133 = x3 & ~x5 ;
  assign n134 = n133 ^ n132 ;
  assign n135 = n134 ^ n132 ;
  assign n138 = n137 ^ n135 ;
  assign n139 = ~x4 & n64 ;
  assign n140 = n32 & n139 ;
  assign n141 = n140 ^ n132 ;
  assign n142 = n141 ^ n132 ;
  assign n143 = n142 ^ n137 ;
  assign n144 = ~n137 & ~n143 ;
  assign n145 = n144 ^ n137 ;
  assign n146 = ~n138 & ~n145 ;
  assign n147 = n146 ^ n144 ;
  assign n148 = n147 ^ n132 ;
  assign n149 = n148 ^ n137 ;
  assign n150 = ~x6 & n149 ;
  assign n151 = n150 ^ n132 ;
  assign n152 = ~n30 & ~n151 ;
  assign n165 = ~x8 & x9 ;
  assign n166 = n49 & n165 ;
  assign n153 = n47 ^ x9 ;
  assign n154 = n153 ^ x8 ;
  assign n155 = n154 ^ n47 ;
  assign n156 = n155 ^ x6 ;
  assign n157 = n49 ^ x8 ;
  assign n158 = n49 & ~n157 ;
  assign n159 = n158 ^ n47 ;
  assign n160 = n159 ^ n49 ;
  assign n161 = n156 & n160 ;
  assign n162 = n161 ^ n158 ;
  assign n163 = n162 ^ n49 ;
  assign n164 = ~x6 & n163 ;
  assign n167 = n166 ^ n164 ;
  assign n168 = n167 ^ n164 ;
  assign n169 = n164 ^ x6 ;
  assign n170 = n169 ^ n164 ;
  assign n171 = n168 & n170 ;
  assign n172 = n171 ^ n164 ;
  assign n173 = ~x3 & n172 ;
  assign n174 = n173 ^ n164 ;
  assign n175 = ~x7 & n174 ;
  assign n176 = ~x6 & n98 ;
  assign n177 = x8 ^ x3 ;
  assign n178 = n177 ^ x8 ;
  assign n179 = n126 ^ x8 ;
  assign n180 = n178 & n179 ;
  assign n181 = n180 ^ x8 ;
  assign n182 = ~x4 & n181 ;
  assign n183 = ~x10 & ~n182 ;
  assign n184 = n176 & ~n183 ;
  assign n185 = ~n175 & ~n184 ;
  assign n186 = ~x13 & ~n80 ;
  assign n187 = x9 & ~x14 ;
  assign n188 = n18 & n187 ;
  assign n189 = n188 ^ x8 ;
  assign n190 = n189 ^ n188 ;
  assign n191 = n190 ^ x10 ;
  assign n192 = n34 ^ x9 ;
  assign n193 = n34 & ~n192 ;
  assign n194 = n193 ^ n188 ;
  assign n195 = n194 ^ n34 ;
  assign n196 = ~n191 & n195 ;
  assign n197 = n196 ^ n193 ;
  assign n198 = n197 ^ n34 ;
  assign n199 = x10 & n198 ;
  assign n200 = n199 ^ x10 ;
  assign n201 = n186 & ~n200 ;
  assign n202 = ~x2 & n201 ;
  assign n203 = ~n185 & n202 ;
  assign n204 = n24 & n45 ;
  assign n205 = n101 & n204 ;
  assign n206 = ~n33 & n80 ;
  assign n207 = x6 & ~n165 ;
  assign n208 = n206 & ~n207 ;
  assign n209 = n205 & n208 ;
  assign n210 = ~n19 & ~n36 ;
  assign n211 = ~x8 & n24 ;
  assign n212 = ~n210 & n211 ;
  assign n213 = ~n209 & ~n212 ;
  assign n214 = ~n203 & n213 ;
  assign n215 = x5 & ~n214 ;
  assign n216 = x2 & n166 ;
  assign n217 = n54 & n216 ;
  assign n218 = x3 & n217 ;
  assign n219 = ~n215 & ~n218 ;
  assign n220 = ~x0 & ~n219 ;
  assign n221 = ~n152 & ~n220 ;
  assign n222 = ~x3 & x6 ;
  assign n223 = ~x7 & ~x10 ;
  assign n224 = n204 & n223 ;
  assign n225 = n224 ^ n16 ;
  assign n226 = n225 ^ x0 ;
  assign n235 = n226 ^ n225 ;
  assign n227 = x10 & n45 ;
  assign n228 = n79 & n227 ;
  assign n229 = n228 ^ n226 ;
  assign n230 = n229 ^ n225 ;
  assign n231 = n226 ^ n224 ;
  assign n232 = n231 ^ n228 ;
  assign n233 = n232 ^ n230 ;
  assign n234 = n230 & ~n233 ;
  assign n236 = n235 ^ n234 ;
  assign n237 = n236 ^ n230 ;
  assign n238 = n225 ^ n25 ;
  assign n239 = n234 ^ n230 ;
  assign n240 = ~n238 & n239 ;
  assign n241 = n240 ^ n225 ;
  assign n242 = ~n237 & n241 ;
  assign n243 = n242 ^ n225 ;
  assign n244 = n243 ^ n16 ;
  assign n245 = n244 ^ n225 ;
  assign n246 = n222 & n245 ;
  assign n247 = ~x6 & ~x9 ;
  assign n248 = n223 & n247 ;
  assign n249 = n79 & n248 ;
  assign n250 = ~x3 & n249 ;
  assign n251 = n99 & n227 ;
  assign n252 = n33 & n251 ;
  assign n253 = ~n250 & ~n252 ;
  assign n254 = ~n246 & n253 ;
  assign n255 = ~x8 & ~n254 ;
  assign n256 = n16 & n83 ;
  assign n257 = ~x14 & n256 ;
  assign n258 = x7 & ~x13 ;
  assign n259 = n258 ^ n83 ;
  assign n260 = n259 ^ x8 ;
  assign n261 = x9 & n78 ;
  assign n262 = n261 ^ n187 ;
  assign n263 = n83 & ~n262 ;
  assign n264 = n263 ^ n261 ;
  assign n265 = n260 & n264 ;
  assign n266 = n265 ^ n263 ;
  assign n267 = n266 ^ n261 ;
  assign n268 = n267 ^ n83 ;
  assign n269 = x8 & n268 ;
  assign n270 = ~x2 & n269 ;
  assign n271 = ~n257 & ~n270 ;
  assign n272 = n82 & ~n271 ;
  assign n273 = ~x13 & n256 ;
  assign n274 = n20 & n273 ;
  assign n275 = ~n272 & ~n274 ;
  assign n276 = x6 & ~n275 ;
  assign n277 = ~n255 & ~n276 ;
  assign n278 = ~x4 & ~n277 ;
  assign n279 = ~x5 & n278 ;
  assign n280 = x8 & ~x9 ;
  assign n281 = x2 & ~x4 ;
  assign n282 = n280 & n281 ;
  assign n283 = n176 & n282 ;
  assign n284 = x10 ^ x6 ;
  assign n285 = x14 ^ x9 ;
  assign n286 = x10 ^ x9 ;
  assign n287 = n286 ^ x9 ;
  assign n288 = n285 & ~n287 ;
  assign n289 = n288 ^ x9 ;
  assign n290 = ~n284 & ~n289 ;
  assign n291 = n98 & n290 ;
  assign n292 = n291 ^ n109 ;
  assign n293 = x4 & ~x9 ;
  assign n294 = n293 ^ n291 ;
  assign n295 = n294 ^ n293 ;
  assign n296 = n295 ^ n292 ;
  assign n297 = x6 & ~x14 ;
  assign n298 = n223 & n297 ;
  assign n299 = n298 ^ x1 ;
  assign n300 = x1 & n299 ;
  assign n301 = n300 ^ n293 ;
  assign n302 = n301 ^ x1 ;
  assign n303 = ~n296 & ~n302 ;
  assign n304 = n303 ^ n300 ;
  assign n305 = n304 ^ x1 ;
  assign n306 = n292 & n305 ;
  assign n307 = n306 ^ n291 ;
  assign n308 = n307 ^ x8 ;
  assign n309 = n308 ^ n307 ;
  assign n310 = n293 & n298 ;
  assign n311 = ~x1 & n310 ;
  assign n312 = n311 ^ n307 ;
  assign n313 = n309 & n312 ;
  assign n314 = n313 ^ n307 ;
  assign n315 = ~x2 & n314 ;
  assign n316 = ~n283 & ~n315 ;
  assign n317 = ~x13 & ~n316 ;
  assign n318 = ~n65 & n216 ;
  assign n319 = ~n317 & ~n318 ;
  assign n320 = n319 ^ x6 ;
  assign n321 = n320 ^ x0 ;
  assign n348 = n321 ^ n320 ;
  assign n322 = ~x2 & n49 ;
  assign n323 = x9 ^ x8 ;
  assign n324 = n286 & n323 ;
  assign n325 = n322 & n324 ;
  assign n326 = ~x10 & n165 ;
  assign n327 = x0 & ~n326 ;
  assign n328 = x4 & ~n280 ;
  assign n329 = n24 & n328 ;
  assign n330 = n327 & n329 ;
  assign n331 = n47 & n280 ;
  assign n332 = n280 ^ x0 ;
  assign n333 = ~x2 & ~x14 ;
  assign n334 = n333 ^ n331 ;
  assign n335 = ~n332 & n334 ;
  assign n336 = n335 ^ n333 ;
  assign n337 = n331 & n336 ;
  assign n338 = ~x10 & n337 ;
  assign n339 = ~n330 & ~n338 ;
  assign n340 = ~n325 & n339 ;
  assign n341 = n258 & ~n340 ;
  assign n342 = n341 ^ n321 ;
  assign n343 = n342 ^ n320 ;
  assign n344 = n321 ^ n319 ;
  assign n345 = n344 ^ n341 ;
  assign n346 = n345 ^ n343 ;
  assign n347 = n343 & ~n346 ;
  assign n349 = n348 ^ n347 ;
  assign n350 = n349 ^ n343 ;
  assign n351 = n127 & n281 ;
  assign n352 = ~n322 & ~n351 ;
  assign n355 = n352 ^ x10 ;
  assign n356 = n355 ^ n352 ;
  assign n353 = n352 ^ n109 ;
  assign n354 = n353 ^ n352 ;
  assign n357 = n356 ^ n354 ;
  assign n358 = x1 & ~x2 ;
  assign n359 = x8 & ~x13 ;
  assign n360 = ~n358 & n359 ;
  assign n361 = n360 ^ n352 ;
  assign n362 = n361 ^ n352 ;
  assign n363 = n362 ^ n356 ;
  assign n364 = ~n356 & ~n363 ;
  assign n365 = n364 ^ n356 ;
  assign n366 = ~n357 & ~n365 ;
  assign n367 = n366 ^ n364 ;
  assign n368 = n367 ^ n352 ;
  assign n369 = n368 ^ n356 ;
  assign n370 = ~x7 & n369 ;
  assign n371 = n370 ^ n352 ;
  assign n372 = n371 ^ n320 ;
  assign n373 = n347 ^ n343 ;
  assign n374 = ~n372 & n373 ;
  assign n375 = n374 ^ n320 ;
  assign n376 = ~n350 & ~n375 ;
  assign n377 = n376 ^ n320 ;
  assign n378 = n377 ^ x6 ;
  assign n379 = n378 ^ n320 ;
  assign n380 = n133 & n379 ;
  assign n381 = ~n279 & ~n380 ;
  assign n382 = n221 & n381 ;
  assign n383 = ~x12 & ~n382 ;
  assign n384 = ~n77 & ~n383 ;
  assign n385 = ~x11 & ~n384 ;
  assign y0 = n385 ;
endmodule
