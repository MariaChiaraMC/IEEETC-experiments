module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 ;
  assign n10 = x7 & x8 ;
  assign n11 = x3 & x4 ;
  assign n12 = x5 & n11 ;
  assign n13 = n10 & n12 ;
  assign n14 = x2 & x5 ;
  assign n15 = n14 ^ x7 ;
  assign n16 = x4 & x8 ;
  assign n17 = n16 ^ x3 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = n16 ^ x4 ;
  assign n20 = n18 & ~n19 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = n21 ^ n14 ;
  assign n23 = ~n15 & n22 ;
  assign n24 = n23 ^ n20 ;
  assign n25 = n24 ^ n16 ;
  assign n26 = n25 ^ x7 ;
  assign n27 = n14 & ~n26 ;
  assign n28 = n27 ^ n14 ;
  assign n29 = ~n13 & ~n28 ;
  assign n30 = ~x2 & ~x5 ;
  assign n31 = ~x4 & ~x8 ;
  assign n32 = x3 & ~n31 ;
  assign n33 = n30 & ~n32 ;
  assign n37 = ~x3 & x5 ;
  assign n34 = ~x2 & ~x3 ;
  assign n35 = ~n30 & ~n34 ;
  assign n36 = n35 ^ x7 ;
  assign n38 = n37 ^ n36 ;
  assign n41 = n38 ^ n16 ;
  assign n42 = n41 ^ n38 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n39 ^ x7 ;
  assign n43 = n42 ^ n40 ;
  assign n44 = n40 ^ x7 ;
  assign n45 = n43 & n44 ;
  assign n46 = n45 ^ n36 ;
  assign n47 = n46 ^ n40 ;
  assign n48 = n47 ^ x7 ;
  assign n49 = ~x2 & x5 ;
  assign n50 = x4 & n49 ;
  assign n51 = x3 & x8 ;
  assign n52 = ~n50 & ~n51 ;
  assign n53 = n52 ^ n36 ;
  assign n54 = n53 ^ x7 ;
  assign n55 = n40 ^ n36 ;
  assign n56 = n55 ^ n42 ;
  assign n57 = n56 ^ x7 ;
  assign n58 = n56 & ~n57 ;
  assign n59 = n58 ^ n36 ;
  assign n60 = n59 ^ n40 ;
  assign n61 = n60 ^ n42 ;
  assign n62 = ~n54 & n61 ;
  assign n63 = n62 ^ x7 ;
  assign n64 = n48 & ~n63 ;
  assign n65 = n64 ^ n45 ;
  assign n66 = n65 ^ n40 ;
  assign n67 = n66 ^ x7 ;
  assign n68 = n67 ^ n35 ;
  assign n69 = n68 ^ n36 ;
  assign n70 = ~n33 & n69 ;
  assign n71 = n70 ^ x6 ;
  assign n72 = n71 ^ n70 ;
  assign n73 = ~x7 & ~n16 ;
  assign n74 = x7 & n16 ;
  assign n75 = ~x3 & ~n74 ;
  assign n76 = ~n73 & ~n75 ;
  assign n77 = n49 & n76 ;
  assign n78 = x2 & ~x5 ;
  assign n79 = ~n11 & ~n78 ;
  assign n80 = n10 & ~n79 ;
  assign n81 = ~n77 & ~n80 ;
  assign n82 = n81 ^ n70 ;
  assign n83 = ~n72 & n82 ;
  assign n84 = n83 ^ n70 ;
  assign n85 = n29 & n84 ;
  assign n86 = x1 & ~n85 ;
  assign n87 = ~x1 & n76 ;
  assign n88 = x3 & n10 ;
  assign n89 = ~n87 & ~n88 ;
  assign n90 = x6 & n78 ;
  assign n91 = ~n89 & n90 ;
  assign n92 = x7 ^ x6 ;
  assign n93 = n92 ^ x4 ;
  assign n94 = n93 ^ x7 ;
  assign n95 = n94 ^ n92 ;
  assign n102 = n92 ^ x8 ;
  assign n103 = n102 ^ x7 ;
  assign n104 = n103 ^ x7 ;
  assign n105 = n104 ^ n92 ;
  assign n97 = x6 ^ x1 ;
  assign n96 = n92 ^ x7 ;
  assign n98 = n97 ^ n96 ;
  assign n106 = n105 ^ n98 ;
  assign n100 = x6 ^ x3 ;
  assign n99 = n98 ^ n97 ;
  assign n101 = n100 ^ n99 ;
  assign n107 = n106 ^ n101 ;
  assign n108 = n107 ^ n95 ;
  assign n109 = ~n95 & n108 ;
  assign n110 = n109 ^ n106 ;
  assign n111 = n100 ^ n98 ;
  assign n112 = n111 ^ n101 ;
  assign n113 = n104 ^ n98 ;
  assign n119 = n113 ^ n101 ;
  assign n120 = n119 ^ n106 ;
  assign n121 = n100 & n120 ;
  assign n114 = n113 ^ n106 ;
  assign n115 = n104 ^ n101 ;
  assign n116 = n115 ^ n106 ;
  assign n117 = n116 ^ n95 ;
  assign n118 = n114 & n117 ;
  assign n122 = n121 ^ n118 ;
  assign n123 = n122 ^ n104 ;
  assign n124 = n123 ^ n100 ;
  assign n125 = n124 ^ n106 ;
  assign n126 = n125 ^ n95 ;
  assign n127 = ~n112 & n126 ;
  assign n128 = n127 ^ n118 ;
  assign n129 = n128 ^ n104 ;
  assign n130 = n129 ^ n100 ;
  assign n131 = n130 ^ n98 ;
  assign n132 = n131 ^ n101 ;
  assign n133 = n132 ^ n106 ;
  assign n134 = n133 ^ n95 ;
  assign n135 = ~n110 & ~n134 ;
  assign n136 = n135 ^ n121 ;
  assign n137 = n136 ^ n109 ;
  assign n138 = n137 ^ n106 ;
  assign n139 = n138 ^ x6 ;
  assign n140 = n139 ^ n100 ;
  assign n141 = n14 & n140 ;
  assign n142 = ~x1 & x6 ;
  assign n143 = n142 ^ x2 ;
  assign n144 = n143 ^ n12 ;
  assign n145 = n10 ^ x7 ;
  assign n146 = ~x2 & ~n145 ;
  assign n147 = n146 ^ x7 ;
  assign n148 = ~n144 & n147 ;
  assign n149 = n148 ^ n146 ;
  assign n150 = n149 ^ x7 ;
  assign n151 = n150 ^ x2 ;
  assign n152 = n12 & ~n151 ;
  assign n153 = ~n141 & ~n152 ;
  assign n154 = ~n91 & n153 ;
  assign n155 = ~n86 & n154 ;
  assign y0 = ~n155 ;
endmodule
