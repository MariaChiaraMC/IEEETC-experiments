module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n12 = ~x0 & ~x1 ;
  assign n13 = ~x2 & x6 ;
  assign n14 = n12 & n13 ;
  assign n15 = ~x3 & ~x10 ;
  assign n16 = ~x9 & n15 ;
  assign n17 = n14 & n16 ;
  assign n18 = x5 ^ x4 ;
  assign n19 = x8 ^ x4 ;
  assign n20 = x8 ^ x7 ;
  assign n21 = ~x8 & ~n20 ;
  assign n22 = n21 ^ x8 ;
  assign n23 = ~n19 & ~n22 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n24 ^ x8 ;
  assign n26 = n25 ^ x7 ;
  assign n27 = n18 & ~n26 ;
  assign n28 = n17 & n27 ;
  assign y0 = n28 ;
endmodule
