module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 ;
  assign n16 = ~x4 & ~x5 ;
  assign n17 = ~x6 & ~x8 ;
  assign n18 = ~x7 & x10 ;
  assign n19 = ~n17 & n18 ;
  assign n20 = n16 & n19 ;
  assign n24 = ~x6 & x14 ;
  assign n21 = ~x0 & ~x12 ;
  assign n22 = x9 & ~x13 ;
  assign n23 = n21 & n22 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = x12 & x13 ;
  assign n28 = n27 ^ n23 ;
  assign n29 = n28 ^ n23 ;
  assign n30 = n26 & n29 ;
  assign n31 = n30 ^ n23 ;
  assign n32 = ~x11 & n31 ;
  assign n33 = n32 ^ n23 ;
  assign n34 = n20 & n33 ;
  assign n35 = ~x10 & ~x11 ;
  assign n36 = ~x13 & n35 ;
  assign n37 = ~x7 & ~x8 ;
  assign n38 = x6 & n16 ;
  assign n39 = ~n37 & n38 ;
  assign n40 = n39 ^ x3 ;
  assign n41 = n40 ^ x12 ;
  assign n48 = n41 ^ n40 ;
  assign n42 = n41 ^ x14 ;
  assign n43 = n42 ^ n40 ;
  assign n44 = n39 ^ x14 ;
  assign n45 = n44 ^ x14 ;
  assign n46 = n45 ^ n43 ;
  assign n47 = n43 & n46 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = n49 ^ n43 ;
  assign n51 = n40 ^ x0 ;
  assign n52 = n47 ^ n43 ;
  assign n53 = n51 & n52 ;
  assign n54 = n53 ^ n40 ;
  assign n55 = n50 & n54 ;
  assign n56 = n55 ^ n40 ;
  assign n57 = n56 ^ n39 ;
  assign n58 = n57 ^ n40 ;
  assign n59 = n36 & n58 ;
  assign n60 = ~n34 & ~n59 ;
  assign n61 = ~x3 & x11 ;
  assign n62 = x5 & ~x13 ;
  assign n63 = x14 & n62 ;
  assign n64 = ~n61 & ~n63 ;
  assign n65 = ~x10 & ~n64 ;
  assign n66 = ~x0 & n63 ;
  assign n67 = x4 & n66 ;
  assign n68 = n67 ^ x11 ;
  assign n69 = n68 ^ n67 ;
  assign n70 = x13 & ~x14 ;
  assign n71 = x4 & x7 ;
  assign n72 = ~x5 & n71 ;
  assign n73 = x1 & x3 ;
  assign n74 = n72 & n73 ;
  assign n75 = n70 & ~n74 ;
  assign n76 = ~x3 & x13 ;
  assign n77 = x1 & n76 ;
  assign n78 = ~x10 & ~n77 ;
  assign n79 = x5 & x6 ;
  assign n80 = x0 & ~n79 ;
  assign n81 = x5 & ~x7 ;
  assign n82 = x10 & x13 ;
  assign n83 = x14 & ~n82 ;
  assign n84 = ~n81 & ~n83 ;
  assign n85 = x4 & n84 ;
  assign n86 = ~n80 & n85 ;
  assign n87 = ~n78 & ~n86 ;
  assign n88 = ~n75 & n87 ;
  assign n89 = n88 ^ n67 ;
  assign n90 = ~n69 & ~n89 ;
  assign n91 = n90 ^ n67 ;
  assign n92 = ~x1 & ~x6 ;
  assign n93 = n67 & ~n92 ;
  assign n94 = n93 ^ n65 ;
  assign n95 = n91 & ~n94 ;
  assign n96 = n95 ^ n93 ;
  assign n97 = ~n65 & n96 ;
  assign n98 = n97 ^ n65 ;
  assign n99 = ~x12 & n98 ;
  assign n100 = x12 & ~x13 ;
  assign n101 = ~x4 & n100 ;
  assign n102 = ~x13 & n16 ;
  assign n103 = x7 & x8 ;
  assign n104 = ~x6 & ~x14 ;
  assign n105 = n103 & n104 ;
  assign n106 = n102 & n105 ;
  assign n107 = ~x2 & n62 ;
  assign n108 = n107 ^ x1 ;
  assign n109 = n107 ^ n72 ;
  assign n110 = n70 & n109 ;
  assign n111 = n110 ^ x6 ;
  assign n112 = ~x1 & ~n111 ;
  assign n113 = n112 ^ n110 ;
  assign n114 = ~n108 & n113 ;
  assign n115 = n114 ^ n107 ;
  assign n116 = n115 ^ n110 ;
  assign n117 = n116 ^ n112 ;
  assign n118 = ~x0 & n117 ;
  assign n119 = x12 & n118 ;
  assign n120 = ~n106 & ~n119 ;
  assign n121 = ~n101 & n120 ;
  assign n122 = x11 & ~n121 ;
  assign n123 = x7 & n16 ;
  assign n124 = ~x8 & n24 ;
  assign n125 = n100 & n124 ;
  assign n126 = n123 & n125 ;
  assign n127 = ~n122 & ~n126 ;
  assign n128 = n127 ^ x10 ;
  assign n129 = n128 ^ n127 ;
  assign n130 = n129 ^ n99 ;
  assign n131 = x4 & x12 ;
  assign n132 = x14 & ~n131 ;
  assign n133 = n132 ^ x11 ;
  assign n134 = ~x11 & n133 ;
  assign n135 = n134 ^ n127 ;
  assign n136 = n135 ^ x11 ;
  assign n137 = n130 & n136 ;
  assign n138 = n137 ^ n134 ;
  assign n139 = n138 ^ x11 ;
  assign n140 = ~n99 & ~n139 ;
  assign n141 = n140 ^ n99 ;
  assign n142 = n141 ^ x9 ;
  assign n143 = n142 ^ n141 ;
  assign n144 = n143 ^ n60 ;
  assign n145 = n24 & n61 ;
  assign n146 = x8 ^ x7 ;
  assign n147 = ~n81 & n146 ;
  assign n148 = n145 & ~n147 ;
  assign n149 = n100 & ~n148 ;
  assign n150 = x13 ^ x11 ;
  assign n151 = n21 ^ x13 ;
  assign n152 = n151 ^ n21 ;
  assign n153 = ~x1 & ~x12 ;
  assign n154 = x14 & n153 ;
  assign n155 = x0 & n154 ;
  assign n156 = n155 ^ n21 ;
  assign n157 = ~n152 & ~n156 ;
  assign n158 = n157 ^ n21 ;
  assign n159 = n150 & n158 ;
  assign n160 = n159 ^ x11 ;
  assign n161 = ~n149 & ~n160 ;
  assign n162 = n161 ^ x10 ;
  assign n163 = ~x10 & n162 ;
  assign n164 = n163 ^ n141 ;
  assign n165 = n164 ^ x10 ;
  assign n166 = n144 & ~n165 ;
  assign n167 = n166 ^ n163 ;
  assign n168 = n167 ^ x10 ;
  assign n169 = n60 & ~n168 ;
  assign n170 = n169 ^ n60 ;
  assign y0 = ~n170 ;
endmodule
