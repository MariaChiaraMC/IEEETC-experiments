// Benchmark "./pla/risc.pla_res_27NonExact" written by ABC on Fri Nov 20 10:29:13 2020

module \./pla/risc.pla_res_27NonExact  ( 
    x0, x1,
    z0  );
  input  x0, x1;
  output z0;
  assign z0 = ~x0 & x1;
endmodule


