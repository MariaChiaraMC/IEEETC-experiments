module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 ;
  assign n20 = x5 ^ x3 ;
  assign n21 = n20 ^ x5 ;
  assign n16 = x5 & ~x8 ;
  assign n22 = n16 ^ x5 ;
  assign n23 = n21 & ~n22 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = x2 & n24 ;
  assign n13 = x2 & x3 ;
  assign n14 = ~x4 & ~x10 ;
  assign n15 = n13 & ~n14 ;
  assign n17 = ~n15 & n16 ;
  assign n26 = n25 ^ n17 ;
  assign n27 = n26 ^ n17 ;
  assign n18 = n17 ^ x4 ;
  assign n19 = n18 ^ n17 ;
  assign n28 = n27 ^ n19 ;
  assign n29 = x8 & ~x10 ;
  assign n30 = n29 ^ x2 ;
  assign n31 = n29 ^ x3 ;
  assign n32 = n31 ^ x3 ;
  assign n33 = ~n20 & n32 ;
  assign n34 = n33 ^ x3 ;
  assign n35 = n30 & ~n34 ;
  assign n36 = n35 ^ x2 ;
  assign n37 = n36 ^ n17 ;
  assign n38 = n37 ^ n17 ;
  assign n39 = n38 ^ n27 ;
  assign n40 = ~n27 & ~n39 ;
  assign n41 = n40 ^ n27 ;
  assign n42 = ~n28 & ~n41 ;
  assign n43 = n42 ^ n40 ;
  assign n44 = n43 ^ n17 ;
  assign n45 = n44 ^ n27 ;
  assign n46 = x7 & ~n45 ;
  assign n47 = n46 ^ n17 ;
  assign y0 = n47 ;
endmodule
