module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 ;
  assign n17 = x4 & ~x5 ;
  assign n18 = ~x3 & ~n17 ;
  assign n36 = x7 & ~n18 ;
  assign n37 = n36 ^ x3 ;
  assign n16 = ~x4 & ~x9 ;
  assign n38 = n36 ^ n16 ;
  assign n39 = n38 ^ n16 ;
  assign n20 = x9 ^ x5 ;
  assign n21 = x4 & ~n20 ;
  assign n22 = n21 ^ x5 ;
  assign n40 = n22 ^ n16 ;
  assign n41 = n39 & n40 ;
  assign n42 = n41 ^ n16 ;
  assign n43 = ~n37 & ~n42 ;
  assign n44 = n43 ^ x3 ;
  assign n45 = n44 ^ x9 ;
  assign n46 = n45 ^ x1 ;
  assign n53 = n46 ^ n45 ;
  assign n47 = n46 ^ x7 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = n46 ^ n44 ;
  assign n50 = n49 ^ x7 ;
  assign n51 = n50 ^ n48 ;
  assign n52 = n48 & n51 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = n54 ^ n48 ;
  assign n56 = n45 ^ x5 ;
  assign n57 = n52 ^ n48 ;
  assign n58 = n56 & n57 ;
  assign n59 = n58 ^ n45 ;
  assign n60 = n55 & n59 ;
  assign n61 = n60 ^ n45 ;
  assign n62 = n61 ^ x9 ;
  assign n63 = n62 ^ n45 ;
  assign n12 = x2 & x8 ;
  assign n13 = n12 ^ x7 ;
  assign n14 = n12 ^ x9 ;
  assign n15 = n14 ^ x9 ;
  assign n19 = ~n16 & n18 ;
  assign n23 = x3 & n22 ;
  assign n24 = n23 ^ x1 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = ~x5 & ~x9 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = ~n25 & ~n27 ;
  assign n29 = n28 ^ n23 ;
  assign n30 = ~n19 & ~n29 ;
  assign n31 = n30 ^ x9 ;
  assign n32 = ~n15 & ~n31 ;
  assign n33 = n32 ^ x9 ;
  assign n34 = n13 & ~n33 ;
  assign n35 = n34 ^ x7 ;
  assign n64 = n63 ^ n35 ;
  assign n65 = n64 ^ n35 ;
  assign n66 = n35 ^ n12 ;
  assign n67 = n66 ^ n35 ;
  assign n68 = ~n65 & ~n67 ;
  assign n69 = n68 ^ n35 ;
  assign n70 = x6 & n69 ;
  assign n71 = n70 ^ n35 ;
  assign n72 = ~x10 & n71 ;
  assign n73 = x7 & x10 ;
  assign n74 = ~x9 & n73 ;
  assign n75 = ~x4 & x5 ;
  assign n76 = x1 & ~x2 ;
  assign n77 = ~n18 & n76 ;
  assign n78 = ~n75 & n77 ;
  assign n79 = ~x0 & ~n78 ;
  assign n80 = n79 ^ x6 ;
  assign n81 = n74 & n80 ;
  assign n82 = ~x8 & n81 ;
  assign n83 = ~n72 & ~n82 ;
  assign y0 = ~n83 ;
endmodule
