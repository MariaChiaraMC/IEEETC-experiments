module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 ;
  assign n11 = ~x2 & x8 ;
  assign n12 = x7 & x9 ;
  assign n13 = n11 & n12 ;
  assign n14 = n13 ^ x6 ;
  assign n15 = x1 & ~x3 ;
  assign n16 = ~x4 & ~x5 ;
  assign n17 = ~n15 & n16 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = n17 ^ x0 ;
  assign n20 = ~n17 & n19 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = ~n18 & ~n21 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n23 ^ n17 ;
  assign n25 = n24 ^ x0 ;
  assign n26 = n14 & n25 ;
  assign y0 = n26 ;
endmodule
