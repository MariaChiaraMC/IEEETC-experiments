module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n13 = x8 & ~x11 ;
  assign n14 = n13 ^ x9 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = n15 ^ x10 ;
  assign n17 = ~x2 & ~x8 ;
  assign n18 = ~x1 & x6 ;
  assign n19 = n17 & n18 ;
  assign n20 = x4 & x7 ;
  assign n21 = ~x3 & n20 ;
  assign n22 = n19 & ~n21 ;
  assign n23 = ~x0 & n22 ;
  assign n24 = n23 ^ x10 ;
  assign n25 = x5 & n24 ;
  assign n26 = n25 ^ n13 ;
  assign n27 = n16 & ~n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = x10 & n28 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n31 ^ x9 ;
  assign y0 = n32 ;
endmodule
