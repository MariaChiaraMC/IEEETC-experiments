module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 ;
  assign n22 = x16 ^ x15 ;
  assign n23 = x18 & x19 ;
  assign n24 = ~x4 & x20 ;
  assign n25 = n23 & n24 ;
  assign n26 = n25 ^ x15 ;
  assign n27 = n26 ^ x15 ;
  assign n28 = n27 ^ n22 ;
  assign n29 = ~n22 & ~n28 ;
  assign n30 = n29 ^ x15 ;
  assign n31 = n30 ^ n22 ;
  assign n32 = x6 & ~x17 ;
  assign n33 = n32 ^ x15 ;
  assign n34 = n33 ^ x0 ;
  assign n35 = n32 & n34 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ x15 ;
  assign n38 = n32 ^ x3 ;
  assign n39 = ~n33 & n38 ;
  assign n40 = n39 ^ x3 ;
  assign n41 = n40 ^ x0 ;
  assign n42 = ~n37 & ~n41 ;
  assign n43 = n42 ^ x0 ;
  assign n44 = n31 & ~n43 ;
  assign n45 = n44 ^ n42 ;
  assign n46 = n45 ^ x0 ;
  assign y0 = ~n46 ;
endmodule
