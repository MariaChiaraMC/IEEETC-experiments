module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 ;
  assign n15 = ~x4 & ~x5 ;
  assign n16 = x1 & x2 ;
  assign n17 = ~x3 & n16 ;
  assign n18 = ~n15 & n17 ;
  assign n19 = ~x1 & ~x10 ;
  assign n20 = x5 ^ x4 ;
  assign n21 = x5 ^ x2 ;
  assign n22 = x5 ^ x3 ;
  assign n23 = ~x5 & ~n22 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = ~n21 & ~n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n26 ^ x5 ;
  assign n28 = n27 ^ x3 ;
  assign n29 = ~n20 & ~n28 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = n19 & ~n30 ;
  assign n32 = ~x7 & x8 ;
  assign n33 = ~x9 & n32 ;
  assign n34 = x11 & x13 ;
  assign n35 = ~x6 & ~n34 ;
  assign n36 = n33 & n35 ;
  assign n37 = ~x11 & ~x13 ;
  assign n38 = n37 ^ x12 ;
  assign n39 = n36 & ~n38 ;
  assign n40 = n31 & n39 ;
  assign n41 = ~n18 & ~n40 ;
  assign n42 = n41 ^ x1 ;
  assign n43 = n42 ^ n41 ;
  assign n44 = n41 ^ x5 ;
  assign n45 = n44 ^ n41 ;
  assign n46 = ~n43 & ~n45 ;
  assign n47 = n46 ^ n41 ;
  assign n48 = x0 & ~n47 ;
  assign n49 = n48 ^ n41 ;
  assign y0 = ~n49 ;
endmodule
