module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 ;
  assign n11 = x6 & x7 ;
  assign n12 = x5 & x9 ;
  assign n13 = ~x2 & x3 ;
  assign n14 = x0 & n13 ;
  assign n15 = n12 & n14 ;
  assign n16 = ~x4 & n15 ;
  assign n17 = n16 ^ x8 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = n18 ^ n11 ;
  assign n20 = x0 & ~x5 ;
  assign n21 = x2 & ~x3 ;
  assign n22 = n21 ^ n13 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = n21 ^ x9 ;
  assign n25 = n21 ^ x4 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = ~n24 & n26 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = n28 ^ n24 ;
  assign n30 = n23 & ~n29 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = n20 & ~n32 ;
  assign n34 = ~x2 & x4 ;
  assign n35 = ~x0 & x3 ;
  assign n36 = x5 & ~x9 ;
  assign n37 = n35 & n36 ;
  assign n38 = n34 & n37 ;
  assign n39 = n38 ^ n33 ;
  assign n40 = ~n33 & n39 ;
  assign n41 = n40 ^ n16 ;
  assign n42 = n41 ^ n33 ;
  assign n43 = n19 & n42 ;
  assign n44 = n43 ^ n40 ;
  assign n45 = n44 ^ n33 ;
  assign n46 = n11 & ~n45 ;
  assign n47 = n46 ^ n11 ;
  assign n48 = ~x4 & ~x9 ;
  assign n49 = ~x3 & ~x5 ;
  assign n50 = x8 & n49 ;
  assign n51 = n48 & n50 ;
  assign n52 = x7 ^ x0 ;
  assign n53 = x2 & n52 ;
  assign n54 = n51 & n53 ;
  assign n61 = ~x7 & ~x8 ;
  assign n55 = x8 & x9 ;
  assign n101 = ~x8 & ~x9 ;
  assign n102 = ~n55 & ~n101 ;
  assign n103 = x3 & x5 ;
  assign n104 = ~n102 & n103 ;
  assign n105 = ~n61 & n104 ;
  assign n106 = n105 ^ x2 ;
  assign n107 = n106 ^ n105 ;
  assign n108 = n105 ^ n49 ;
  assign n109 = n108 ^ n106 ;
  assign n116 = n109 ^ n106 ;
  assign n117 = n116 ^ n105 ;
  assign n110 = x7 & ~x9 ;
  assign n111 = n110 ^ n109 ;
  assign n112 = n111 ^ x8 ;
  assign n113 = n112 ^ n111 ;
  assign n114 = n113 ^ n105 ;
  assign n115 = n114 ^ n107 ;
  assign n118 = n117 ^ n115 ;
  assign n119 = ~n107 & n118 ;
  assign n120 = n119 ^ n113 ;
  assign n121 = n120 ^ n117 ;
  assign n127 = n111 ^ n109 ;
  assign n122 = ~x7 & x9 ;
  assign n123 = n122 ^ n111 ;
  assign n124 = n117 ^ n113 ;
  assign n125 = ~n123 & ~n124 ;
  assign n126 = n125 ^ n119 ;
  assign n128 = n127 ^ n126 ;
  assign n129 = n128 ^ n123 ;
  assign n130 = n129 ^ n113 ;
  assign n131 = n117 & n130 ;
  assign n132 = n131 ^ n107 ;
  assign n133 = ~n121 & ~n132 ;
  assign n134 = n133 ^ n107 ;
  assign n135 = n134 ^ x2 ;
  assign n136 = n135 ^ n107 ;
  assign n137 = x0 & ~n136 ;
  assign n56 = x2 & x3 ;
  assign n57 = n20 & n56 ;
  assign n58 = n55 & n57 ;
  assign n59 = x7 & n58 ;
  assign n60 = x7 & x8 ;
  assign n62 = ~n60 & ~n61 ;
  assign n63 = ~x2 & ~x9 ;
  assign n64 = x3 & ~x7 ;
  assign n65 = ~x0 & ~x5 ;
  assign n66 = ~n64 & n65 ;
  assign n67 = n63 & n66 ;
  assign n68 = ~n62 & n67 ;
  assign n69 = x8 ^ x0 ;
  assign n70 = n21 ^ x8 ;
  assign n71 = n70 ^ n21 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = ~x2 & ~x7 ;
  assign n74 = x2 & x7 ;
  assign n75 = ~n73 & ~n74 ;
  assign n76 = n75 ^ x3 ;
  assign n77 = ~n75 & ~n76 ;
  assign n78 = n77 ^ n21 ;
  assign n79 = n78 ^ n75 ;
  assign n80 = n72 & ~n79 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n81 ^ n75 ;
  assign n83 = ~n69 & ~n82 ;
  assign n84 = n36 & n83 ;
  assign n85 = ~n68 & ~n84 ;
  assign n86 = ~n59 & n85 ;
  assign n87 = ~x7 & x8 ;
  assign n88 = x0 & x5 ;
  assign n89 = n56 & n88 ;
  assign n90 = ~x0 & ~x3 ;
  assign n91 = ~x2 & ~x5 ;
  assign n92 = x9 & n91 ;
  assign n93 = ~n90 & n92 ;
  assign n94 = ~n89 & ~n93 ;
  assign n95 = n87 & ~n94 ;
  assign n96 = x2 & n35 ;
  assign n97 = n12 & n61 ;
  assign n98 = n96 & n97 ;
  assign n99 = ~n95 & ~n98 ;
  assign n100 = n86 & n99 ;
  assign n138 = n137 ^ n100 ;
  assign n139 = n138 ^ n100 ;
  assign n140 = ~x2 & ~x3 ;
  assign n141 = n60 & n140 ;
  assign n142 = n12 & n141 ;
  assign n143 = x9 & n87 ;
  assign n144 = n96 & n143 ;
  assign n145 = ~n142 & ~n144 ;
  assign n146 = n145 ^ n100 ;
  assign n147 = n146 ^ n100 ;
  assign n148 = ~n139 & n147 ;
  assign n149 = n148 ^ n100 ;
  assign n150 = ~x4 & n149 ;
  assign n151 = n150 ^ n100 ;
  assign n152 = ~x6 & ~n151 ;
  assign n153 = x2 & ~x7 ;
  assign n154 = n101 & n153 ;
  assign n155 = x7 & x9 ;
  assign n156 = ~x0 & x2 ;
  assign n157 = ~n155 & n156 ;
  assign n158 = ~n102 & n157 ;
  assign n159 = ~n154 & ~n158 ;
  assign n160 = x5 & ~n159 ;
  assign n161 = x7 ^ x2 ;
  assign n162 = n161 ^ x2 ;
  assign n163 = n91 ^ x2 ;
  assign n164 = n162 & n163 ;
  assign n165 = n164 ^ x2 ;
  assign n166 = n101 & n165 ;
  assign n167 = ~x0 & n166 ;
  assign n168 = ~n160 & ~n167 ;
  assign n169 = ~x4 & ~n168 ;
  assign n170 = n169 ^ x3 ;
  assign n171 = n170 ^ n169 ;
  assign n172 = n171 ^ x6 ;
  assign n173 = n12 & n34 ;
  assign n174 = n48 & n156 ;
  assign n175 = ~x5 & n174 ;
  assign n176 = ~n173 & ~n175 ;
  assign n177 = n87 & ~n176 ;
  assign n178 = ~x4 & ~x5 ;
  assign n179 = x2 & x9 ;
  assign n180 = n178 & n179 ;
  assign n181 = ~n62 & n180 ;
  assign n182 = x0 & n181 ;
  assign n183 = ~n177 & ~n182 ;
  assign n185 = x7 ^ x4 ;
  assign n184 = x8 ^ x4 ;
  assign n186 = n185 ^ n184 ;
  assign n191 = n186 ^ x2 ;
  assign n192 = n191 ^ n186 ;
  assign n187 = n186 ^ x9 ;
  assign n188 = n187 ^ n185 ;
  assign n189 = n188 ^ x4 ;
  assign n190 = n189 ^ n186 ;
  assign n193 = n192 ^ n190 ;
  assign n196 = n189 ^ x4 ;
  assign n194 = n185 ^ x4 ;
  assign n195 = n194 ^ n190 ;
  assign n197 = n196 ^ n195 ;
  assign n198 = ~n193 & n197 ;
  assign n199 = n198 ^ n189 ;
  assign n200 = n199 ^ n194 ;
  assign n201 = n200 ^ n196 ;
  assign n202 = n195 ^ n192 ;
  assign n203 = ~n199 & ~n202 ;
  assign n204 = n203 ^ n189 ;
  assign n205 = n204 ^ n190 ;
  assign n206 = n205 ^ n192 ;
  assign n207 = n201 & n206 ;
  assign n208 = n88 & n207 ;
  assign n209 = n208 ^ n183 ;
  assign n210 = n183 & ~n209 ;
  assign n211 = n210 ^ n169 ;
  assign n212 = n211 ^ n183 ;
  assign n213 = n172 & ~n212 ;
  assign n214 = n213 ^ n210 ;
  assign n215 = n214 ^ n183 ;
  assign n216 = x6 & n215 ;
  assign n217 = n216 ^ x6 ;
  assign n218 = ~n152 & ~n217 ;
  assign n219 = ~n54 & n218 ;
  assign n220 = n219 ^ x1 ;
  assign n221 = n220 ^ n219 ;
  assign n222 = ~x6 & ~x7 ;
  assign n223 = n35 & n173 ;
  assign n224 = n222 & n223 ;
  assign n225 = ~x2 & n90 ;
  assign n226 = n36 & n225 ;
  assign n227 = n222 & n226 ;
  assign n260 = n14 & n122 ;
  assign n261 = x5 & n260 ;
  assign n262 = n35 & n92 ;
  assign n263 = x7 & n90 ;
  assign n264 = n12 & n263 ;
  assign n265 = x9 ^ x7 ;
  assign n266 = n265 ^ x9 ;
  assign n267 = ~x3 & ~x9 ;
  assign n268 = n267 ^ x9 ;
  assign n269 = n266 & n268 ;
  assign n270 = n269 ^ x9 ;
  assign n271 = n88 & n270 ;
  assign n272 = ~n264 & ~n271 ;
  assign n273 = n272 ^ n12 ;
  assign n274 = n273 ^ n272 ;
  assign n275 = n263 ^ n64 ;
  assign n276 = n263 ^ x5 ;
  assign n277 = n276 ^ n275 ;
  assign n278 = x9 ^ x0 ;
  assign n279 = x5 & n278 ;
  assign n280 = n279 ^ x9 ;
  assign n281 = n277 & n280 ;
  assign n282 = n281 ^ n279 ;
  assign n283 = n282 ^ x9 ;
  assign n284 = n283 ^ x5 ;
  assign n285 = n275 & n284 ;
  assign n286 = n285 ^ n64 ;
  assign n287 = n286 ^ n272 ;
  assign n288 = n287 ^ n272 ;
  assign n289 = ~n274 & n288 ;
  assign n290 = n289 ^ n272 ;
  assign n291 = x2 & ~n290 ;
  assign n292 = n291 ^ n272 ;
  assign n293 = ~n262 & n292 ;
  assign n294 = n293 ^ x6 ;
  assign n295 = n294 ^ n293 ;
  assign n296 = ~n63 & ~n153 ;
  assign n235 = ~x7 & ~x9 ;
  assign n297 = n49 & ~n235 ;
  assign n298 = ~x0 & n297 ;
  assign n299 = ~n296 & n298 ;
  assign n300 = ~n14 & ~n88 ;
  assign n301 = x3 ^ x2 ;
  assign n302 = x5 & n301 ;
  assign n303 = n155 & ~n302 ;
  assign n304 = ~n300 & n303 ;
  assign n305 = ~n299 & ~n304 ;
  assign n306 = n305 ^ n293 ;
  assign n307 = n295 & n306 ;
  assign n308 = n307 ^ n293 ;
  assign n309 = ~n261 & n308 ;
  assign n228 = x6 & n56 ;
  assign n229 = ~n225 & ~n228 ;
  assign n230 = n36 & ~n229 ;
  assign n231 = ~x7 & n230 ;
  assign n232 = n35 & n91 ;
  assign n233 = n222 & n232 ;
  assign n234 = ~n231 & ~n233 ;
  assign n236 = ~x5 & n140 ;
  assign n237 = x6 & n103 ;
  assign n238 = ~n236 & ~n237 ;
  assign n239 = n235 & ~n238 ;
  assign n240 = n239 ^ x0 ;
  assign n241 = n240 ^ n239 ;
  assign n242 = n241 ^ n234 ;
  assign n243 = n155 & n228 ;
  assign n244 = x3 & ~n11 ;
  assign n245 = x6 ^ x3 ;
  assign n246 = x9 & ~n245 ;
  assign n247 = n246 ^ x3 ;
  assign n248 = ~n244 & n247 ;
  assign n249 = ~x2 & n248 ;
  assign n250 = ~n243 & ~n249 ;
  assign n251 = n250 ^ x5 ;
  assign n252 = ~n250 & n251 ;
  assign n253 = n252 ^ n239 ;
  assign n254 = n253 ^ n250 ;
  assign n255 = ~n242 & ~n254 ;
  assign n256 = n255 ^ n252 ;
  assign n257 = n256 ^ n250 ;
  assign n258 = n234 & ~n257 ;
  assign n259 = n258 ^ n234 ;
  assign n310 = n309 ^ n259 ;
  assign n311 = ~x4 & n310 ;
  assign n312 = n311 ^ n309 ;
  assign n313 = ~n227 & n312 ;
  assign n314 = n313 ^ x8 ;
  assign n315 = n314 ^ n313 ;
  assign n316 = n13 & n222 ;
  assign n317 = n122 ^ x6 ;
  assign n318 = n317 ^ n122 ;
  assign n319 = n122 ^ n110 ;
  assign n320 = n318 & n319 ;
  assign n321 = n320 ^ n122 ;
  assign n322 = n21 & n321 ;
  assign n323 = ~n316 & ~n322 ;
  assign n324 = n20 & ~n323 ;
  assign n325 = n155 & n237 ;
  assign n326 = n325 ^ x0 ;
  assign n327 = n326 ^ n325 ;
  assign n328 = n327 ^ n324 ;
  assign n329 = n268 ^ x9 ;
  assign n330 = n73 ^ x9 ;
  assign n331 = n330 ^ x9 ;
  assign n332 = n329 & ~n331 ;
  assign n333 = n332 ^ x9 ;
  assign n334 = ~n74 & n333 ;
  assign n335 = n334 ^ x9 ;
  assign n336 = n335 ^ n140 ;
  assign n337 = n336 ^ n335 ;
  assign n338 = n335 ^ n235 ;
  assign n339 = n338 ^ n335 ;
  assign n340 = n337 & n339 ;
  assign n341 = n340 ^ n335 ;
  assign n342 = ~x5 & n341 ;
  assign n343 = n342 ^ n335 ;
  assign n344 = n343 ^ x6 ;
  assign n345 = n343 & ~n344 ;
  assign n346 = n345 ^ n325 ;
  assign n347 = n346 ^ n343 ;
  assign n348 = n328 & n347 ;
  assign n349 = n348 ^ n345 ;
  assign n350 = n349 ^ n343 ;
  assign n351 = ~n324 & n350 ;
  assign n352 = n351 ^ n324 ;
  assign n353 = ~x4 & n352 ;
  assign n354 = n88 & ~n155 ;
  assign n355 = ~n222 & ~n354 ;
  assign n356 = x4 & n355 ;
  assign n357 = x6 & ~n122 ;
  assign n358 = n140 & ~n357 ;
  assign n359 = n358 ^ x0 ;
  assign n360 = n359 ^ n358 ;
  assign n361 = n360 ^ n356 ;
  assign n362 = n91 ^ x6 ;
  assign n363 = n155 ^ x3 ;
  assign n364 = n363 ^ n155 ;
  assign n365 = n235 ^ n155 ;
  assign n366 = n364 & n365 ;
  assign n367 = n366 ^ n155 ;
  assign n368 = n367 ^ n91 ;
  assign n369 = n362 & n368 ;
  assign n370 = n369 ^ n366 ;
  assign n371 = n370 ^ n155 ;
  assign n372 = n371 ^ x6 ;
  assign n373 = n91 & n372 ;
  assign n374 = n373 ^ n91 ;
  assign n375 = n36 & n56 ;
  assign n376 = ~x6 & n375 ;
  assign n377 = n376 ^ n374 ;
  assign n378 = ~n374 & n377 ;
  assign n379 = n378 ^ n358 ;
  assign n380 = n379 ^ n374 ;
  assign n381 = ~n361 & n380 ;
  assign n382 = n381 ^ n378 ;
  assign n383 = n382 ^ n374 ;
  assign n384 = n356 & ~n383 ;
  assign n385 = n384 ^ n356 ;
  assign n386 = ~n353 & ~n385 ;
  assign n387 = n386 ^ n313 ;
  assign n388 = n315 & n387 ;
  assign n389 = n388 ^ n313 ;
  assign n390 = ~n224 & n389 ;
  assign n391 = n390 ^ n219 ;
  assign n392 = n221 & n391 ;
  assign n393 = n392 ^ n219 ;
  assign n394 = ~n47 & n393 ;
  assign y0 = ~n394 ;
endmodule
