module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 ;
  assign n17 = ~x3 & x4 ;
  assign n18 = x1 ^ x0 ;
  assign n19 = ~x8 & ~x15 ;
  assign n20 = n19 ^ x14 ;
  assign n21 = n20 ^ x13 ;
  assign n22 = n19 ^ x13 ;
  assign n23 = ~x11 & ~x12 ;
  assign n24 = x10 ^ x9 ;
  assign n25 = n24 ^ x8 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = x15 ^ x9 ;
  assign n28 = ~x8 & n27 ;
  assign n29 = n28 ^ x15 ;
  assign n30 = ~n26 & ~n29 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n31 ^ x15 ;
  assign n33 = n32 ^ x8 ;
  assign n34 = n23 & n33 ;
  assign n35 = n34 ^ x13 ;
  assign n36 = x13 & n35 ;
  assign n37 = n36 ^ x13 ;
  assign n38 = ~n22 & n37 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n39 ^ x13 ;
  assign n41 = n40 ^ n34 ;
  assign n42 = ~n21 & n41 ;
  assign n43 = ~x7 & ~n42 ;
  assign n44 = ~x2 & ~x5 ;
  assign n45 = ~n43 & n44 ;
  assign n46 = x1 & ~n45 ;
  assign n47 = n18 & n46 ;
  assign n48 = n47 ^ n18 ;
  assign n49 = n17 & n48 ;
  assign y0 = n49 ;
endmodule
