module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 ;
  output y0 ;
  wire n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 ;
  assign n26 = ~x6 & ~x23 ;
  assign n27 = ~x8 & n26 ;
  assign n28 = ~x7 & ~x9 ;
  assign n29 = ~x1 & ~x2 ;
  assign n37 = ~x0 & ~x3 ;
  assign n31 = ~x4 & ~x5 ;
  assign n38 = x4 & x5 ;
  assign n39 = ~x3 & ~n38 ;
  assign n40 = ~n31 & ~n39 ;
  assign n41 = ~n37 & ~n40 ;
  assign n30 = x0 & ~x16 ;
  assign n32 = ~x3 & n31 ;
  assign n33 = x13 & ~x14 ;
  assign n34 = ~x15 & n33 ;
  assign n35 = n32 & n34 ;
  assign n36 = n30 & n35 ;
  assign n42 = n41 ^ n36 ;
  assign n43 = n42 ^ x17 ;
  assign n54 = n43 ^ n42 ;
  assign n44 = ~x13 & x14 ;
  assign n45 = x15 & x17 ;
  assign n46 = x16 & n45 ;
  assign n47 = n44 & n46 ;
  assign n48 = n47 ^ n43 ;
  assign n49 = n48 ^ n42 ;
  assign n50 = n43 ^ n36 ;
  assign n51 = n50 ^ n47 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = ~n49 & ~n52 ;
  assign n55 = n54 ^ n53 ;
  assign n56 = n55 ^ n49 ;
  assign n57 = ~x15 & ~x16 ;
  assign n58 = x13 & n57 ;
  assign n59 = x14 & n58 ;
  assign n60 = n59 ^ n42 ;
  assign n61 = n53 ^ n49 ;
  assign n62 = ~n60 & ~n61 ;
  assign n63 = n62 ^ n42 ;
  assign n64 = ~n56 & n63 ;
  assign n65 = n64 ^ n42 ;
  assign n66 = n65 ^ n41 ;
  assign n67 = n66 ^ n42 ;
  assign n68 = n29 & n67 ;
  assign n69 = ~x1 & n58 ;
  assign n70 = ~n47 & ~n69 ;
  assign n71 = ~x2 & n39 ;
  assign n72 = ~n70 & ~n71 ;
  assign n73 = x24 & n31 ;
  assign n74 = ~x1 & ~n73 ;
  assign n75 = n44 & ~n74 ;
  assign n76 = n44 & n57 ;
  assign n77 = ~n33 & ~n76 ;
  assign n78 = ~n75 & n77 ;
  assign n79 = ~x3 & n29 ;
  assign n80 = n73 & n79 ;
  assign n81 = n80 ^ n46 ;
  assign n82 = n81 ^ n74 ;
  assign n83 = n76 ^ n44 ;
  assign n84 = n46 & ~n83 ;
  assign n85 = n84 ^ n76 ;
  assign n86 = ~n82 & n85 ;
  assign n87 = n86 ^ n84 ;
  assign n88 = n87 ^ n76 ;
  assign n89 = n88 ^ n46 ;
  assign n90 = ~n74 & n89 ;
  assign n91 = ~n78 & n90 ;
  assign n92 = x17 ^ x14 ;
  assign n93 = ~n74 & n92 ;
  assign n95 = x14 & x17 ;
  assign n96 = x5 & ~n95 ;
  assign n97 = ~x4 & ~n96 ;
  assign n94 = ~x1 & ~n92 ;
  assign n98 = n97 ^ n94 ;
  assign n99 = n98 ^ n94 ;
  assign n100 = ~x1 & ~x5 ;
  assign n101 = ~x3 & ~n100 ;
  assign n102 = ~x2 & n101 ;
  assign n103 = n102 ^ n94 ;
  assign n104 = n99 & n103 ;
  assign n105 = n104 ^ n94 ;
  assign n106 = ~n93 & ~n105 ;
  assign n107 = n58 & ~n106 ;
  assign n108 = ~n91 & ~n107 ;
  assign n109 = ~n72 & n108 ;
  assign n110 = ~x0 & ~n109 ;
  assign n111 = ~n68 & ~n110 ;
  assign n112 = ~x10 & ~n111 ;
  assign n113 = ~x0 & x10 ;
  assign n114 = n80 & n113 ;
  assign n115 = x22 ^ x13 ;
  assign n116 = n115 ^ x22 ;
  assign n117 = n116 ^ n114 ;
  assign n118 = ~x20 & x21 ;
  assign n119 = x19 & n118 ;
  assign n120 = n119 ^ x18 ;
  assign n121 = n119 & n120 ;
  assign n122 = n121 ^ x22 ;
  assign n123 = n122 ^ n119 ;
  assign n124 = ~n117 & ~n123 ;
  assign n125 = n124 ^ n121 ;
  assign n126 = n125 ^ n119 ;
  assign n127 = n114 & n126 ;
  assign n128 = n127 ^ n114 ;
  assign n129 = ~n112 & ~n128 ;
  assign n130 = x11 & ~n129 ;
  assign n131 = x14 ^ x13 ;
  assign n132 = ~x0 & n131 ;
  assign n133 = x16 & ~n132 ;
  assign n134 = x10 & x15 ;
  assign n135 = ~x11 & ~x17 ;
  assign n136 = n134 & n135 ;
  assign n137 = ~x13 & ~x14 ;
  assign n138 = ~x16 & ~n137 ;
  assign n139 = n31 & ~n138 ;
  assign n140 = n136 & n139 ;
  assign n141 = x16 ^ x3 ;
  assign n142 = n141 ^ x16 ;
  assign n143 = x24 ^ x16 ;
  assign n144 = ~n142 & n143 ;
  assign n145 = n144 ^ x16 ;
  assign n146 = ~x0 & ~n145 ;
  assign n147 = n146 ^ x3 ;
  assign n148 = n29 & ~n147 ;
  assign n149 = n140 & n148 ;
  assign n150 = ~n133 & n149 ;
  assign n151 = ~n130 & ~n150 ;
  assign n154 = n151 ^ n114 ;
  assign n155 = n154 ^ n151 ;
  assign n152 = n151 ^ n34 ;
  assign n153 = n152 ^ n151 ;
  assign n156 = n155 ^ n153 ;
  assign n157 = n151 ^ x11 ;
  assign n158 = n157 ^ n151 ;
  assign n159 = n158 ^ n155 ;
  assign n160 = n155 & n159 ;
  assign n161 = n160 ^ n155 ;
  assign n162 = n156 & n161 ;
  assign n163 = n162 ^ n160 ;
  assign n164 = n163 ^ n151 ;
  assign n165 = n164 ^ n155 ;
  assign n166 = x12 & ~n165 ;
  assign n167 = n166 ^ n151 ;
  assign n168 = n28 & ~n167 ;
  assign n169 = n27 & n168 ;
  assign y0 = n169 ;
endmodule
