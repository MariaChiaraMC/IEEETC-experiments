module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n13 = x11 ^ x4 ;
  assign n14 = x0 & x7 ;
  assign n15 = x1 & x8 ;
  assign n16 = n14 & n15 ;
  assign n17 = x9 & n16 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = ~x2 & ~x6 ;
  assign n20 = ~x3 & x5 ;
  assign n21 = n19 & n20 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = x5 & x10 ;
  assign n25 = x6 & ~n24 ;
  assign n26 = x2 & x3 ;
  assign n27 = n25 & n26 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = n23 & n28 ;
  assign n30 = n29 ^ n21 ;
  assign n31 = n30 ^ n13 ;
  assign n32 = n18 & n31 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ n21 ;
  assign n35 = n34 ^ n17 ;
  assign n36 = n13 & n35 ;
  assign n37 = n36 ^ n13 ;
  assign y0 = n37 ;
endmodule
