module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 ;
  assign n17 = ~x9 & ~x10 ;
  assign n18 = ~x12 & ~x13 ;
  assign n19 = ~n17 & n18 ;
  assign n20 = ~x8 & x15 ;
  assign n21 = ~x11 & ~x14 ;
  assign n22 = n20 & n21 ;
  assign n23 = n19 & n22 ;
  assign n24 = n23 ^ x6 ;
  assign n25 = n24 ^ x6 ;
  assign n26 = n25 ^ x0 ;
  assign n30 = ~x4 & x5 ;
  assign n31 = ~x7 & ~n30 ;
  assign n27 = x9 & x10 ;
  assign n28 = x5 & ~n27 ;
  assign n29 = x7 & ~n28 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = ~x6 & ~n32 ;
  assign n34 = n33 ^ n29 ;
  assign n35 = ~n26 & ~n34 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = n36 ^ n29 ;
  assign n38 = n37 ^ x6 ;
  assign n39 = ~x0 & n38 ;
  assign n40 = n39 ^ x6 ;
  assign y0 = ~n40 ;
endmodule
