module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 ;
  assign n16 = x5 ^ x4 ;
  assign n26 = x5 ^ x3 ;
  assign n18 = x5 ^ x2 ;
  assign n19 = n18 ^ x5 ;
  assign n27 = n26 ^ n19 ;
  assign n28 = n27 ^ x5 ;
  assign n17 = n16 ^ x1 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n20 ^ n16 ;
  assign n29 = n28 ^ n21 ;
  assign n30 = n29 ^ n16 ;
  assign n31 = ~n16 & n30 ;
  assign n32 = n31 ^ n19 ;
  assign n33 = n32 ^ n21 ;
  assign n34 = n33 ^ n16 ;
  assign n35 = n34 ^ x5 ;
  assign n36 = n21 ^ n16 ;
  assign n37 = n36 ^ x5 ;
  assign n38 = ~n33 & n37 ;
  assign n39 = n38 ^ n19 ;
  assign n40 = n39 ^ n21 ;
  assign n41 = n40 ^ n16 ;
  assign n42 = n41 ^ x5 ;
  assign n43 = ~n35 & ~n42 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ n16 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n23 & ~n24 ;
  assign n44 = n43 ^ n25 ;
  assign n45 = n44 ^ n31 ;
  assign n46 = n45 ^ n19 ;
  assign n47 = n46 ^ n21 ;
  assign n48 = n47 ^ n16 ;
  assign n49 = n48 ^ x5 ;
  assign n50 = n49 ^ x4 ;
  assign n51 = ~x4 & x5 ;
  assign n52 = ~x2 & n51 ;
  assign n53 = n26 ^ x5 ;
  assign n55 = ~x8 & ~x12 ;
  assign n56 = x1 & ~x13 ;
  assign n57 = n55 & n56 ;
  assign n58 = ~x10 & n57 ;
  assign n54 = ~x1 & x11 ;
  assign n59 = n58 ^ n54 ;
  assign n60 = n59 ^ n54 ;
  assign n61 = ~x7 & ~x9 ;
  assign n62 = x2 & ~x14 ;
  assign n63 = ~n61 & n62 ;
  assign n64 = n63 ^ n54 ;
  assign n65 = n64 ^ n54 ;
  assign n66 = n60 & n65 ;
  assign n67 = n66 ^ n54 ;
  assign n68 = x4 & n67 ;
  assign n69 = n68 ^ n54 ;
  assign n70 = n69 ^ x5 ;
  assign n71 = n53 & ~n70 ;
  assign n72 = n71 ^ x5 ;
  assign n73 = ~x1 & ~x5 ;
  assign n74 = n73 ^ n52 ;
  assign n75 = ~n72 & ~n74 ;
  assign n76 = n75 ^ n73 ;
  assign n77 = ~n52 & n76 ;
  assign n78 = n77 ^ n52 ;
  assign n79 = n78 ^ x6 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = ~x3 & x4 ;
  assign n82 = x1 & ~x5 ;
  assign n83 = ~x2 & n82 ;
  assign n84 = x3 & n51 ;
  assign n85 = ~n83 & ~n84 ;
  assign n86 = ~n81 & n85 ;
  assign n87 = n86 ^ n78 ;
  assign n88 = ~n80 & ~n87 ;
  assign n89 = n88 ^ n78 ;
  assign n90 = n50 & ~n89 ;
  assign n91 = ~x0 & ~n90 ;
  assign y0 = n91 ;
endmodule
