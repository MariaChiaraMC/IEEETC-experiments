module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 ;
  assign n11 = x4 & x7 ;
  assign n87 = x2 & ~n11 ;
  assign n86 = ~x4 & ~x7 ;
  assign n133 = ~x1 & ~x3 ;
  assign n134 = ~n86 & n133 ;
  assign n135 = ~n87 & n134 ;
  assign n10 = x1 & x2 ;
  assign n16 = x4 & ~x7 ;
  assign n136 = x3 & n16 ;
  assign n137 = n10 & n136 ;
  assign n138 = ~n135 & ~n137 ;
  assign n139 = x0 & ~n138 ;
  assign n140 = x1 & x3 ;
  assign n141 = ~x2 & n140 ;
  assign n142 = n141 ^ x7 ;
  assign n143 = n142 ^ x4 ;
  assign n144 = ~x1 & x2 ;
  assign n145 = ~x0 & ~x3 ;
  assign n146 = n144 & n145 ;
  assign n147 = n146 ^ x0 ;
  assign n148 = ~x7 & n147 ;
  assign n149 = n148 ^ x0 ;
  assign n150 = n143 & ~n149 ;
  assign n151 = n150 ^ n148 ;
  assign n152 = n151 ^ x0 ;
  assign n153 = n152 ^ x7 ;
  assign n154 = ~x4 & n153 ;
  assign n155 = ~n139 & ~n154 ;
  assign n119 = ~x0 & ~x2 ;
  assign n120 = n86 & n119 ;
  assign n72 = x2 & x3 ;
  assign n121 = x0 & x7 ;
  assign n122 = n72 & n121 ;
  assign n123 = x4 & n122 ;
  assign n124 = ~n120 & ~n123 ;
  assign n125 = ~x1 & ~n124 ;
  assign n17 = x0 & ~x1 ;
  assign n92 = ~x4 & x7 ;
  assign n126 = ~n17 & n92 ;
  assign n127 = x3 ^ x2 ;
  assign n128 = n126 & ~n127 ;
  assign n129 = ~n10 & n128 ;
  assign n130 = ~n125 & ~n129 ;
  assign n9 = x5 ^ x3 ;
  assign n12 = n10 & n11 ;
  assign n13 = n12 ^ x5 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n14 ^ n9 ;
  assign n18 = n17 ^ n16 ;
  assign n19 = n16 & n18 ;
  assign n20 = n19 ^ n12 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = ~n15 & n21 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = n23 ^ n16 ;
  assign n25 = n9 & n24 ;
  assign n26 = x5 ^ x1 ;
  assign n27 = n26 ^ x7 ;
  assign n31 = n27 ^ x3 ;
  assign n32 = n31 ^ n27 ;
  assign n33 = n32 ^ x5 ;
  assign n35 = n33 ^ x5 ;
  assign n28 = x5 ^ x4 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ x5 ;
  assign n36 = n35 ^ n30 ;
  assign n34 = ~n30 & n33 ;
  assign n37 = n36 ^ n34 ;
  assign n41 = x5 ^ x2 ;
  assign n42 = n41 ^ n31 ;
  assign n38 = n27 ^ x7 ;
  assign n39 = n38 ^ n31 ;
  assign n40 = n39 ^ n27 ;
  assign n43 = n42 ^ n40 ;
  assign n44 = n43 ^ n31 ;
  assign n45 = n44 ^ x5 ;
  assign n46 = n45 ^ n30 ;
  assign n47 = n40 ^ n30 ;
  assign n48 = ~n46 & n47 ;
  assign n49 = n48 ^ n40 ;
  assign n50 = n49 ^ n33 ;
  assign n51 = n50 ^ n45 ;
  assign n52 = n45 ^ n33 ;
  assign n53 = n52 ^ n36 ;
  assign n54 = n45 ^ n27 ;
  assign n55 = n54 ^ n36 ;
  assign n56 = ~n53 & n55 ;
  assign n57 = n56 ^ n40 ;
  assign n58 = n57 ^ n27 ;
  assign n59 = n58 ^ n33 ;
  assign n60 = ~n51 & n59 ;
  assign n61 = n60 ^ n27 ;
  assign n62 = ~n37 & ~n61 ;
  assign n63 = n62 ^ n34 ;
  assign n64 = n63 ^ n60 ;
  assign n65 = n64 ^ n36 ;
  assign n66 = n65 ^ n27 ;
  assign n67 = n66 ^ x0 ;
  assign n68 = n67 ^ n66 ;
  assign n83 = ~x2 & n11 ;
  assign n84 = ~x3 & x5 ;
  assign n85 = n83 & n84 ;
  assign n88 = ~n86 & n87 ;
  assign n89 = x3 & ~n88 ;
  assign n90 = ~x2 & ~x5 ;
  assign n91 = n86 & n90 ;
  assign n93 = n92 ^ x2 ;
  assign n94 = ~x2 & ~n41 ;
  assign n95 = n94 ^ x2 ;
  assign n96 = n93 & ~n95 ;
  assign n97 = n96 ^ n94 ;
  assign n98 = n97 ^ x2 ;
  assign n99 = n98 ^ x5 ;
  assign n100 = ~n91 & ~n99 ;
  assign n101 = n100 ^ n91 ;
  assign n102 = n89 & n101 ;
  assign n103 = ~n85 & ~n102 ;
  assign n69 = ~x2 & ~x3 ;
  assign n70 = ~x7 & n69 ;
  assign n71 = n70 ^ x5 ;
  assign n73 = n72 ^ n70 ;
  assign n74 = n72 ^ n28 ;
  assign n75 = ~n72 & n74 ;
  assign n76 = n75 ^ n72 ;
  assign n77 = n73 & ~n76 ;
  assign n78 = n77 ^ n75 ;
  assign n79 = n78 ^ n72 ;
  assign n80 = n79 ^ n28 ;
  assign n81 = ~n71 & n80 ;
  assign n82 = n81 ^ n70 ;
  assign n104 = n103 ^ n82 ;
  assign n105 = n82 ^ x7 ;
  assign n106 = n82 ^ x1 ;
  assign n107 = n82 & ~n106 ;
  assign n108 = n107 ^ n82 ;
  assign n109 = n105 & n108 ;
  assign n110 = n109 ^ n107 ;
  assign n111 = n110 ^ n82 ;
  assign n112 = n111 ^ x1 ;
  assign n113 = ~n104 & ~n112 ;
  assign n114 = n113 ^ n82 ;
  assign n115 = n114 ^ n66 ;
  assign n116 = ~n68 & ~n115 ;
  assign n117 = n116 ^ n66 ;
  assign n118 = ~n25 & n117 ;
  assign n131 = n130 ^ n118 ;
  assign n132 = n131 ^ n130 ;
  assign n156 = n155 ^ n132 ;
  assign n157 = n156 ^ n131 ;
  assign n158 = n131 ^ x5 ;
  assign n159 = n158 ^ n131 ;
  assign n160 = n157 & ~n159 ;
  assign n161 = n160 ^ n131 ;
  assign n162 = ~x6 & n161 ;
  assign n163 = n162 ^ n118 ;
  assign y0 = ~n163 ;
endmodule
