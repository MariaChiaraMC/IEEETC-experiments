module top( x0 , x1 , x2 , x3 , x4 , y0 );
  input x0 , x1 , x2 , x3 , x4 ;
  output y0 ;
  wire n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n9 = x3 ^ x2 ;
  assign n6 = x4 ^ x1 ;
  assign n7 = n6 ^ x0 ;
  assign n8 = n7 ^ x2 ;
  assign n10 = n9 ^ n8 ;
  assign n13 = n7 ^ x0 ;
  assign n11 = x1 ^ x0 ;
  assign n12 = n11 ^ n8 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n10 & n14 ;
  assign n16 = n15 ^ n7 ;
  assign n17 = n16 ^ n11 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = n12 ^ n9 ;
  assign n20 = n16 & n19 ;
  assign n21 = n20 ^ n7 ;
  assign n22 = n21 ^ n8 ;
  assign n23 = n22 ^ n9 ;
  assign n24 = n18 & n23 ;
  assign y0 = n24 ;
endmodule
