module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 ;
  assign n7 = x3 ^ x2 ;
  assign n8 = n7 ^ x2 ;
  assign n9 = x0 & x1 ;
  assign n10 = n9 ^ x2 ;
  assign n11 = ~n8 & n10 ;
  assign n12 = n11 ^ x2 ;
  assign n13 = ~x4 & ~n12 ;
  assign n15 = ~x0 & x5 ;
  assign n16 = ~x1 & ~n15 ;
  assign n14 = x0 & x2 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = n14 ^ x5 ;
  assign n19 = n18 ^ x3 ;
  assign n20 = n19 ^ n14 ;
  assign n21 = ~n17 & ~n20 ;
  assign n22 = n21 ^ n14 ;
  assign n23 = ~x3 & n14 ;
  assign n24 = n23 ^ x4 ;
  assign n25 = n22 & n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = x4 & n26 ;
  assign n28 = n27 ^ x4 ;
  assign n29 = ~n13 & ~n28 ;
  assign n30 = x5 ^ x3 ;
  assign n31 = ~x0 & n30 ;
  assign n32 = n31 ^ x3 ;
  assign n33 = ~x1 & n32 ;
  assign n34 = ~x3 & ~x5 ;
  assign n35 = ~x4 & n34 ;
  assign n36 = ~n33 & ~n35 ;
  assign n37 = n36 ^ x0 ;
  assign n38 = n37 ^ x2 ;
  assign n47 = n38 ^ n37 ;
  assign n39 = x1 & ~x5 ;
  assign n40 = x3 & n39 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n41 ^ n37 ;
  assign n43 = n38 ^ n36 ;
  assign n44 = n43 ^ n40 ;
  assign n45 = n44 ^ n42 ;
  assign n46 = n42 & n45 ;
  assign n48 = n47 ^ n46 ;
  assign n49 = n48 ^ n42 ;
  assign n50 = ~x4 & x5 ;
  assign n51 = n50 ^ n37 ;
  assign n52 = n46 ^ n42 ;
  assign n53 = ~n51 & n52 ;
  assign n54 = n53 ^ n37 ;
  assign n55 = ~n49 & n54 ;
  assign n56 = n55 ^ n37 ;
  assign n57 = n56 ^ x0 ;
  assign n58 = n57 ^ n37 ;
  assign n59 = ~n29 & n58 ;
  assign y0 = ~n59 ;
endmodule
