module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n8 = x3 & x4 ;
  assign n9 = ~x2 & ~n8 ;
  assign n10 = ~x1 & ~n9 ;
  assign n12 = ~x3 & ~x5 ;
  assign n13 = ~x4 & n12 ;
  assign n11 = x2 ^ x0 ;
  assign n14 = n13 ^ n11 ;
  assign n15 = n14 ^ n11 ;
  assign n16 = n11 ^ x0 ;
  assign n17 = n15 & n16 ;
  assign n18 = n17 ^ n11 ;
  assign n19 = x6 & ~n11 ;
  assign n20 = n19 ^ n10 ;
  assign n21 = ~n18 & ~n20 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = ~n10 & n22 ;
  assign n24 = n23 ^ n10 ;
  assign y0 = n24 ;
endmodule
