module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 ;
  assign n9 = x2 & x3 ;
  assign n10 = n9 ^ x1 ;
  assign n11 = n10 ^ n9 ;
  assign n12 = n11 ^ x0 ;
  assign n38 = x4 & ~x5 ;
  assign n15 = x4 ^ x2 ;
  assign n16 = n15 ^ x6 ;
  assign n13 = x5 ^ x4 ;
  assign n14 = n13 ^ x6 ;
  assign n17 = n16 ^ n14 ;
  assign n18 = n17 ^ x4 ;
  assign n19 = x6 ^ x4 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = n20 ^ n16 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = n22 ^ x7 ;
  assign n24 = n23 ^ n14 ;
  assign n25 = ~n16 & ~n24 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = n26 ^ n18 ;
  assign n28 = n22 ^ n16 ;
  assign n29 = n28 ^ n18 ;
  assign n30 = x4 & n29 ;
  assign n31 = n30 ^ n16 ;
  assign n32 = ~n27 & ~n31 ;
  assign n33 = ~n18 & n32 ;
  assign n34 = n33 ^ n25 ;
  assign n35 = n34 ^ n30 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = ~x3 & ~n36 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = ~n9 & ~n39 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n12 & n41 ;
  assign n43 = n42 ^ n40 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = n44 ^ n9 ;
  assign n46 = ~x0 & ~n45 ;
  assign y0 = n46 ;
endmodule
