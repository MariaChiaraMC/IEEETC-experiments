module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 ;
  assign n249 = ~x5 & x9 ;
  assign n83 = x13 & x14 ;
  assign n18 = ~x15 & ~x16 ;
  assign n225 = x2 & n18 ;
  assign n250 = n83 & n225 ;
  assign n251 = ~x8 & n250 ;
  assign n49 = x15 & x16 ;
  assign n148 = x2 & n49 ;
  assign n232 = ~x11 & ~x13 ;
  assign n252 = n148 & n232 ;
  assign n125 = x13 & n49 ;
  assign n104 = x3 & x8 ;
  assign n105 = ~x2 & n104 ;
  assign n184 = ~x8 & x14 ;
  assign n253 = ~n105 & ~n184 ;
  assign n254 = n125 & ~n253 ;
  assign n255 = ~x4 & n254 ;
  assign n256 = ~n252 & ~n255 ;
  assign n257 = ~n251 & n256 ;
  assign n258 = n249 & ~n257 ;
  assign n149 = x10 & x11 ;
  assign n150 = ~x13 & n149 ;
  assign n259 = n148 & n150 ;
  assign n160 = ~x8 & n49 ;
  assign n161 = ~x13 & n160 ;
  assign n19 = x14 & n18 ;
  assign n260 = x8 & n19 ;
  assign n261 = ~n161 & ~n260 ;
  assign n262 = ~x4 & ~n261 ;
  assign n263 = ~x5 & n184 ;
  assign n264 = n18 & n263 ;
  assign n265 = ~n262 & ~n264 ;
  assign n266 = ~n149 & ~n265 ;
  assign n267 = x2 & n266 ;
  assign n268 = ~x5 & x13 ;
  assign n269 = ~x4 & x14 ;
  assign n270 = n160 & n269 ;
  assign n271 = n18 & n149 ;
  assign n272 = x14 & n271 ;
  assign n273 = ~n270 & ~n272 ;
  assign n274 = n273 ^ x2 ;
  assign n275 = n274 ^ n273 ;
  assign n276 = n275 ^ n268 ;
  assign n199 = ~x10 & n49 ;
  assign n277 = ~n160 & ~n199 ;
  assign n278 = n269 & ~n277 ;
  assign n279 = ~x10 & x14 ;
  assign n280 = ~x4 & n49 ;
  assign n281 = ~n199 & ~n280 ;
  assign n282 = ~n279 & ~n281 ;
  assign n283 = n104 & n282 ;
  assign n284 = n283 ^ n278 ;
  assign n285 = ~n278 & n284 ;
  assign n286 = n285 ^ n273 ;
  assign n287 = n286 ^ n278 ;
  assign n288 = ~n276 & ~n287 ;
  assign n289 = n288 ^ n285 ;
  assign n290 = n289 ^ n278 ;
  assign n291 = n268 & ~n290 ;
  assign n292 = n291 ^ n268 ;
  assign n293 = ~n267 & ~n292 ;
  assign n294 = ~n259 & n293 ;
  assign n295 = ~x9 & ~n294 ;
  assign n296 = ~n258 & ~n295 ;
  assign n297 = x6 & ~n296 ;
  assign n25 = x5 & ~x6 ;
  assign n92 = ~x7 & n25 ;
  assign n113 = ~x4 & x6 ;
  assign n298 = ~n92 & ~n113 ;
  assign n299 = x2 & ~x9 ;
  assign n300 = ~n149 & n299 ;
  assign n301 = ~x9 & n279 ;
  assign n302 = ~x2 & ~x3 ;
  assign n303 = x13 & n302 ;
  assign n304 = ~n301 & n303 ;
  assign n305 = ~n300 & ~n304 ;
  assign n306 = n49 & ~n305 ;
  assign n108 = n18 & n83 ;
  assign n307 = x2 & x9 ;
  assign n308 = ~x11 & n307 ;
  assign n309 = n108 & n308 ;
  assign n310 = ~n306 & ~n309 ;
  assign n311 = x8 & ~n310 ;
  assign n155 = ~n19 & ~n49 ;
  assign n21 = ~x8 & x13 ;
  assign n219 = x11 & ~n21 ;
  assign n312 = n219 & n307 ;
  assign n313 = ~n155 & n312 ;
  assign n314 = ~n311 & ~n313 ;
  assign n315 = ~n298 & ~n314 ;
  assign n316 = x4 & x9 ;
  assign n131 = ~x7 & x8 ;
  assign n132 = ~x6 & n131 ;
  assign n109 = ~x2 & n108 ;
  assign n317 = ~n109 & ~n252 ;
  assign n318 = n132 & ~n317 ;
  assign n319 = n316 & n318 ;
  assign n320 = ~n315 & ~n319 ;
  assign n321 = ~n297 & n320 ;
  assign n20 = x2 & x6 ;
  assign n22 = ~x4 & x5 ;
  assign n23 = n21 & n22 ;
  assign n24 = n20 & ~n23 ;
  assign n32 = x6 & ~x13 ;
  assign n26 = ~x7 & ~x8 ;
  assign n27 = x4 & ~x6 ;
  assign n28 = ~n26 & n27 ;
  assign n29 = ~n25 & ~n28 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n33 ^ n29 ;
  assign n30 = n29 ^ n22 ;
  assign n31 = n30 ^ n29 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = n29 ^ x3 ;
  assign n37 = n36 ^ n29 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = n34 & n38 ;
  assign n40 = n39 ^ n34 ;
  assign n41 = n35 & n40 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = n42 ^ n29 ;
  assign n44 = n43 ^ n34 ;
  assign n45 = ~x2 & ~n44 ;
  assign n46 = n45 ^ n29 ;
  assign n47 = ~n24 & n46 ;
  assign n48 = n19 & ~n47 ;
  assign n50 = x4 & x5 ;
  assign n51 = x6 & ~n21 ;
  assign n52 = ~x5 & n28 ;
  assign n53 = ~n51 & ~n52 ;
  assign n54 = ~n50 & ~n53 ;
  assign n55 = x2 & n54 ;
  assign n56 = ~x6 & x8 ;
  assign n57 = ~n32 & ~n56 ;
  assign n58 = ~x2 & x3 ;
  assign n59 = ~x14 & n58 ;
  assign n60 = x5 & ~x7 ;
  assign n61 = ~x4 & n60 ;
  assign n62 = n59 & n61 ;
  assign n63 = ~n57 & n62 ;
  assign n64 = x2 & x5 ;
  assign n65 = ~x6 & x7 ;
  assign n66 = ~n56 & ~n65 ;
  assign n67 = x4 & x6 ;
  assign n68 = n66 & ~n67 ;
  assign n69 = n64 & ~n68 ;
  assign n70 = ~n63 & ~n69 ;
  assign n71 = ~n55 & n70 ;
  assign n72 = x4 & ~x5 ;
  assign n73 = ~x6 & ~x7 ;
  assign n74 = n72 & n73 ;
  assign n75 = x5 & x6 ;
  assign n76 = ~x4 & n75 ;
  assign n77 = ~n74 & ~n76 ;
  assign n78 = ~x5 & ~x14 ;
  assign n79 = n20 & n78 ;
  assign n80 = x4 & n79 ;
  assign n81 = n77 & ~n80 ;
  assign n82 = n21 & ~n81 ;
  assign n84 = ~x4 & x8 ;
  assign n85 = ~x3 & n84 ;
  assign n86 = ~n65 & ~n85 ;
  assign n87 = ~x2 & x5 ;
  assign n88 = ~x3 & ~x6 ;
  assign n89 = n87 & ~n88 ;
  assign n90 = ~n86 & n89 ;
  assign n91 = ~x5 & x6 ;
  assign n93 = ~n91 & ~n92 ;
  assign n94 = x4 & ~x8 ;
  assign n95 = x2 & x8 ;
  assign n96 = ~n94 & ~n95 ;
  assign n97 = ~n93 & n96 ;
  assign n98 = ~n90 & ~n97 ;
  assign n99 = n83 & ~n98 ;
  assign n100 = ~n82 & ~n99 ;
  assign n101 = n71 & n100 ;
  assign n102 = n49 & ~n101 ;
  assign n103 = ~n48 & ~n102 ;
  assign n106 = n19 & n74 ;
  assign n107 = n105 & n106 ;
  assign n110 = x4 & x8 ;
  assign n111 = ~x7 & n110 ;
  assign n112 = n111 ^ x5 ;
  assign n114 = x8 & n113 ;
  assign n115 = ~n67 & ~n114 ;
  assign n116 = n115 ^ n88 ;
  assign n117 = n111 ^ n88 ;
  assign n118 = n117 ^ n88 ;
  assign n119 = n116 & ~n118 ;
  assign n120 = n119 ^ n88 ;
  assign n121 = n112 & n120 ;
  assign n122 = n121 ^ x5 ;
  assign n123 = n109 & n122 ;
  assign n124 = ~n107 & ~n123 ;
  assign n126 = ~n72 & ~n85 ;
  assign n127 = x6 & ~n126 ;
  assign n128 = x3 & ~x7 ;
  assign n129 = x3 & ~x4 ;
  assign n130 = ~n128 & ~n129 ;
  assign n133 = ~x3 & ~n132 ;
  assign n134 = n130 & ~n133 ;
  assign n135 = x5 & n134 ;
  assign n136 = ~n127 & ~n135 ;
  assign n137 = ~x14 & ~n136 ;
  assign n138 = x6 & n104 ;
  assign n139 = ~x5 & x14 ;
  assign n140 = ~n50 & ~n139 ;
  assign n141 = n138 & n140 ;
  assign n142 = ~n52 & ~n141 ;
  assign n143 = ~n137 & n142 ;
  assign n144 = ~x2 & ~n143 ;
  assign n145 = n125 & n144 ;
  assign n146 = n124 & ~n145 ;
  assign n147 = n103 & n146 ;
  assign n322 = n321 ^ n147 ;
  assign n323 = n322 ^ n147 ;
  assign n151 = ~x6 & n150 ;
  assign n152 = n148 & n151 ;
  assign n153 = n19 & n132 ;
  assign n154 = n58 & n153 ;
  assign n156 = x6 & ~x8 ;
  assign n157 = x2 & ~n156 ;
  assign n158 = ~n26 & n157 ;
  assign n159 = ~n155 & n158 ;
  assign n162 = n20 & n161 ;
  assign n163 = ~n159 & ~n162 ;
  assign n164 = ~n154 & n163 ;
  assign n165 = ~n149 & ~n164 ;
  assign n166 = ~n152 & ~n165 ;
  assign n167 = ~x5 & ~n166 ;
  assign n168 = ~x5 & n49 ;
  assign n169 = n26 & n168 ;
  assign n170 = x7 & n49 ;
  assign n171 = ~x5 & n170 ;
  assign n172 = n19 & n131 ;
  assign n173 = ~n171 & ~n172 ;
  assign n174 = n149 & ~n173 ;
  assign n175 = x2 & n174 ;
  assign n176 = ~n169 & ~n175 ;
  assign n177 = ~x6 & ~n176 ;
  assign n178 = n79 & n160 ;
  assign n180 = ~x10 & ~x14 ;
  assign n179 = x3 & n156 ;
  assign n181 = n180 ^ n179 ;
  assign n182 = n181 ^ n179 ;
  assign n183 = n182 ^ n66 ;
  assign n185 = n184 ^ x6 ;
  assign n186 = ~n184 & ~n185 ;
  assign n187 = n186 ^ n179 ;
  assign n188 = n187 ^ n184 ;
  assign n189 = ~n183 & ~n188 ;
  assign n190 = n189 ^ n186 ;
  assign n191 = n190 ^ n184 ;
  assign n192 = n66 & ~n191 ;
  assign n193 = n192 ^ n66 ;
  assign n194 = n168 & ~n193 ;
  assign n195 = n153 ^ x3 ;
  assign n196 = n153 ^ n149 ;
  assign n197 = n196 ^ n149 ;
  assign n198 = n197 ^ n195 ;
  assign n200 = n78 & n199 ;
  assign n201 = n200 ^ x6 ;
  assign n202 = x6 & n201 ;
  assign n203 = n202 ^ n149 ;
  assign n204 = n203 ^ x6 ;
  assign n205 = n198 & ~n204 ;
  assign n206 = n205 ^ n202 ;
  assign n207 = n206 ^ x6 ;
  assign n208 = ~n195 & n207 ;
  assign n209 = n208 ^ n153 ;
  assign n210 = ~n194 & ~n209 ;
  assign n211 = ~x2 & ~n210 ;
  assign n212 = ~n178 & ~n211 ;
  assign n213 = ~n177 & n212 ;
  assign n214 = x13 & ~n213 ;
  assign n215 = ~n167 & ~n214 ;
  assign n216 = n215 ^ x5 ;
  assign n217 = n216 ^ n215 ;
  assign n218 = ~x6 & ~n131 ;
  assign n220 = ~n218 & ~n219 ;
  assign n221 = n148 & ~n220 ;
  assign n222 = x6 & n184 ;
  assign n223 = n125 & ~n222 ;
  assign n224 = ~n157 & n223 ;
  assign n226 = x14 & n225 ;
  assign n227 = n21 ^ x11 ;
  assign n228 = n65 ^ x11 ;
  assign n229 = n228 ^ x11 ;
  assign n230 = ~n227 & ~n229 ;
  assign n231 = n230 ^ x11 ;
  assign n233 = n232 ^ n226 ;
  assign n234 = ~n231 & n233 ;
  assign n235 = n234 ^ n232 ;
  assign n236 = n226 & n235 ;
  assign n237 = n236 ^ n226 ;
  assign n238 = ~n224 & ~n237 ;
  assign n239 = ~n221 & n238 ;
  assign n240 = n239 ^ n215 ;
  assign n241 = n240 ^ n215 ;
  assign n242 = ~n217 & ~n241 ;
  assign n243 = n242 ^ n215 ;
  assign n244 = x9 & ~n243 ;
  assign n245 = n244 ^ n215 ;
  assign n246 = x4 & ~n245 ;
  assign n247 = n246 ^ n147 ;
  assign n248 = n247 ^ n147 ;
  assign n324 = n323 ^ n248 ;
  assign n325 = ~x9 & n199 ;
  assign n326 = ~n18 & ~n325 ;
  assign n327 = ~x3 & x6 ;
  assign n328 = x8 & n327 ;
  assign n329 = ~n326 & n328 ;
  assign n330 = n73 & ~n277 ;
  assign n331 = ~x9 & n330 ;
  assign n332 = ~n329 & ~n331 ;
  assign n333 = n269 & ~n332 ;
  assign n334 = ~x8 & n113 ;
  assign n335 = n49 & n334 ;
  assign n336 = x4 & n19 ;
  assign n337 = n327 & n336 ;
  assign n338 = x4 & x14 ;
  assign n339 = n132 & n338 ;
  assign n340 = n325 & n339 ;
  assign n341 = ~n337 & ~n340 ;
  assign n342 = ~n335 & n341 ;
  assign n343 = ~n333 & n342 ;
  assign n344 = x13 & ~n343 ;
  assign n345 = x9 & ~x11 ;
  assign n346 = ~x9 & n149 ;
  assign n347 = ~n128 & n346 ;
  assign n348 = ~n345 & ~n347 ;
  assign n349 = ~x13 & n18 ;
  assign n350 = ~x6 & n349 ;
  assign n351 = ~n348 & n350 ;
  assign n352 = ~x14 & n351 ;
  assign n353 = ~n344 & ~n352 ;
  assign n354 = n65 & n83 ;
  assign n355 = ~x7 & ~x14 ;
  assign n356 = ~x13 & ~n355 ;
  assign n357 = n51 & ~n356 ;
  assign n358 = n357 ^ n131 ;
  assign n359 = n358 ^ n357 ;
  assign n360 = ~x13 & x14 ;
  assign n361 = n360 ^ n357 ;
  assign n362 = n359 & ~n361 ;
  assign n363 = n362 ^ n357 ;
  assign n364 = ~n354 & ~n363 ;
  assign n365 = n280 & ~n364 ;
  assign n366 = n108 & n114 ;
  assign n367 = x14 & n49 ;
  assign n368 = x13 & n170 ;
  assign n369 = ~n367 & ~n368 ;
  assign n370 = n28 & ~n369 ;
  assign n371 = ~n366 & ~n370 ;
  assign n372 = ~n365 & n371 ;
  assign n373 = n372 ^ x9 ;
  assign n374 = n373 ^ n372 ;
  assign n375 = n374 ^ x3 ;
  assign n376 = x6 & x10 ;
  assign n377 = ~x14 & ~n376 ;
  assign n378 = n368 & n377 ;
  assign n379 = ~x6 & x10 ;
  assign n380 = ~n26 & n367 ;
  assign n381 = x11 & ~x13 ;
  assign n382 = n355 & n381 ;
  assign n383 = n18 & n382 ;
  assign n384 = ~n380 & ~n383 ;
  assign n385 = n379 & ~n384 ;
  assign n386 = n73 & ~n149 ;
  assign n387 = n260 & n386 ;
  assign n388 = x13 & n387 ;
  assign n389 = ~n385 & ~n388 ;
  assign n390 = ~n378 & n389 ;
  assign n391 = n390 ^ n199 ;
  assign n392 = n391 ^ x4 ;
  assign n399 = n392 ^ n391 ;
  assign n393 = n392 ^ n354 ;
  assign n394 = n393 ^ n391 ;
  assign n395 = n392 ^ n390 ;
  assign n396 = n395 ^ n354 ;
  assign n397 = n396 ^ n394 ;
  assign n398 = ~n394 & ~n397 ;
  assign n400 = n399 ^ n398 ;
  assign n401 = n400 ^ n394 ;
  assign n402 = n391 ^ n357 ;
  assign n403 = n398 ^ n394 ;
  assign n404 = n402 & ~n403 ;
  assign n405 = n404 ^ n391 ;
  assign n406 = ~n401 & ~n405 ;
  assign n407 = n406 ^ n391 ;
  assign n408 = n407 ^ n199 ;
  assign n409 = n408 ^ n391 ;
  assign n410 = n56 & n355 ;
  assign n411 = ~x7 & x14 ;
  assign n412 = n411 ^ n357 ;
  assign n413 = n412 ^ n357 ;
  assign n414 = x8 & x13 ;
  assign n415 = n414 ^ n357 ;
  assign n416 = n413 & n415 ;
  assign n417 = n416 ^ n357 ;
  assign n418 = ~n354 & ~n417 ;
  assign n419 = x10 & ~n418 ;
  assign n420 = ~n410 & ~n419 ;
  assign n421 = n49 & ~n420 ;
  assign n422 = x7 & n150 ;
  assign n423 = n19 & n51 ;
  assign n424 = ~n422 & n423 ;
  assign n425 = n349 & n355 ;
  assign n426 = n149 & n425 ;
  assign n427 = ~n424 & ~n426 ;
  assign n428 = ~n421 & n427 ;
  assign n429 = ~x4 & ~n428 ;
  assign n430 = n429 ^ n409 ;
  assign n431 = ~n409 & n430 ;
  assign n432 = n431 ^ n372 ;
  assign n433 = n432 ^ n409 ;
  assign n434 = ~n375 & ~n433 ;
  assign n435 = n434 ^ n431 ;
  assign n436 = n435 ^ n409 ;
  assign n437 = x3 & ~n436 ;
  assign n438 = n437 ^ x3 ;
  assign n439 = n353 & ~n438 ;
  assign n440 = ~x2 & ~n439 ;
  assign n441 = n73 & n251 ;
  assign n442 = ~n73 & ~n113 ;
  assign n443 = ~x11 & ~n49 ;
  assign n444 = n442 & ~n443 ;
  assign n445 = ~n155 & n444 ;
  assign n446 = ~x13 & n73 ;
  assign n447 = ~n156 & ~n446 ;
  assign n448 = n280 & ~n381 ;
  assign n449 = ~n447 & n448 ;
  assign n450 = x9 & ~n449 ;
  assign n451 = ~n445 & n450 ;
  assign n452 = x2 & ~n451 ;
  assign n453 = ~n441 & ~n452 ;
  assign n454 = n442 ^ x13 ;
  assign n455 = n442 ^ n149 ;
  assign n456 = n455 ^ n149 ;
  assign n457 = n26 & n269 ;
  assign n458 = ~n334 & ~n457 ;
  assign n459 = n458 ^ n149 ;
  assign n460 = ~n456 & ~n459 ;
  assign n461 = n460 ^ n149 ;
  assign n462 = n454 & ~n461 ;
  assign n463 = n462 ^ x13 ;
  assign n464 = ~n151 & ~n463 ;
  assign n465 = n49 & ~n464 ;
  assign n466 = x10 ^ x8 ;
  assign n467 = n466 ^ x8 ;
  assign n468 = x11 ^ x8 ;
  assign n469 = n468 ^ x8 ;
  assign n470 = n467 & n469 ;
  assign n471 = n470 ^ x8 ;
  assign n472 = x13 & ~n471 ;
  assign n473 = n472 ^ x8 ;
  assign n474 = n113 & n473 ;
  assign n475 = x13 & ~n65 ;
  assign n476 = ~n110 & ~n156 ;
  assign n477 = n475 & n476 ;
  assign n478 = n149 & ~n477 ;
  assign n479 = n19 & ~n478 ;
  assign n480 = ~n474 & n479 ;
  assign n481 = ~n465 & ~n480 ;
  assign n482 = ~x9 & n481 ;
  assign n483 = ~n453 & ~n482 ;
  assign n484 = n73 & n83 ;
  assign n485 = x9 & n484 ;
  assign n486 = n160 & n485 ;
  assign n487 = ~x4 & n486 ;
  assign n488 = ~n483 & ~n487 ;
  assign n489 = ~n440 & n488 ;
  assign n490 = x5 & ~n489 ;
  assign n491 = n490 ^ n147 ;
  assign n492 = n491 ^ n147 ;
  assign n493 = n492 ^ n323 ;
  assign n494 = n323 & ~n493 ;
  assign n495 = n494 ^ n323 ;
  assign n496 = ~n324 & n495 ;
  assign n497 = n496 ^ n494 ;
  assign n498 = n497 ^ n147 ;
  assign n499 = n498 ^ n323 ;
  assign n500 = x0 & n499 ;
  assign n501 = n500 ^ n147 ;
  assign n502 = x5 & n49 ;
  assign n503 = ~x14 & n502 ;
  assign n504 = x4 & n414 ;
  assign n505 = ~x7 & ~n504 ;
  assign n506 = n503 & ~n505 ;
  assign n507 = ~n130 & n506 ;
  assign n508 = n108 & ~n111 ;
  assign n509 = ~x3 & n368 ;
  assign n510 = ~n508 & ~n509 ;
  assign n511 = n510 ^ x5 ;
  assign n512 = n511 ^ n510 ;
  assign n513 = n512 ^ n507 ;
  assign n514 = ~x4 & ~n155 ;
  assign n515 = x7 & n19 ;
  assign n516 = ~n514 & ~n515 ;
  assign n517 = n516 ^ x13 ;
  assign n518 = x13 & ~n517 ;
  assign n519 = n518 ^ n510 ;
  assign n520 = n519 ^ x13 ;
  assign n521 = n513 & ~n520 ;
  assign n522 = n521 ^ n518 ;
  assign n523 = n522 ^ x13 ;
  assign n524 = ~n507 & n523 ;
  assign n525 = n524 ^ n507 ;
  assign n526 = ~x2 & n525 ;
  assign n527 = ~x4 & ~x14 ;
  assign n528 = ~n338 & ~n527 ;
  assign n529 = ~x14 & x16 ;
  assign n530 = n528 & ~n529 ;
  assign n531 = x15 & n60 ;
  assign n532 = n21 & n531 ;
  assign n533 = ~n530 & n532 ;
  assign n534 = ~n526 & ~n533 ;
  assign n535 = n534 ^ x6 ;
  assign n536 = n535 ^ n534 ;
  assign n537 = n536 ^ n501 ;
  assign n538 = ~x2 & ~x5 ;
  assign n539 = n19 & n538 ;
  assign n540 = n49 & n50 ;
  assign n541 = n302 & n540 ;
  assign n542 = ~n539 & ~n541 ;
  assign n543 = ~x5 & x15 ;
  assign n544 = ~x8 & n543 ;
  assign n545 = ~n528 & n544 ;
  assign n546 = n542 & ~n545 ;
  assign n547 = n546 ^ x13 ;
  assign n548 = x13 & ~n547 ;
  assign n549 = n548 ^ n534 ;
  assign n550 = n549 ^ x13 ;
  assign n551 = n537 & ~n550 ;
  assign n552 = n551 ^ n548 ;
  assign n553 = n552 ^ x13 ;
  assign n554 = n501 & n553 ;
  assign n555 = n554 ^ n501 ;
  assign n556 = ~x1 & ~n555 ;
  assign n557 = x0 & n58 ;
  assign n558 = ~x9 & n180 ;
  assign n559 = n368 & ~n558 ;
  assign n560 = ~n108 & ~n559 ;
  assign n561 = x4 & ~n560 ;
  assign n562 = ~x4 & n18 ;
  assign n563 = n422 ^ x9 ;
  assign n564 = n563 ^ n422 ;
  assign n565 = ~n232 & ~n360 ;
  assign n566 = n565 ^ n422 ;
  assign n567 = n564 & ~n566 ;
  assign n568 = n567 ^ n422 ;
  assign n569 = n562 & n568 ;
  assign n570 = ~n561 & ~n569 ;
  assign n571 = n75 & ~n570 ;
  assign n572 = n106 & n381 ;
  assign n573 = ~x6 & n502 ;
  assign n574 = n338 & n573 ;
  assign n575 = n268 & n336 ;
  assign n576 = n76 & n368 ;
  assign n577 = x6 & n18 ;
  assign n578 = x6 & x7 ;
  assign n579 = n49 & ~n578 ;
  assign n580 = ~n577 & ~n579 ;
  assign n581 = n22 & n83 ;
  assign n582 = ~n580 & n581 ;
  assign n583 = ~n576 & ~n582 ;
  assign n584 = ~n575 & n583 ;
  assign n585 = ~n574 & n584 ;
  assign n586 = x1 & ~n585 ;
  assign n587 = ~n572 & ~n586 ;
  assign n588 = n587 ^ x1 ;
  assign n589 = n588 ^ n587 ;
  assign n590 = ~x13 & ~n386 ;
  assign n591 = n19 & ~n590 ;
  assign n592 = n72 & n591 ;
  assign n593 = x14 & ~n149 ;
  assign n594 = ~x7 & n150 ;
  assign n595 = ~n593 & ~n594 ;
  assign n596 = n22 & n577 ;
  assign n597 = ~n595 & n596 ;
  assign n598 = ~x6 & n367 ;
  assign n599 = x10 & ~x13 ;
  assign n600 = x4 & n599 ;
  assign n601 = n600 ^ x13 ;
  assign n602 = n598 & n601 ;
  assign n603 = x6 & x13 ;
  assign n604 = ~n338 & ~n355 ;
  assign n605 = ~n281 & n604 ;
  assign n606 = n269 & n271 ;
  assign n607 = ~n605 & ~n606 ;
  assign n608 = n603 & ~n607 ;
  assign n609 = ~n602 & ~n608 ;
  assign n610 = x5 & ~n609 ;
  assign n611 = ~n597 & ~n610 ;
  assign n612 = ~n592 & n611 ;
  assign n613 = n612 ^ n587 ;
  assign n614 = n613 ^ n587 ;
  assign n615 = n589 & ~n614 ;
  assign n616 = n615 ^ n587 ;
  assign n617 = ~x9 & ~n616 ;
  assign n618 = n617 ^ n587 ;
  assign n619 = ~n571 & n618 ;
  assign n620 = n557 & ~n619 ;
  assign n621 = ~x0 & x14 ;
  assign n622 = ~n67 & n502 ;
  assign n623 = n621 & n622 ;
  assign n624 = ~x0 & n578 ;
  assign n625 = ~n27 & ~n624 ;
  assign n626 = n503 & ~n625 ;
  assign n627 = ~n168 & ~n626 ;
  assign n628 = ~x0 & x4 ;
  assign n629 = ~n73 & n628 ;
  assign n630 = n629 ^ n18 ;
  assign n631 = ~n72 & ~n75 ;
  assign n632 = n631 ^ n19 ;
  assign n633 = ~n630 & n632 ;
  assign n634 = n633 ^ n631 ;
  assign n635 = n19 & n634 ;
  assign n636 = n627 & ~n635 ;
  assign n637 = ~n623 & n636 ;
  assign n638 = x13 & ~n637 ;
  assign n639 = n527 & ~n578 ;
  assign n640 = n502 & n639 ;
  assign n641 = n18 & n621 ;
  assign n642 = ~n77 & n641 ;
  assign n643 = ~n640 & ~n642 ;
  assign n644 = n58 & n643 ;
  assign n645 = ~n638 & n644 ;
  assign n646 = x2 & ~n641 ;
  assign n647 = ~n49 & n646 ;
  assign n648 = ~x4 & ~x5 ;
  assign n649 = ~x6 & n648 ;
  assign n650 = x2 & n649 ;
  assign n651 = ~n125 & n302 ;
  assign n652 = ~n108 & n651 ;
  assign n653 = ~n650 & ~n652 ;
  assign n654 = x1 & n653 ;
  assign n655 = ~n647 & n654 ;
  assign n656 = ~n645 & n655 ;
  assign n657 = ~x2 & n50 ;
  assign n658 = x3 & n657 ;
  assign n659 = x6 & ~x7 ;
  assign n660 = n367 & n659 ;
  assign n661 = n125 & n578 ;
  assign n662 = n621 & n661 ;
  assign n663 = n662 ^ n658 ;
  assign n664 = n660 & n663 ;
  assign n665 = n664 ^ n662 ;
  assign n666 = n658 & n665 ;
  assign n667 = n650 ^ n49 ;
  assign n668 = n667 ^ n666 ;
  assign n669 = n603 & n658 ;
  assign n670 = n355 & n669 ;
  assign n671 = n670 ^ n641 ;
  assign n672 = ~n650 & ~n671 ;
  assign n673 = n672 ^ n641 ;
  assign n674 = ~n668 & ~n673 ;
  assign n675 = n674 ^ n672 ;
  assign n676 = n675 ^ n641 ;
  assign n677 = n676 ^ n650 ;
  assign n678 = ~n666 & n677 ;
  assign n679 = ~n656 & n678 ;
  assign n680 = ~x1 & ~n649 ;
  assign n681 = n226 & ~n680 ;
  assign n682 = ~n345 & ~n346 ;
  assign n683 = ~n681 & n682 ;
  assign n684 = n87 ^ x14 ;
  assign n685 = n27 & n128 ;
  assign n686 = ~x2 & ~n685 ;
  assign n687 = n686 ^ n87 ;
  assign n688 = n687 ^ n686 ;
  assign n689 = n688 ^ n684 ;
  assign n690 = x4 ^ x1 ;
  assign n691 = x6 & n690 ;
  assign n692 = n691 ^ x1 ;
  assign n693 = n692 ^ n327 ;
  assign n694 = ~n692 & n693 ;
  assign n695 = n694 ^ n686 ;
  assign n696 = n695 ^ n692 ;
  assign n697 = n689 & n696 ;
  assign n698 = n697 ^ n694 ;
  assign n699 = n698 ^ n692 ;
  assign n700 = n684 & ~n699 ;
  assign n701 = n700 ^ x14 ;
  assign n702 = n349 & ~n701 ;
  assign n703 = ~n91 & n442 ;
  assign n704 = ~n91 & n648 ;
  assign n705 = n95 & n125 ;
  assign n706 = ~n704 & n705 ;
  assign n707 = ~n703 & n706 ;
  assign n708 = ~x1 & n707 ;
  assign n709 = n680 & ~n703 ;
  assign n710 = n250 & ~n709 ;
  assign n711 = ~n682 & ~n710 ;
  assign n712 = ~n708 & n711 ;
  assign n713 = ~n702 & n712 ;
  assign n714 = ~n683 & ~n713 ;
  assign n715 = x0 & n714 ;
  assign n716 = n679 & ~n715 ;
  assign n717 = ~n620 & n716 ;
  assign n718 = ~n556 & n717 ;
  assign n719 = n718 ^ x13 ;
  assign n720 = n719 ^ x12 ;
  assign n871 = n720 ^ n719 ;
  assign n721 = x12 & n19 ;
  assign n722 = n91 & n721 ;
  assign n723 = ~x2 & n722 ;
  assign n724 = x0 & x9 ;
  assign n725 = ~x7 & ~n724 ;
  assign n726 = ~n110 & ~n302 ;
  assign n727 = n19 & n726 ;
  assign n728 = n727 ^ x4 ;
  assign n729 = n728 ^ n727 ;
  assign n730 = ~x2 & n49 ;
  assign n731 = n730 ^ n727 ;
  assign n732 = n731 ^ n727 ;
  assign n733 = n729 & n732 ;
  assign n734 = n733 ^ n727 ;
  assign n735 = ~x5 & n734 ;
  assign n736 = n735 ^ n727 ;
  assign n737 = n725 & n736 ;
  assign n738 = n514 & n538 ;
  assign n739 = x0 & ~x5 ;
  assign n740 = n316 & n739 ;
  assign n741 = n49 & n740 ;
  assign n742 = ~n738 & ~n741 ;
  assign n743 = ~x11 & n94 ;
  assign n744 = n307 & ~n743 ;
  assign n745 = n105 & ~n301 ;
  assign n746 = ~n744 & ~n745 ;
  assign n747 = n746 ^ n59 ;
  assign n748 = n747 ^ x0 ;
  assign n755 = n748 ^ n747 ;
  assign n749 = n748 ^ n94 ;
  assign n750 = n749 ^ n747 ;
  assign n751 = n94 ^ n59 ;
  assign n752 = n751 ^ n94 ;
  assign n753 = n752 ^ n750 ;
  assign n754 = ~n750 & ~n753 ;
  assign n756 = n755 ^ n754 ;
  assign n757 = n756 ^ n750 ;
  assign n758 = n747 ^ x8 ;
  assign n759 = n754 ^ n750 ;
  assign n760 = n758 & ~n759 ;
  assign n761 = n760 ^ n747 ;
  assign n762 = ~n757 & ~n761 ;
  assign n763 = n762 ^ n747 ;
  assign n764 = n763 ^ n59 ;
  assign n765 = n764 ^ n747 ;
  assign n766 = n502 & n765 ;
  assign n767 = x5 & ~x8 ;
  assign n773 = n58 & n280 ;
  assign n774 = x14 & n773 ;
  assign n769 = x0 & x10 ;
  assign n770 = ~n724 & ~n769 ;
  assign n771 = x5 & n770 ;
  assign n775 = n774 ^ n771 ;
  assign n786 = n775 ^ n771 ;
  assign n787 = n786 ^ n771 ;
  assign n788 = n786 & n787 ;
  assign n777 = x11 & n769 ;
  assign n778 = ~x8 & ~n777 ;
  assign n779 = n336 & ~n778 ;
  assign n768 = ~n302 & ~n724 ;
  assign n772 = n771 ^ n768 ;
  assign n776 = n775 ^ n772 ;
  assign n780 = n779 ^ n776 ;
  assign n781 = n780 ^ n776 ;
  assign n782 = n776 ^ n775 ;
  assign n783 = n782 ^ n771 ;
  assign n784 = n781 & n783 ;
  assign n791 = n788 ^ n784 ;
  assign n785 = n784 ^ n767 ;
  assign n789 = n788 ^ n786 ;
  assign n790 = n785 & n789 ;
  assign n792 = n791 ^ n790 ;
  assign n793 = n767 & n792 ;
  assign n794 = n793 ^ n784 ;
  assign n795 = n794 ^ n788 ;
  assign n796 = n795 ^ n790 ;
  assign n797 = n796 ^ n774 ;
  assign n798 = ~n766 & ~n797 ;
  assign n799 = n798 ^ x7 ;
  assign n800 = n799 ^ n798 ;
  assign n801 = n800 ^ n742 ;
  assign n802 = n72 & ~n724 ;
  assign n803 = ~n64 & ~n802 ;
  assign n804 = n803 ^ n49 ;
  assign n805 = ~n803 & ~n804 ;
  assign n806 = n805 ^ n798 ;
  assign n807 = n806 ^ n803 ;
  assign n808 = n801 & n807 ;
  assign n809 = n808 ^ n805 ;
  assign n810 = n809 ^ n803 ;
  assign n811 = n742 & ~n810 ;
  assign n812 = n811 ^ n742 ;
  assign n813 = ~n737 & n812 ;
  assign n814 = x12 & ~n813 ;
  assign n815 = x0 & n50 ;
  assign n816 = n308 & n815 ;
  assign n817 = n49 & n816 ;
  assign n818 = ~n593 & ~n621 ;
  assign n819 = n72 & n768 ;
  assign n820 = n18 & n819 ;
  assign n821 = ~n818 & n820 ;
  assign n822 = n338 & ~n770 ;
  assign n823 = ~n527 & ~n822 ;
  assign n824 = n58 & n502 ;
  assign n825 = ~n823 & n824 ;
  assign n826 = ~n821 & ~n825 ;
  assign n827 = ~n817 & n826 ;
  assign n828 = n26 & ~n827 ;
  assign n829 = x2 & n725 ;
  assign n830 = ~n721 & ~n829 ;
  assign n831 = ~n302 & n725 ;
  assign n832 = ~n148 & n831 ;
  assign n833 = ~x12 & ~n778 ;
  assign n834 = ~n832 & ~n833 ;
  assign n835 = ~n648 & n834 ;
  assign n836 = ~n830 & n835 ;
  assign n837 = ~n828 & ~n836 ;
  assign n838 = ~n814 & n837 ;
  assign n839 = ~x6 & ~n838 ;
  assign n840 = x3 & ~n659 ;
  assign n841 = n338 & n770 ;
  assign n842 = x7 & ~n841 ;
  assign n843 = n840 & ~n842 ;
  assign n844 = n730 & ~n843 ;
  assign n845 = n336 & ~n557 ;
  assign n846 = ~x11 & n724 ;
  assign n847 = x8 & n846 ;
  assign n848 = ~n316 & n847 ;
  assign n849 = n148 & ~n848 ;
  assign n850 = ~n845 & ~n849 ;
  assign n851 = x6 & ~n850 ;
  assign n852 = ~n844 & ~n851 ;
  assign n853 = x12 & ~n852 ;
  assign n854 = x6 & n95 ;
  assign n855 = n846 & n854 ;
  assign n856 = n280 & n855 ;
  assign n857 = ~n853 & ~n856 ;
  assign n858 = x5 & ~n857 ;
  assign n859 = ~n839 & ~n858 ;
  assign n860 = ~n723 & n859 ;
  assign n861 = ~x1 & ~n860 ;
  assign n862 = n658 & n770 ;
  assign n863 = n598 & n862 ;
  assign n864 = ~n861 & ~n863 ;
  assign n865 = n864 ^ n720 ;
  assign n866 = n865 ^ n719 ;
  assign n867 = n720 ^ n718 ;
  assign n868 = n867 ^ n864 ;
  assign n869 = n868 ^ n866 ;
  assign n870 = ~n866 & n869 ;
  assign n872 = n871 ^ n870 ;
  assign n873 = n872 ^ n866 ;
  assign n874 = ~n155 & n650 ;
  assign n875 = n502 ^ x4 ;
  assign n876 = n875 ^ x2 ;
  assign n883 = n876 ^ n875 ;
  assign n878 = n19 & n25 ;
  assign n877 = n876 ^ n502 ;
  assign n879 = n878 ^ n877 ;
  assign n880 = n878 ^ n876 ;
  assign n881 = n880 ^ n875 ;
  assign n882 = ~n879 & ~n881 ;
  assign n884 = n883 ^ n882 ;
  assign n885 = n49 & ~n91 ;
  assign n886 = n885 ^ n876 ;
  assign n887 = n883 & ~n886 ;
  assign n888 = n887 ^ n885 ;
  assign n889 = n884 & n888 ;
  assign n890 = n889 ^ n882 ;
  assign n891 = n890 ^ n876 ;
  assign n892 = n891 ^ x4 ;
  assign n893 = n892 ^ n875 ;
  assign n894 = ~n539 & n893 ;
  assign n895 = x14 & n840 ;
  assign n896 = n771 & n895 ;
  assign n897 = n49 & n72 ;
  assign n898 = ~n730 & ~n897 ;
  assign n899 = ~n896 & ~n898 ;
  assign n900 = ~n845 & ~n899 ;
  assign n901 = n900 ^ x6 ;
  assign n902 = n900 ^ x5 ;
  assign n903 = n902 ^ x5 ;
  assign n904 = n336 ^ x5 ;
  assign n905 = n903 & ~n904 ;
  assign n906 = n905 ^ x5 ;
  assign n907 = n901 & n906 ;
  assign n908 = n907 ^ x6 ;
  assign n909 = n894 & n908 ;
  assign n910 = x1 & ~n909 ;
  assign n911 = ~n530 & n543 ;
  assign n912 = ~n225 & ~n280 ;
  assign n913 = n139 & ~n912 ;
  assign n914 = n170 & n770 ;
  assign n915 = x0 & n18 ;
  assign n916 = ~n914 & ~n915 ;
  assign n917 = x14 & n658 ;
  assign n918 = ~n916 & n917 ;
  assign n919 = ~n913 & ~n918 ;
  assign n920 = ~n911 & n919 ;
  assign n921 = x6 & ~n920 ;
  assign n922 = ~n910 & ~n921 ;
  assign n923 = ~n874 & n922 ;
  assign n924 = n923 ^ n719 ;
  assign n925 = n870 ^ n866 ;
  assign n926 = n924 & ~n925 ;
  assign n927 = n926 ^ n719 ;
  assign n928 = n873 & n927 ;
  assign n929 = n928 ^ n719 ;
  assign n930 = n929 ^ x13 ;
  assign n931 = n930 ^ n719 ;
  assign y0 = ~n931 ;
endmodule
