// Benchmark "./inc.pla" written by ABC on Thu Apr 23 10:59:53 2020

module \./inc.pla  ( 
    x0, x1, x2, x3, x4, x5, x6,
    z6  );
  input  x0, x1, x2, x3, x4, x5, x6;
  output z6;
  assign z6 = 1'b1;
endmodule


