module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 ;
  assign n15 = ~x6 & ~x7 ;
  assign n16 = x5 & x12 ;
  assign n17 = ~n15 & n16 ;
  assign n18 = ~x8 & x11 ;
  assign n19 = ~x9 & n18 ;
  assign n21 = n19 ^ x5 ;
  assign n30 = n21 ^ n19 ;
  assign n20 = n19 ^ x10 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n23 ^ n19 ;
  assign n25 = n22 ^ x7 ;
  assign n26 = n25 ^ x6 ;
  assign n27 = n26 ^ n22 ;
  assign n28 = n27 ^ n24 ;
  assign n29 = n24 & ~n28 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = n19 ^ x6 ;
  assign n34 = n29 ^ n24 ;
  assign n35 = n33 & n34 ;
  assign n36 = n35 ^ n19 ;
  assign n37 = ~n32 & ~n36 ;
  assign n38 = n37 ^ n19 ;
  assign n39 = n38 ^ x5 ;
  assign n40 = n39 ^ n19 ;
  assign n41 = ~n17 & n40 ;
  assign n42 = x2 & x13 ;
  assign n43 = x0 & x1 ;
  assign n44 = x4 & n43 ;
  assign n45 = x3 & n44 ;
  assign n46 = n42 & n45 ;
  assign n47 = ~n41 & n46 ;
  assign y0 = n47 ;
endmodule
