module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 ;
  assign n8 = ~x1 & x3 ;
  assign n18 = x1 & ~x3 ;
  assign n19 = x4 & x5 ;
  assign n20 = ~n18 & n19 ;
  assign n9 = x5 & x6 ;
  assign n10 = n9 ^ x1 ;
  assign n11 = n10 ^ x1 ;
  assign n12 = x4 ^ x1 ;
  assign n13 = n12 ^ x1 ;
  assign n14 = ~n11 & ~n13 ;
  assign n15 = n14 ^ x1 ;
  assign n16 = x3 & n15 ;
  assign n17 = n16 ^ x1 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = n21 ^ x0 ;
  assign n29 = n22 ^ n21 ;
  assign n23 = n22 ^ x1 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n22 ^ n17 ;
  assign n26 = n25 ^ x1 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = ~n24 & ~n27 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = n30 ^ n24 ;
  assign n32 = n21 ^ x6 ;
  assign n33 = n28 ^ n24 ;
  assign n34 = ~n32 & ~n33 ;
  assign n35 = n34 ^ n21 ;
  assign n36 = n31 & n35 ;
  assign n37 = n36 ^ n21 ;
  assign n38 = n37 ^ n20 ;
  assign n39 = n38 ^ n21 ;
  assign n40 = ~n8 & ~n39 ;
  assign n41 = ~x2 & ~n40 ;
  assign n42 = x1 ^ x0 ;
  assign n43 = n42 ^ x1 ;
  assign n44 = n43 ^ x2 ;
  assign n45 = n8 ^ x4 ;
  assign n46 = x4 & n45 ;
  assign n47 = n46 ^ x1 ;
  assign n48 = n47 ^ x4 ;
  assign n49 = n44 & n48 ;
  assign n50 = n49 ^ n46 ;
  assign n51 = n50 ^ x4 ;
  assign n52 = x2 & n51 ;
  assign n53 = n52 ^ x2 ;
  assign n54 = ~n41 & ~n53 ;
  assign y0 = ~n54 ;
endmodule
