module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 ;
  assign n9 = x7 ^ x6 ;
  assign n10 = ~x2 & n9 ;
  assign n11 = n10 ^ x6 ;
  assign n13 = n11 ^ x4 ;
  assign n12 = n11 ^ x5 ;
  assign n14 = n13 ^ n12 ;
  assign n15 = n13 ^ x2 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = n14 & ~n16 ;
  assign n18 = n17 ^ n13 ;
  assign n19 = x1 & n18 ;
  assign n20 = n19 ^ n11 ;
  assign n21 = n20 ^ x3 ;
  assign n22 = ~x0 & n21 ;
  assign n23 = n22 ^ x3 ;
  assign y0 = n23 ;
endmodule
