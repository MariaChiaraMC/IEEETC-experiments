module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 ;
  assign n9 = ~x3 & ~x5 ;
  assign n10 = x6 & n9 ;
  assign n11 = x6 & x7 ;
  assign n12 = ~x5 & ~n11 ;
  assign n13 = x3 & ~n12 ;
  assign n14 = ~x2 & n13 ;
  assign n15 = ~n10 & ~n14 ;
  assign n16 = ~x4 & ~n15 ;
  assign n20 = x3 ^ x2 ;
  assign n17 = x6 ^ x3 ;
  assign n18 = n17 ^ x5 ;
  assign n19 = n18 ^ n17 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = n20 ^ x6 ;
  assign n23 = n22 ^ n17 ;
  assign n24 = n23 ^ n18 ;
  assign n25 = n24 ^ n17 ;
  assign n29 = n25 ^ n17 ;
  assign n30 = n29 ^ n21 ;
  assign n26 = n20 ^ x7 ;
  assign n27 = n26 ^ n20 ;
  assign n28 = n27 ^ n25 ;
  assign n31 = n30 ^ n28 ;
  assign n32 = n21 & n31 ;
  assign n33 = n32 ^ n25 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = n34 ^ n20 ;
  assign n36 = n20 ^ x4 ;
  assign n37 = n36 ^ n18 ;
  assign n38 = n37 ^ n20 ;
  assign n39 = n38 ^ n25 ;
  assign n40 = n39 ^ n27 ;
  assign n41 = n40 ^ n21 ;
  assign n42 = n41 ^ n30 ;
  assign n43 = n30 & n42 ;
  assign n44 = n43 ^ n25 ;
  assign n45 = n44 ^ n38 ;
  assign n46 = n45 ^ n20 ;
  assign n47 = n27 ^ n21 ;
  assign n48 = n47 ^ n30 ;
  assign n49 = n25 ^ n21 ;
  assign n50 = n49 ^ n20 ;
  assign n51 = n48 & n50 ;
  assign n52 = n51 ^ n25 ;
  assign n53 = n52 ^ n27 ;
  assign n54 = n53 ^ n21 ;
  assign n55 = n46 & n54 ;
  assign n56 = n55 ^ n25 ;
  assign n57 = n56 ^ n30 ;
  assign n58 = n35 & n57 ;
  assign n59 = n58 ^ x3 ;
  assign n60 = ~n16 & n59 ;
  assign n61 = ~x0 & ~n60 ;
  assign n62 = ~x1 & n61 ;
  assign y0 = n62 ;
endmodule
