module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n7 = x2 ^ x1 ;
  assign n8 = x5 & n7 ;
  assign n9 = x4 ^ x3 ;
  assign n10 = n9 ^ x0 ;
  assign n12 = n10 ^ x4 ;
  assign n13 = n12 ^ n10 ;
  assign n11 = n10 ^ x2 ;
  assign n14 = n13 ^ n11 ;
  assign n15 = n10 ^ x0 ;
  assign n16 = n15 ^ n10 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = ~n13 & n17 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = n14 & ~n19 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = n21 ^ n10 ;
  assign n23 = n22 ^ n13 ;
  assign n24 = n8 & ~n23 ;
  assign y0 = ~n24 ;
endmodule
