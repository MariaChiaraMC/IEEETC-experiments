module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ;
  assign n8 = ~x5 & ~x6 ;
  assign n9 = x1 & ~x4 ;
  assign n10 = ~n8 & ~n9 ;
  assign n11 = n10 ^ x0 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = ~x4 & ~x5 ;
  assign n14 = n13 ^ n10 ;
  assign n15 = n12 & n14 ;
  assign n16 = n15 ^ n10 ;
  assign n17 = ~x3 & n16 ;
  assign n18 = x5 & x6 ;
  assign n19 = x2 ^ x1 ;
  assign n20 = n19 ^ x2 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = x2 ^ x0 ;
  assign n23 = n22 ^ x4 ;
  assign n24 = ~x4 & n23 ;
  assign n25 = n24 ^ x2 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = n21 & n26 ;
  assign n28 = n27 ^ n24 ;
  assign n29 = n28 ^ x4 ;
  assign n30 = ~n18 & ~n29 ;
  assign n31 = n17 & n30 ;
  assign n32 = ~x1 & x2 ;
  assign n33 = ~x0 & n32 ;
  assign n34 = n18 ^ n8 ;
  assign n35 = ~x4 & n34 ;
  assign n36 = n35 ^ n8 ;
  assign n37 = n33 & n36 ;
  assign n38 = x3 & n37 ;
  assign n39 = ~n31 & ~n38 ;
  assign y0 = ~n39 ;
endmodule
