module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 ;
  assign n9 = x3 ^ x2 ;
  assign n10 = n9 ^ x2 ;
  assign n13 = x4 ^ x2 ;
  assign n14 = n13 ^ x6 ;
  assign n11 = x5 ^ x4 ;
  assign n12 = n11 ^ x6 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n15 ^ x4 ;
  assign n17 = x6 ^ x4 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = n18 ^ n14 ;
  assign n20 = n19 ^ x4 ;
  assign n21 = n20 ^ x7 ;
  assign n22 = n21 ^ n12 ;
  assign n23 = ~n14 & ~n22 ;
  assign n24 = n23 ^ x4 ;
  assign n25 = n24 ^ n16 ;
  assign n26 = n20 ^ n14 ;
  assign n27 = n26 ^ n16 ;
  assign n28 = x4 & n27 ;
  assign n29 = n28 ^ n14 ;
  assign n30 = ~n25 & ~n29 ;
  assign n31 = ~n16 & n30 ;
  assign n32 = n31 ^ n23 ;
  assign n33 = n32 ^ n28 ;
  assign n34 = n33 ^ n30 ;
  assign n35 = x3 ^ x1 ;
  assign n36 = n35 ^ n10 ;
  assign n37 = n36 ^ n10 ;
  assign n38 = ~n34 & ~n37 ;
  assign n39 = n38 ^ x2 ;
  assign n40 = x4 & ~x5 ;
  assign n41 = n40 ^ x2 ;
  assign n42 = ~n36 & ~n41 ;
  assign n43 = n42 ^ n10 ;
  assign n44 = n43 ^ n36 ;
  assign n45 = n39 & ~n44 ;
  assign n46 = n10 & n45 ;
  assign n47 = n46 ^ n38 ;
  assign n48 = n47 ^ x1 ;
  assign y0 = n48 ;
endmodule
