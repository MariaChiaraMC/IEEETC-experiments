// Benchmark "./newcwp.pla" written by ABC on Thu Apr 23 10:59:58 2020

module \./newcwp.pla  ( 
    x0, x1, x2, x3,
    z3  );
  input  x0, x1, x2, x3;
  output z3;
  assign z3 = 1'b1;
endmodule


