module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 ;
  assign n18 = ~x0 & ~x8 ;
  assign n19 = n18 ^ x0 ;
  assign n20 = ~x1 & n19 ;
  assign n21 = n20 ^ x0 ;
  assign n22 = n21 ^ x13 ;
  assign n23 = n22 ^ x13 ;
  assign n16 = x13 ^ x12 ;
  assign n17 = n16 ^ x13 ;
  assign n24 = n23 ^ n17 ;
  assign n25 = x9 & ~x13 ;
  assign n26 = n25 ^ x13 ;
  assign n27 = n26 ^ x13 ;
  assign n28 = n27 ^ n23 ;
  assign n29 = ~n23 & ~n28 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = ~n24 & ~n30 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = n32 ^ x13 ;
  assign n34 = n33 ^ n23 ;
  assign n35 = x11 & ~n34 ;
  assign n36 = n35 ^ x13 ;
  assign n37 = x10 & n36 ;
  assign n38 = x14 ^ x0 ;
  assign n39 = x14 ^ x8 ;
  assign n40 = n39 ^ x8 ;
  assign n41 = ~x2 & ~x3 ;
  assign n42 = n41 ^ x8 ;
  assign n43 = n40 & n42 ;
  assign n44 = n43 ^ x8 ;
  assign n45 = ~n38 & ~n44 ;
  assign n46 = ~x1 & n45 ;
  assign n47 = x0 & x1 ;
  assign n48 = x9 & ~n47 ;
  assign n49 = ~x11 & n48 ;
  assign n50 = ~x14 & ~n49 ;
  assign n51 = x10 & ~n50 ;
  assign n52 = ~n46 & n51 ;
  assign n53 = ~x13 & ~x14 ;
  assign n54 = n53 ^ x9 ;
  assign n55 = n54 ^ x11 ;
  assign n67 = n55 ^ n54 ;
  assign n57 = n41 ^ x4 ;
  assign n58 = n57 ^ x4 ;
  assign n59 = n21 ^ x4 ;
  assign n60 = ~n58 & n59 ;
  assign n61 = n60 ^ x4 ;
  assign n62 = x13 & ~n61 ;
  assign n56 = n55 ^ n53 ;
  assign n63 = n62 ^ n56 ;
  assign n64 = n62 ^ n55 ;
  assign n65 = n64 ^ n54 ;
  assign n66 = ~n63 & ~n65 ;
  assign n68 = n67 ^ n66 ;
  assign n69 = ~x13 & n47 ;
  assign n70 = x5 & x6 ;
  assign n71 = ~x2 & ~x4 ;
  assign n72 = ~n70 & n71 ;
  assign n73 = n72 ^ x3 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = n74 ^ n69 ;
  assign n76 = ~x5 & ~x7 ;
  assign n77 = ~x4 & ~x6 ;
  assign n78 = n76 & ~n77 ;
  assign n79 = x4 & x5 ;
  assign n80 = x2 & ~n79 ;
  assign n81 = n80 ^ n78 ;
  assign n82 = ~n78 & n81 ;
  assign n83 = n82 ^ n72 ;
  assign n84 = n83 ^ n78 ;
  assign n85 = ~n75 & n84 ;
  assign n86 = n85 ^ n82 ;
  assign n87 = n86 ^ n78 ;
  assign n88 = n69 & ~n87 ;
  assign n89 = n88 ^ n69 ;
  assign n90 = ~x0 & x1 ;
  assign n91 = x13 & ~n90 ;
  assign n92 = x1 ^ x0 ;
  assign n93 = x6 ^ x1 ;
  assign n94 = n93 ^ n92 ;
  assign n95 = n79 ^ x5 ;
  assign n96 = ~x1 & n95 ;
  assign n97 = n96 ^ n79 ;
  assign n98 = n94 & n97 ;
  assign n99 = n98 ^ n96 ;
  assign n100 = n99 ^ n79 ;
  assign n101 = n100 ^ x1 ;
  assign n102 = ~n92 & ~n101 ;
  assign n103 = n102 ^ x0 ;
  assign n104 = ~n91 & ~n103 ;
  assign n105 = n104 ^ x1 ;
  assign n106 = n105 ^ n89 ;
  assign n121 = ~x4 & n76 ;
  assign n122 = ~x3 & ~n121 ;
  assign n123 = x2 & ~n122 ;
  assign n107 = x3 ^ x2 ;
  assign n108 = n107 ^ x0 ;
  assign n109 = x4 & x6 ;
  assign n110 = n109 ^ x2 ;
  assign n111 = n76 ^ x5 ;
  assign n112 = x2 ^ x0 ;
  assign n113 = ~n111 & n112 ;
  assign n114 = n113 ^ n76 ;
  assign n115 = n114 ^ n111 ;
  assign n116 = n110 & ~n115 ;
  assign n117 = n116 ^ x2 ;
  assign n118 = n108 & n117 ;
  assign n119 = n118 ^ n116 ;
  assign n120 = x0 & n119 ;
  assign n124 = n123 ^ n120 ;
  assign n125 = ~n104 & ~n124 ;
  assign n126 = n125 ^ n123 ;
  assign n127 = n106 & ~n126 ;
  assign n128 = n127 ^ n125 ;
  assign n129 = n128 ^ n123 ;
  assign n130 = n129 ^ n104 ;
  assign n131 = ~n89 & n130 ;
  assign n132 = ~x10 & ~n131 ;
  assign n133 = n132 ^ n55 ;
  assign n134 = n67 & n133 ;
  assign n135 = n134 ^ n132 ;
  assign n136 = n68 & n135 ;
  assign n137 = n136 ^ n66 ;
  assign n138 = n137 ^ n55 ;
  assign n139 = n138 ^ x9 ;
  assign n140 = n139 ^ n54 ;
  assign n141 = ~n52 & n140 ;
  assign n142 = ~x12 & ~n141 ;
  assign n143 = ~n37 & ~n142 ;
  assign y0 = ~n143 ;
endmodule
