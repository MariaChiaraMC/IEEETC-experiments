module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 ;
  assign n9 = ~x6 & x7 ;
  assign n10 = ~x2 & ~x5 ;
  assign n11 = n9 & n10 ;
  assign n12 = ~x1 & n11 ;
  assign n13 = x3 & ~x5 ;
  assign n14 = x6 & ~x7 ;
  assign n15 = n13 & ~n14 ;
  assign n16 = x1 & n15 ;
  assign n19 = ~x3 & x5 ;
  assign n17 = n13 ^ x6 ;
  assign n18 = n17 ^ x1 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = n20 ^ n19 ;
  assign n31 = n21 ^ n20 ;
  assign n28 = n17 ^ n13 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = n32 ^ n28 ;
  assign n22 = x5 & ~x7 ;
  assign n24 = n22 ^ n13 ;
  assign n34 = n24 ^ n20 ;
  assign n35 = n34 ^ n28 ;
  assign n36 = ~n33 & ~n35 ;
  assign n23 = n22 ^ n20 ;
  assign n25 = n24 ^ n23 ;
  assign n26 = n25 ^ n20 ;
  assign n27 = n26 ^ n21 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n21 & ~n29 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = n37 ^ n21 ;
  assign n39 = n30 ^ n28 ;
  assign n40 = n39 ^ n32 ;
  assign n41 = ~n28 & ~n40 ;
  assign n42 = n41 ^ n30 ;
  assign n43 = n38 & n42 ;
  assign n44 = n43 ^ n36 ;
  assign n45 = n44 ^ n41 ;
  assign n46 = n45 ^ n21 ;
  assign n47 = n46 ^ n28 ;
  assign n48 = n47 ^ n32 ;
  assign n49 = n48 ^ n17 ;
  assign n50 = n49 ^ x2 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = x7 ^ x6 ;
  assign n53 = x5 ^ x3 ;
  assign n54 = x7 ^ x5 ;
  assign n55 = n54 ^ x5 ;
  assign n56 = n53 & n55 ;
  assign n57 = n56 ^ x5 ;
  assign n58 = n52 & ~n57 ;
  assign n59 = x1 & n58 ;
  assign n60 = ~x5 & ~x7 ;
  assign n61 = x5 & x7 ;
  assign n62 = ~n60 & ~n61 ;
  assign n63 = x1 & ~x7 ;
  assign n64 = ~n9 & ~n63 ;
  assign n65 = x3 & n64 ;
  assign n66 = n62 & n65 ;
  assign n67 = ~n59 & ~n66 ;
  assign n68 = n67 ^ n49 ;
  assign n69 = n51 & n68 ;
  assign n70 = n69 ^ n49 ;
  assign n71 = ~n16 & n70 ;
  assign n72 = n71 ^ x4 ;
  assign n73 = n72 ^ n71 ;
  assign n74 = x3 ^ x2 ;
  assign n84 = n74 ^ x5 ;
  assign n81 = n74 ^ x6 ;
  assign n79 = n74 ^ x3 ;
  assign n82 = n81 ^ n79 ;
  assign n85 = n84 ^ n82 ;
  assign n76 = n74 ^ x1 ;
  assign n77 = n76 ^ x6 ;
  assign n75 = n74 ^ x7 ;
  assign n78 = n77 ^ n75 ;
  assign n80 = n79 ^ n78 ;
  assign n83 = n82 ^ n80 ;
  assign n86 = n85 ^ n83 ;
  assign n87 = n86 ^ n82 ;
  assign n88 = n87 ^ n79 ;
  assign n89 = n88 ^ n77 ;
  assign n90 = n89 ^ n74 ;
  assign n96 = n90 ^ n82 ;
  assign n92 = n85 ^ n79 ;
  assign n93 = n92 ^ n77 ;
  assign n94 = n93 ^ n79 ;
  assign n91 = n90 ^ n74 ;
  assign n95 = n94 ^ n91 ;
  assign n97 = n96 ^ n95 ;
  assign n98 = n97 ^ n90 ;
  assign n99 = n98 ^ n96 ;
  assign n107 = n93 ^ n90 ;
  assign n101 = n90 ^ n77 ;
  assign n102 = n101 ^ n96 ;
  assign n103 = n102 ^ n74 ;
  assign n108 = n107 ^ n103 ;
  assign n109 = ~n99 & n108 ;
  assign n100 = n99 ^ n96 ;
  assign n104 = n103 ^ n93 ;
  assign n105 = n104 ^ n99 ;
  assign n106 = ~n100 & ~n105 ;
  assign n110 = n109 ^ n106 ;
  assign n111 = n110 ^ n93 ;
  assign n112 = n111 ^ n94 ;
  assign n113 = n112 ^ n103 ;
  assign n114 = n109 ^ n96 ;
  assign n115 = n107 ^ n94 ;
  assign n116 = n115 ^ n96 ;
  assign n117 = n107 ^ n96 ;
  assign n118 = n117 ^ n99 ;
  assign n119 = ~n116 & n118 ;
  assign n120 = n119 ^ n90 ;
  assign n121 = n120 ^ n93 ;
  assign n122 = n121 ^ n96 ;
  assign n123 = n122 ^ n103 ;
  assign n124 = n123 ^ n99 ;
  assign n125 = n114 & ~n124 ;
  assign n126 = n125 ^ n93 ;
  assign n127 = n126 ^ n99 ;
  assign n128 = n113 & n127 ;
  assign n129 = n128 ^ n109 ;
  assign n130 = n129 ^ n119 ;
  assign n131 = n130 ^ n106 ;
  assign n132 = n131 ^ n125 ;
  assign n133 = n132 ^ n90 ;
  assign n134 = n133 ^ n96 ;
  assign n135 = n134 ^ n103 ;
  assign n136 = n135 ^ n99 ;
  assign n137 = n136 ^ x3 ;
  assign n138 = n137 ^ n97 ;
  assign n139 = n138 ^ n71 ;
  assign n140 = n73 & ~n139 ;
  assign n141 = n140 ^ n71 ;
  assign n142 = ~n12 & n141 ;
  assign n143 = ~x0 & ~n142 ;
  assign n144 = x6 & x7 ;
  assign n145 = x0 & x1 ;
  assign n146 = ~n144 & ~n145 ;
  assign n147 = x1 & x6 ;
  assign n148 = ~x4 & n10 ;
  assign n149 = ~n147 & n148 ;
  assign n150 = ~n146 & n149 ;
  assign n151 = ~x3 & n150 ;
  assign n152 = ~n143 & ~n151 ;
  assign y0 = ~n152 ;
endmodule
