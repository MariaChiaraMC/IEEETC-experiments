module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 ;
  assign n9 = x1 & x4 ;
  assign n10 = ~x3 & n9 ;
  assign n11 = ~x6 & ~x7 ;
  assign n12 = ~x2 & n11 ;
  assign n13 = n12 ^ x5 ;
  assign n14 = n13 ^ n10 ;
  assign n15 = x6 & x7 ;
  assign n16 = ~x0 & x2 ;
  assign n17 = n15 & n16 ;
  assign n18 = n17 ^ x0 ;
  assign n19 = ~x5 & n18 ;
  assign n20 = n19 ^ x0 ;
  assign n21 = ~n14 & ~n20 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ x0 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = n10 & n24 ;
  assign n26 = ~x6 & x7 ;
  assign n27 = x0 & x5 ;
  assign n28 = x2 & n27 ;
  assign n29 = n26 & n28 ;
  assign n30 = ~x3 & n29 ;
  assign n42 = ~x5 & ~x7 ;
  assign n43 = x6 & n42 ;
  assign n44 = x2 & ~n43 ;
  assign n31 = ~x3 & x5 ;
  assign n32 = n15 & n31 ;
  assign n33 = n32 ^ n11 ;
  assign n34 = n33 ^ n32 ;
  assign n35 = x3 & ~x5 ;
  assign n36 = n35 ^ n32 ;
  assign n37 = n36 ^ n32 ;
  assign n38 = n34 & n37 ;
  assign n39 = n38 ^ n32 ;
  assign n40 = x2 & n39 ;
  assign n41 = n40 ^ n32 ;
  assign n45 = n44 ^ n41 ;
  assign n46 = n45 ^ n41 ;
  assign n47 = x3 & x5 ;
  assign n48 = n26 & n47 ;
  assign n49 = ~x2 & x3 ;
  assign n50 = n42 & ~n49 ;
  assign n51 = ~n48 & ~n50 ;
  assign n52 = n51 ^ n41 ;
  assign n53 = n52 ^ n41 ;
  assign n54 = ~n46 & ~n53 ;
  assign n55 = n54 ^ n41 ;
  assign n56 = x0 & n55 ;
  assign n57 = n56 ^ n41 ;
  assign n58 = x1 & n57 ;
  assign n59 = n16 ^ x3 ;
  assign n60 = x6 ^ x5 ;
  assign n61 = n60 ^ x5 ;
  assign n62 = x2 & x5 ;
  assign n63 = n62 ^ x5 ;
  assign n64 = n61 & ~n63 ;
  assign n65 = n64 ^ x5 ;
  assign n66 = n65 ^ n16 ;
  assign n67 = ~n59 & n66 ;
  assign n68 = n67 ^ n64 ;
  assign n69 = n68 ^ x5 ;
  assign n70 = n69 ^ x3 ;
  assign n71 = ~n16 & ~n70 ;
  assign n72 = n71 ^ n16 ;
  assign n73 = n72 ^ x7 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = n74 ^ x1 ;
  assign n76 = x5 & ~x6 ;
  assign n77 = ~n49 & ~n76 ;
  assign n78 = x0 & ~n77 ;
  assign n79 = ~n47 & n78 ;
  assign n80 = ~x2 & ~x3 ;
  assign n81 = ~x0 & x6 ;
  assign n82 = ~n80 & n81 ;
  assign n83 = x5 ^ x3 ;
  assign n84 = n82 & ~n83 ;
  assign n85 = n84 ^ n79 ;
  assign n86 = ~n79 & n85 ;
  assign n87 = n86 ^ n72 ;
  assign n88 = n87 ^ n79 ;
  assign n89 = ~n75 & ~n88 ;
  assign n90 = n89 ^ n86 ;
  assign n91 = n90 ^ n79 ;
  assign n92 = ~x1 & ~n91 ;
  assign n93 = n92 ^ x1 ;
  assign n94 = ~n58 & n93 ;
  assign n95 = ~n30 & n94 ;
  assign n96 = n95 ^ x1 ;
  assign n97 = n96 ^ x4 ;
  assign n106 = n97 ^ n96 ;
  assign n98 = n12 & n27 ;
  assign n99 = ~x3 & n98 ;
  assign n100 = n99 ^ n97 ;
  assign n101 = n100 ^ n96 ;
  assign n102 = n97 ^ n95 ;
  assign n103 = n102 ^ n99 ;
  assign n104 = n103 ^ n101 ;
  assign n105 = n101 & n104 ;
  assign n107 = n106 ^ n105 ;
  assign n108 = n107 ^ n101 ;
  assign n113 = ~x2 & x5 ;
  assign n110 = n26 & ~n62 ;
  assign n114 = n113 ^ n110 ;
  assign n115 = n114 ^ n110 ;
  assign n109 = x7 ^ x2 ;
  assign n111 = n110 ^ n109 ;
  assign n112 = n111 ^ n110 ;
  assign n116 = n115 ^ n112 ;
  assign n117 = n110 ^ x6 ;
  assign n118 = n117 ^ n110 ;
  assign n119 = n118 ^ n115 ;
  assign n120 = ~n115 & ~n119 ;
  assign n121 = n120 ^ n115 ;
  assign n122 = n116 & ~n121 ;
  assign n123 = n122 ^ n120 ;
  assign n124 = n123 ^ n110 ;
  assign n125 = n124 ^ n115 ;
  assign n126 = x0 & ~n125 ;
  assign n127 = n126 ^ n110 ;
  assign n128 = x3 & n127 ;
  assign n129 = n81 & n109 ;
  assign n130 = n31 & n129 ;
  assign n131 = ~n128 & ~n130 ;
  assign n132 = n131 ^ n96 ;
  assign n133 = n105 ^ n101 ;
  assign n134 = n132 & n133 ;
  assign n135 = n134 ^ n96 ;
  assign n136 = ~n108 & n135 ;
  assign n137 = n136 ^ n96 ;
  assign n138 = n137 ^ x1 ;
  assign n139 = n138 ^ n96 ;
  assign n140 = ~n25 & n139 ;
  assign y0 = ~n140 ;
endmodule
