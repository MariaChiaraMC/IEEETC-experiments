module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 ;
  assign n9 = x7 ^ x6 ;
  assign n10 = x4 & ~n9 ;
  assign n11 = ~x5 & ~n10 ;
  assign n12 = x3 & ~n11 ;
  assign n13 = x6 & x7 ;
  assign n14 = ~x4 & ~n13 ;
  assign n15 = ~x2 & ~x5 ;
  assign n16 = ~n14 & ~n15 ;
  assign n17 = x4 ^ x2 ;
  assign n18 = n17 ^ x3 ;
  assign n19 = n18 ^ x6 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = n18 ^ x3 ;
  assign n22 = n21 ^ x2 ;
  assign n23 = n20 & n22 ;
  assign n24 = n23 ^ x3 ;
  assign n25 = ~x3 & ~x5 ;
  assign n26 = n25 ^ x2 ;
  assign n27 = ~n24 & n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = x2 & n28 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = n30 ^ x3 ;
  assign n32 = n31 ^ x3 ;
  assign n33 = n16 & ~n32 ;
  assign n34 = ~n12 & n33 ;
  assign n48 = x5 & n13 ;
  assign n49 = ~n14 & ~n48 ;
  assign n50 = x2 & x3 ;
  assign n51 = ~n49 & n50 ;
  assign n35 = x5 & ~x7 ;
  assign n36 = ~x2 & n35 ;
  assign n52 = x6 & n36 ;
  assign n53 = ~x3 & n52 ;
  assign n54 = x2 & ~x3 ;
  assign n55 = n54 ^ x4 ;
  assign n56 = n55 ^ n54 ;
  assign n57 = n56 ^ n53 ;
  assign n58 = ~x5 & x6 ;
  assign n59 = x3 & x7 ;
  assign n60 = x5 & ~x6 ;
  assign n61 = n59 & ~n60 ;
  assign n62 = ~n58 & ~n61 ;
  assign n63 = n58 & n59 ;
  assign n64 = x2 & ~n63 ;
  assign n65 = ~n62 & n64 ;
  assign n66 = n13 ^ x3 ;
  assign n67 = x5 & ~n66 ;
  assign n68 = n67 ^ x3 ;
  assign n69 = ~x2 & n68 ;
  assign n70 = n69 ^ n65 ;
  assign n71 = ~n65 & n70 ;
  assign n72 = n71 ^ n54 ;
  assign n73 = n72 ^ n65 ;
  assign n74 = ~n57 & ~n73 ;
  assign n75 = n74 ^ n71 ;
  assign n76 = n75 ^ n65 ;
  assign n77 = ~n53 & ~n76 ;
  assign n78 = n77 ^ n53 ;
  assign n79 = ~n51 & ~n78 ;
  assign n37 = x2 & ~x7 ;
  assign n38 = ~n9 & ~n37 ;
  assign n39 = ~x5 & ~n38 ;
  assign n40 = ~n36 & ~n39 ;
  assign n41 = n40 ^ x3 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = n37 ^ x6 ;
  assign n44 = n43 ^ n40 ;
  assign n45 = ~n42 & n44 ;
  assign n46 = n45 ^ n40 ;
  assign n47 = ~x4 & n46 ;
  assign n80 = n79 ^ n47 ;
  assign n81 = n80 ^ n79 ;
  assign n82 = n60 ^ n59 ;
  assign n83 = n60 ^ n37 ;
  assign n84 = n83 ^ n37 ;
  assign n85 = n58 ^ n37 ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = n86 ^ n37 ;
  assign n88 = n82 & n87 ;
  assign n89 = n88 ^ n59 ;
  assign n90 = ~n52 & ~n89 ;
  assign n91 = x7 ^ x3 ;
  assign n92 = n15 & n91 ;
  assign n93 = n90 & ~n92 ;
  assign n94 = x4 & n93 ;
  assign n95 = n94 ^ n79 ;
  assign n96 = n95 ^ n79 ;
  assign n97 = ~n81 & ~n96 ;
  assign n98 = n97 ^ n79 ;
  assign n99 = ~x1 & ~n98 ;
  assign n100 = n99 ^ n79 ;
  assign n101 = ~n34 & n100 ;
  assign n102 = ~x0 & ~n101 ;
  assign y0 = n102 ;
endmodule
