module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n7 = x5 ^ x3 ;
  assign n8 = ~x1 & x4 ;
  assign n9 = n8 ^ x0 ;
  assign n10 = n8 ^ x3 ;
  assign n11 = n8 ^ x2 ;
  assign n12 = n8 & ~n11 ;
  assign n13 = n12 ^ n8 ;
  assign n14 = n10 & n13 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n15 ^ n8 ;
  assign n17 = n16 ^ x2 ;
  assign n18 = n9 & ~n17 ;
  assign n19 = n18 ^ x0 ;
  assign n20 = n19 ^ n7 ;
  assign n21 = x1 & ~x4 ;
  assign n22 = n21 ^ x3 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = x0 & ~x1 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = ~n23 & n25 ;
  assign n27 = n26 ^ n21 ;
  assign n28 = n27 ^ n7 ;
  assign n29 = ~n20 & n28 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n30 ^ n21 ;
  assign n32 = n31 ^ n19 ;
  assign n33 = ~n7 & ~n32 ;
  assign n34 = n33 ^ n7 ;
  assign y0 = ~n34 ;
endmodule
