module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 ;
  assign n10 = x4 & x8 ;
  assign n11 = ~x6 & ~x7 ;
  assign n12 = ~x1 & ~x3 ;
  assign n13 = n11 & n12 ;
  assign n14 = n10 & n13 ;
  assign n15 = x1 & x7 ;
  assign n16 = x8 ^ x4 ;
  assign n17 = n15 & ~n16 ;
  assign n18 = n17 ^ x6 ;
  assign n19 = n18 ^ n17 ;
  assign n20 = n19 ^ n14 ;
  assign n21 = ~x7 & x8 ;
  assign n22 = x7 & ~x8 ;
  assign n23 = ~x1 & n22 ;
  assign n24 = ~n21 & ~n23 ;
  assign n25 = ~x3 & ~x4 ;
  assign n26 = n25 ^ n24 ;
  assign n27 = ~n24 & ~n26 ;
  assign n28 = n27 ^ n17 ;
  assign n29 = n28 ^ n24 ;
  assign n30 = ~n20 & ~n29 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n31 ^ n24 ;
  assign n33 = ~n14 & ~n32 ;
  assign n34 = n33 ^ n14 ;
  assign n35 = ~x5 & n34 ;
  assign n36 = x5 & n25 ;
  assign n37 = n11 & n36 ;
  assign n50 = x3 & ~x6 ;
  assign n38 = x3 & x8 ;
  assign n39 = x5 & ~x7 ;
  assign n40 = n39 ^ x5 ;
  assign n41 = n40 ^ n39 ;
  assign n42 = x6 & x7 ;
  assign n43 = n42 ^ n39 ;
  assign n44 = n43 ^ n39 ;
  assign n45 = ~n41 & n44 ;
  assign n46 = n45 ^ n39 ;
  assign n47 = ~x4 & n46 ;
  assign n48 = n47 ^ n39 ;
  assign n49 = n38 & n48 ;
  assign n51 = n50 ^ n49 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = x4 & ~x8 ;
  assign n54 = n39 & n53 ;
  assign n55 = x5 & x8 ;
  assign n56 = ~x4 & x7 ;
  assign n57 = ~n55 & n56 ;
  assign n58 = ~n54 & ~n57 ;
  assign n59 = n58 ^ n49 ;
  assign n60 = n59 ^ n49 ;
  assign n61 = n52 & ~n60 ;
  assign n62 = n61 ^ n49 ;
  assign n63 = ~x1 & n62 ;
  assign n64 = n63 ^ n49 ;
  assign n65 = ~n37 & ~n64 ;
  assign n66 = ~x5 & ~x7 ;
  assign n67 = ~x1 & n50 ;
  assign n68 = n67 ^ x3 ;
  assign n69 = n68 ^ x8 ;
  assign n78 = n69 ^ n68 ;
  assign n70 = ~x4 & x6 ;
  assign n71 = ~x1 & n70 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = n72 ^ n68 ;
  assign n74 = n69 ^ n67 ;
  assign n75 = n74 ^ n71 ;
  assign n76 = n75 ^ n73 ;
  assign n77 = n73 & ~n76 ;
  assign n79 = n78 ^ n77 ;
  assign n80 = n79 ^ n73 ;
  assign n81 = x4 & ~x6 ;
  assign n82 = n81 ^ n68 ;
  assign n83 = n77 ^ n73 ;
  assign n84 = ~n82 & n83 ;
  assign n85 = n84 ^ n68 ;
  assign n86 = ~n80 & n85 ;
  assign n87 = n86 ^ n68 ;
  assign n88 = n87 ^ x3 ;
  assign n89 = n88 ^ n68 ;
  assign n90 = n66 & n89 ;
  assign n91 = x4 & n42 ;
  assign n92 = x7 & n50 ;
  assign n93 = ~n91 & ~n92 ;
  assign n94 = ~x5 & ~x8 ;
  assign n95 = ~n93 & n94 ;
  assign n96 = ~x6 & x7 ;
  assign n97 = ~x5 & n96 ;
  assign n98 = x8 & n97 ;
  assign n99 = x6 ^ x4 ;
  assign n102 = n99 ^ x6 ;
  assign n103 = n102 ^ x8 ;
  assign n100 = n99 ^ x8 ;
  assign n101 = n100 ^ x5 ;
  assign n104 = n103 ^ n101 ;
  assign n105 = n104 ^ x7 ;
  assign n106 = ~x7 & ~n105 ;
  assign n107 = n106 ^ n99 ;
  assign n108 = n107 ^ x7 ;
  assign n109 = x5 & n103 ;
  assign n110 = n109 ^ n99 ;
  assign n111 = n108 & ~n110 ;
  assign n112 = n111 ^ n99 ;
  assign n113 = n112 ^ x5 ;
  assign n114 = ~n98 & n113 ;
  assign n115 = ~x3 & ~n114 ;
  assign n116 = ~n95 & ~n115 ;
  assign n117 = x1 & ~n116 ;
  assign n118 = ~x1 & x8 ;
  assign n119 = x6 & ~n66 ;
  assign n120 = x3 & n119 ;
  assign n121 = x7 & n81 ;
  assign n122 = x5 & n121 ;
  assign n123 = ~n120 & ~n122 ;
  assign n124 = n118 & ~n123 ;
  assign n125 = ~x4 & ~x8 ;
  assign n126 = ~n42 & ~n66 ;
  assign n127 = n125 & n126 ;
  assign n128 = n11 & n55 ;
  assign n129 = ~n127 & ~n128 ;
  assign n130 = ~x3 & ~n129 ;
  assign n133 = x1 & n11 ;
  assign n131 = ~x3 & x8 ;
  assign n132 = ~x4 & ~n131 ;
  assign n134 = n133 ^ n132 ;
  assign n135 = ~x8 & n42 ;
  assign n136 = n135 ^ n132 ;
  assign n137 = x3 & x5 ;
  assign n138 = n137 ^ n133 ;
  assign n139 = n138 ^ n135 ;
  assign n140 = ~n135 & ~n139 ;
  assign n141 = n140 ^ n135 ;
  assign n142 = ~n136 & ~n141 ;
  assign n143 = n142 ^ n140 ;
  assign n144 = n143 ^ n135 ;
  assign n145 = n144 ^ n138 ;
  assign n146 = n134 & ~n145 ;
  assign n147 = n146 ^ n133 ;
  assign n148 = ~n130 & ~n147 ;
  assign n149 = ~n124 & n148 ;
  assign n150 = ~n117 & n149 ;
  assign n151 = ~n90 & n150 ;
  assign n152 = n151 ^ x2 ;
  assign n153 = n152 ^ n151 ;
  assign n159 = ~n39 & ~n81 ;
  assign n157 = x8 ^ x1 ;
  assign n154 = ~x4 & n21 ;
  assign n155 = ~n135 & ~n154 ;
  assign n156 = n155 ^ x1 ;
  assign n158 = n157 ^ n156 ;
  assign n160 = n159 ^ n158 ;
  assign n161 = n160 ^ n158 ;
  assign n162 = n158 ^ n156 ;
  assign n163 = n162 ^ x1 ;
  assign n164 = ~n161 & ~n163 ;
  assign n165 = n164 ^ n156 ;
  assign n166 = n66 & ~n156 ;
  assign n167 = n166 ^ x1 ;
  assign n168 = ~n165 & n167 ;
  assign n169 = n168 ^ n166 ;
  assign n170 = x1 & n169 ;
  assign n171 = n170 ^ n164 ;
  assign n172 = n171 ^ n155 ;
  assign n173 = n172 ^ n156 ;
  assign n174 = x6 & n66 ;
  assign n175 = n174 ^ x8 ;
  assign n176 = ~x4 & ~x5 ;
  assign n177 = ~n91 & ~n176 ;
  assign n178 = ~x1 & ~n177 ;
  assign n179 = n178 ^ n131 ;
  assign n180 = ~n175 & n179 ;
  assign n181 = n180 ^ n178 ;
  assign n182 = n131 & n181 ;
  assign n183 = n182 ^ x3 ;
  assign n184 = ~n173 & ~n183 ;
  assign n185 = n96 ^ x8 ;
  assign n186 = n185 ^ n96 ;
  assign n187 = n96 ^ n66 ;
  assign n188 = n187 ^ n96 ;
  assign n189 = ~n186 & n188 ;
  assign n190 = n189 ^ n96 ;
  assign n191 = x4 & n190 ;
  assign n192 = n191 ^ n96 ;
  assign n193 = x1 & n192 ;
  assign n194 = x3 & ~n98 ;
  assign n195 = ~n193 & n194 ;
  assign n196 = ~n184 & ~n195 ;
  assign n197 = ~x4 & ~x7 ;
  assign n198 = n197 ^ n42 ;
  assign n199 = n198 ^ x8 ;
  assign n206 = n199 ^ n198 ;
  assign n200 = n199 ^ x1 ;
  assign n201 = n200 ^ n198 ;
  assign n202 = n197 ^ x1 ;
  assign n203 = n202 ^ x1 ;
  assign n204 = n203 ^ n201 ;
  assign n205 = n201 & n204 ;
  assign n207 = n206 ^ n205 ;
  assign n208 = n207 ^ n201 ;
  assign n209 = n198 ^ x6 ;
  assign n210 = n205 ^ n201 ;
  assign n211 = ~n209 & n210 ;
  assign n212 = n211 ^ n198 ;
  assign n213 = n208 & n212 ;
  assign n214 = n213 ^ n198 ;
  assign n215 = n214 ^ n197 ;
  assign n216 = n215 ^ n198 ;
  assign n217 = n137 & n216 ;
  assign n218 = n154 ^ x6 ;
  assign n219 = n218 ^ n154 ;
  assign n220 = n15 & n53 ;
  assign n221 = n220 ^ n154 ;
  assign n222 = n219 & n221 ;
  assign n223 = n222 ^ n154 ;
  assign n224 = x5 & n223 ;
  assign n225 = ~n217 & ~n224 ;
  assign n226 = ~n196 & n225 ;
  assign n227 = n226 ^ n151 ;
  assign n228 = n153 & n227 ;
  assign n229 = n228 ^ n151 ;
  assign n230 = n65 & n229 ;
  assign n231 = ~n35 & n230 ;
  assign n232 = ~x0 & ~n231 ;
  assign n233 = x0 & n94 ;
  assign n234 = n42 & n55 ;
  assign n235 = ~n233 & ~n234 ;
  assign n236 = ~x4 & ~n235 ;
  assign n237 = n10 & n96 ;
  assign n238 = x4 & n119 ;
  assign n239 = ~n54 & ~n238 ;
  assign n240 = ~n97 & n239 ;
  assign n241 = x0 & ~n240 ;
  assign n242 = ~n237 & ~n241 ;
  assign n243 = ~n236 & n242 ;
  assign n244 = n12 & ~n243 ;
  assign n245 = ~x2 & n244 ;
  assign n246 = ~n232 & ~n245 ;
  assign y0 = ~n246 ;
endmodule
