module top( x0 , x1 , x2 , x3 , x4 , y0 );
  input x0 , x1 , x2 , x3 , x4 ;
  output y0 ;
  wire n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 ;
  assign n6 = x4 ^ x3 ;
  assign n7 = x1 ^ x0 ;
  assign n8 = n7 ^ n6 ;
  assign n9 = x2 ^ x1 ;
  assign n10 = n9 ^ x1 ;
  assign n11 = x4 ^ x1 ;
  assign n12 = ~n10 & ~n11 ;
  assign n13 = n12 ^ x1 ;
  assign n14 = n13 ^ n6 ;
  assign n15 = ~n8 & ~n14 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = n16 ^ x1 ;
  assign n18 = n17 ^ n7 ;
  assign n19 = n6 & n18 ;
  assign n20 = n19 ^ n6 ;
  assign y0 = n20 ;
endmodule
