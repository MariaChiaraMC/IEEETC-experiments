module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n8 = ~x2 & ~x3 ;
  assign n9 = ~x1 & n8 ;
  assign n12 = ~x5 & ~x6 ;
  assign n13 = n12 ^ x3 ;
  assign n14 = n13 ^ x4 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = n15 ^ x3 ;
  assign n18 = n16 ^ x3 ;
  assign n10 = x3 ^ x1 ;
  assign n11 = ~x0 & n10 ;
  assign n17 = n16 ^ n11 ;
  assign n19 = n18 ^ n17 ;
  assign n22 = n13 ^ x3 ;
  assign n20 = n18 ^ n16 ;
  assign n21 = x2 & n20 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = ~n18 & ~n23 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n19 & n25 ;
  assign n27 = n26 ^ n21 ;
  assign n28 = n27 ^ n11 ;
  assign n29 = n28 ^ n24 ;
  assign n30 = n29 ^ x3 ;
  assign n31 = ~n9 & ~n30 ;
  assign y0 = ~n31 ;
endmodule
