module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 ;
  assign n15 = x2 & ~x12 ;
  assign n16 = x9 & n15 ;
  assign n17 = ~x7 & ~x10 ;
  assign n18 = ~x8 & ~x11 ;
  assign n19 = n17 & n18 ;
  assign n20 = x5 & ~x13 ;
  assign n21 = n19 & n20 ;
  assign n22 = n16 & n21 ;
  assign n23 = x3 & ~n22 ;
  assign n24 = x4 ^ x0 ;
  assign n25 = ~x3 & x5 ;
  assign n26 = x1 & ~n25 ;
  assign n27 = n26 ^ x6 ;
  assign n28 = n27 ^ n26 ;
  assign n29 = ~x1 & ~x3 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = ~n28 & n30 ;
  assign n32 = n31 ^ n26 ;
  assign n33 = n32 ^ x4 ;
  assign n34 = ~n24 & n33 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = n35 ^ n26 ;
  assign n37 = n36 ^ x0 ;
  assign n38 = x4 & ~n37 ;
  assign n39 = n38 ^ x4 ;
  assign n40 = ~n23 & n39 ;
  assign y0 = n40 ;
endmodule
