module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 ;
  assign n9 = x0 & ~x2 ;
  assign n10 = x1 & x7 ;
  assign n11 = ~x4 & n10 ;
  assign n12 = x3 & ~x6 ;
  assign n13 = n11 & n12 ;
  assign n14 = n9 & n13 ;
  assign n15 = x3 & ~x7 ;
  assign n16 = ~x0 & ~x3 ;
  assign n17 = x6 & n16 ;
  assign n18 = ~n15 & ~n17 ;
  assign n19 = ~x2 & ~n18 ;
  assign n20 = n15 ^ x0 ;
  assign n21 = ~x3 & x7 ;
  assign n22 = n21 ^ n15 ;
  assign n23 = n21 ^ x6 ;
  assign n24 = ~n21 & ~n23 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n22 & ~n25 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = n28 ^ x6 ;
  assign n30 = n20 & ~n29 ;
  assign n31 = n30 ^ n15 ;
  assign n32 = ~n19 & ~n31 ;
  assign n35 = n32 ^ x6 ;
  assign n36 = n35 ^ n32 ;
  assign n33 = n32 ^ n16 ;
  assign n34 = n33 ^ n32 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = x7 ^ x2 ;
  assign n39 = n38 ^ n32 ;
  assign n40 = n39 ^ n32 ;
  assign n41 = n40 ^ n36 ;
  assign n42 = ~n36 & n41 ;
  assign n43 = n42 ^ n36 ;
  assign n44 = ~n37 & ~n43 ;
  assign n45 = n44 ^ n42 ;
  assign n46 = n45 ^ n32 ;
  assign n47 = n46 ^ n36 ;
  assign n48 = ~x1 & n47 ;
  assign n49 = n48 ^ n32 ;
  assign n50 = ~x4 & ~n49 ;
  assign n51 = ~x1 & x6 ;
  assign n52 = x3 & n51 ;
  assign n53 = x7 & n52 ;
  assign n54 = ~x0 & x4 ;
  assign n55 = ~x0 & ~x2 ;
  assign n56 = ~n54 & ~n55 ;
  assign n57 = n53 & ~n56 ;
  assign n58 = ~x2 & ~x3 ;
  assign n59 = x4 & n58 ;
  assign n60 = x0 & ~x1 ;
  assign n61 = x6 & ~x7 ;
  assign n62 = n60 & n61 ;
  assign n63 = n59 & n62 ;
  assign n64 = x2 & ~x6 ;
  assign n65 = x7 ^ x3 ;
  assign n66 = n65 ^ x3 ;
  assign n67 = x3 ^ x1 ;
  assign n68 = ~n66 & ~n67 ;
  assign n69 = n68 ^ x3 ;
  assign n70 = n64 & n69 ;
  assign n71 = n54 & n70 ;
  assign n72 = ~n63 & ~n71 ;
  assign n73 = ~n57 & n72 ;
  assign n74 = ~n50 & n73 ;
  assign n75 = n74 ^ x5 ;
  assign n76 = n75 ^ n74 ;
  assign n77 = n58 ^ x3 ;
  assign n78 = n77 ^ n58 ;
  assign n79 = n58 ^ x0 ;
  assign n80 = n79 ^ n58 ;
  assign n81 = n78 & ~n80 ;
  assign n82 = n81 ^ n58 ;
  assign n83 = ~x7 & n82 ;
  assign n84 = n83 ^ n58 ;
  assign n85 = ~n54 & n84 ;
  assign n86 = n51 & n85 ;
  assign n87 = ~x1 & ~n9 ;
  assign n88 = x4 & ~n87 ;
  assign n89 = ~x0 & x2 ;
  assign n90 = n89 ^ x7 ;
  assign n92 = n90 ^ n55 ;
  assign n93 = n92 ^ n90 ;
  assign n91 = n90 ^ n89 ;
  assign n94 = n93 ^ n91 ;
  assign n95 = n90 ^ x1 ;
  assign n96 = n95 ^ n90 ;
  assign n97 = n96 ^ n93 ;
  assign n98 = n93 & n97 ;
  assign n99 = n98 ^ n93 ;
  assign n100 = n94 & n99 ;
  assign n101 = n100 ^ n98 ;
  assign n102 = n101 ^ n90 ;
  assign n103 = n102 ^ n93 ;
  assign n104 = ~x3 & ~n103 ;
  assign n105 = n104 ^ n90 ;
  assign n106 = n88 & ~n105 ;
  assign n107 = n106 ^ x6 ;
  assign n108 = n107 ^ n106 ;
  assign n109 = ~x2 & ~x7 ;
  assign n110 = n16 & n109 ;
  assign n111 = x3 ^ x2 ;
  assign n112 = n60 & n111 ;
  assign n113 = x7 & n112 ;
  assign n114 = ~n110 & ~n113 ;
  assign n115 = x4 & ~n114 ;
  assign n116 = ~x7 & n89 ;
  assign n117 = x2 & x3 ;
  assign n118 = x4 & ~n58 ;
  assign n119 = ~n117 & ~n118 ;
  assign n120 = x0 & n21 ;
  assign n121 = n120 ^ x3 ;
  assign n122 = n119 & n121 ;
  assign n123 = ~n116 & ~n122 ;
  assign n124 = x1 & ~n123 ;
  assign n125 = n124 ^ n60 ;
  assign n126 = n125 ^ n15 ;
  assign n127 = n126 ^ n125 ;
  assign n128 = n127 ^ x4 ;
  assign n129 = n124 ^ n58 ;
  assign n130 = n58 & n129 ;
  assign n131 = n130 ^ n125 ;
  assign n132 = n131 ^ n58 ;
  assign n133 = n128 & n132 ;
  assign n134 = n133 ^ n130 ;
  assign n135 = n134 ^ n58 ;
  assign n136 = ~x4 & n135 ;
  assign n137 = n136 ^ n124 ;
  assign n138 = ~n115 & ~n137 ;
  assign n139 = n138 ^ n106 ;
  assign n140 = ~n108 & ~n139 ;
  assign n141 = n140 ^ n106 ;
  assign n142 = ~n86 & ~n141 ;
  assign n143 = n142 ^ n74 ;
  assign n144 = ~n76 & n143 ;
  assign n145 = n144 ^ n74 ;
  assign n146 = ~n14 & n145 ;
  assign y0 = ~n146 ;
endmodule
