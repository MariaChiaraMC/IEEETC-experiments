module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 ;
  assign n22 = x1 & ~x3 ;
  assign n23 = ~x0 & ~x4 ;
  assign n24 = ~x2 & n23 ;
  assign n25 = n22 & n24 ;
  assign n26 = x1 & ~x2 ;
  assign n27 = ~x2 & ~x3 ;
  assign n28 = x0 & ~n27 ;
  assign n29 = ~n26 & ~n28 ;
  assign n30 = x0 & x1 ;
  assign n31 = ~x4 & ~n30 ;
  assign n32 = x5 & n31 ;
  assign n33 = ~n29 & n32 ;
  assign n34 = n33 ^ x14 ;
  assign n185 = ~x19 & ~x20 ;
  assign n35 = ~x12 & ~x13 ;
  assign n36 = x8 & x9 ;
  assign n37 = x10 & ~x11 ;
  assign n38 = n36 & n37 ;
  assign n39 = ~x4 & n38 ;
  assign n40 = n30 & n39 ;
  assign n41 = x2 & n40 ;
  assign n42 = ~x6 & ~x7 ;
  assign n43 = ~x0 & ~x1 ;
  assign n44 = ~x10 & x11 ;
  assign n45 = n36 & n44 ;
  assign n46 = ~x8 & n37 ;
  assign n47 = ~n45 & ~n46 ;
  assign n48 = ~n43 & ~n47 ;
  assign n49 = n42 & n48 ;
  assign n50 = n49 ^ n23 ;
  assign n51 = n49 ^ x1 ;
  assign n52 = n51 ^ n50 ;
  assign n53 = ~x8 & x9 ;
  assign n54 = ~x11 & n53 ;
  assign n55 = n42 & n54 ;
  assign n56 = n55 ^ x2 ;
  assign n57 = ~x1 & n56 ;
  assign n58 = n57 ^ n55 ;
  assign n59 = n52 & ~n58 ;
  assign n60 = n59 ^ n57 ;
  assign n61 = n60 ^ n55 ;
  assign n62 = n61 ^ x1 ;
  assign n63 = n50 & n62 ;
  assign n64 = n63 ^ n23 ;
  assign n65 = ~n41 & ~n64 ;
  assign n66 = n35 & ~n65 ;
  assign n67 = n23 ^ x5 ;
  assign n68 = n67 ^ x2 ;
  assign n101 = n68 ^ n67 ;
  assign n69 = x11 & ~x12 ;
  assign n70 = n53 & n69 ;
  assign n71 = n43 & ~n70 ;
  assign n72 = ~n30 & ~n71 ;
  assign n73 = x4 & ~n72 ;
  assign n74 = x13 & n54 ;
  assign n75 = ~x10 & n74 ;
  assign n76 = x10 & ~x12 ;
  assign n77 = n76 ^ x13 ;
  assign n78 = x9 & x11 ;
  assign n79 = n78 ^ n76 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = ~x1 & x2 ;
  assign n83 = ~x1 & x12 ;
  assign n84 = n83 ^ n82 ;
  assign n85 = ~n82 & n84 ;
  assign n86 = n85 ^ n78 ;
  assign n87 = n86 ^ n82 ;
  assign n88 = ~n81 & n87 ;
  assign n89 = n88 ^ n85 ;
  assign n90 = n89 ^ n82 ;
  assign n91 = n77 & ~n90 ;
  assign n92 = n91 ^ n76 ;
  assign n93 = ~n75 & ~n92 ;
  assign n94 = n73 & n93 ;
  assign n95 = n94 ^ n68 ;
  assign n96 = n95 ^ n67 ;
  assign n97 = n68 ^ n23 ;
  assign n98 = n97 ^ n94 ;
  assign n99 = n98 ^ n96 ;
  assign n100 = ~n96 & ~n99 ;
  assign n102 = n101 ^ n100 ;
  assign n103 = n102 ^ n96 ;
  assign n104 = ~x6 & ~x17 ;
  assign n105 = x12 & ~x13 ;
  assign n106 = n104 & ~n105 ;
  assign n107 = ~x8 & n106 ;
  assign n108 = ~x9 & ~x15 ;
  assign n109 = n108 ^ x7 ;
  assign n110 = n108 ^ x13 ;
  assign n111 = n110 ^ n109 ;
  assign n112 = x11 ^ x10 ;
  assign n113 = x13 & n112 ;
  assign n114 = n113 ^ x10 ;
  assign n115 = n111 & n114 ;
  assign n116 = n115 ^ n113 ;
  assign n117 = n116 ^ x10 ;
  assign n118 = n117 ^ x13 ;
  assign n119 = ~n109 & n118 ;
  assign n120 = n119 ^ x7 ;
  assign n121 = n107 & ~n120 ;
  assign n122 = x12 ^ x11 ;
  assign n123 = n122 ^ x12 ;
  assign n129 = ~x10 & x16 ;
  assign n125 = ~x10 & ~x13 ;
  assign n126 = ~x9 & n125 ;
  assign n130 = n129 ^ n126 ;
  assign n124 = n123 ^ x12 ;
  assign n127 = n126 ^ n123 ;
  assign n128 = n124 & ~n127 ;
  assign n131 = n130 ^ n128 ;
  assign n132 = ~n123 & n131 ;
  assign n133 = n132 ^ n129 ;
  assign n134 = n133 ^ n123 ;
  assign n135 = n121 & ~n134 ;
  assign n136 = n135 ^ n67 ;
  assign n137 = n100 ^ n96 ;
  assign n138 = n136 & ~n137 ;
  assign n139 = n138 ^ n67 ;
  assign n140 = n103 & n139 ;
  assign n141 = n140 ^ n67 ;
  assign n142 = n141 ^ x5 ;
  assign n143 = n142 ^ n67 ;
  assign n144 = ~n66 & ~n143 ;
  assign n145 = ~x3 & ~n144 ;
  assign n146 = x2 & x5 ;
  assign n147 = ~n38 & ~n55 ;
  assign n148 = n146 & ~n147 ;
  assign n149 = x5 & ~x9 ;
  assign n150 = ~x8 & n149 ;
  assign n151 = ~n37 & ~n44 ;
  assign n152 = n150 & ~n151 ;
  assign n153 = x3 & ~x5 ;
  assign n154 = n82 & n153 ;
  assign n155 = ~n26 & ~n154 ;
  assign n156 = n45 & ~n155 ;
  assign n157 = ~x0 & n156 ;
  assign n158 = ~n152 & ~n157 ;
  assign n159 = n42 & ~n158 ;
  assign n160 = ~n148 & ~n159 ;
  assign n161 = n35 & ~n160 ;
  assign n162 = ~x2 & x13 ;
  assign n163 = n150 & n162 ;
  assign n164 = n44 & n163 ;
  assign n165 = ~n161 & ~n164 ;
  assign n166 = ~x4 & ~n165 ;
  assign n167 = x4 & ~n22 ;
  assign n168 = ~x5 & ~n167 ;
  assign n169 = ~x0 & ~x5 ;
  assign n170 = n169 ^ x1 ;
  assign n171 = n170 ^ x1 ;
  assign n172 = n171 ^ n168 ;
  assign n173 = ~x3 & x5 ;
  assign n174 = ~n146 & ~n173 ;
  assign n175 = n174 ^ x2 ;
  assign n176 = x1 & ~n175 ;
  assign n177 = n176 ^ n174 ;
  assign n178 = n172 & n177 ;
  assign n179 = n178 ^ n176 ;
  assign n180 = n179 ^ n174 ;
  assign n181 = n180 ^ x1 ;
  assign n182 = ~n168 & n181 ;
  assign n183 = ~n166 & ~n182 ;
  assign n184 = ~n145 & n183 ;
  assign n186 = n185 ^ n184 ;
  assign n187 = n186 ^ n184 ;
  assign n188 = n184 ^ x18 ;
  assign n189 = ~n187 & n188 ;
  assign n190 = n189 ^ n184 ;
  assign n191 = n190 ^ n33 ;
  assign n192 = ~n34 & ~n191 ;
  assign n193 = n192 ^ n189 ;
  assign n194 = n193 ^ n184 ;
  assign n195 = n194 ^ x14 ;
  assign n196 = ~n33 & n195 ;
  assign n197 = n196 ^ n33 ;
  assign n198 = ~n25 & ~n197 ;
  assign y0 = ~n198 ;
endmodule
