module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 ;
  assign n11 = ~x4 & x7 ;
  assign n12 = x3 & x5 ;
  assign n13 = n11 & n12 ;
  assign n14 = x1 & x2 ;
  assign n15 = x8 & ~x9 ;
  assign n16 = n14 & n15 ;
  assign n17 = n13 & n16 ;
  assign n18 = ~x7 & x9 ;
  assign n19 = x3 & ~n18 ;
  assign n20 = x7 & ~x9 ;
  assign n21 = ~x3 & ~n20 ;
  assign n22 = x4 & ~x5 ;
  assign n23 = ~x8 & n22 ;
  assign n24 = ~x1 & ~x2 ;
  assign n25 = n23 & n24 ;
  assign n26 = ~n21 & n25 ;
  assign n27 = ~n19 & n26 ;
  assign n28 = ~n17 & ~n27 ;
  assign n29 = x5 & x9 ;
  assign n30 = x8 ^ x7 ;
  assign n31 = x7 ^ x4 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = x8 ^ x2 ;
  assign n34 = x3 ^ x2 ;
  assign n35 = n34 ^ x2 ;
  assign n36 = n33 & n35 ;
  assign n37 = n36 ^ x2 ;
  assign n38 = n37 ^ n30 ;
  assign n39 = ~n32 & n38 ;
  assign n40 = n39 ^ n36 ;
  assign n41 = n40 ^ x2 ;
  assign n42 = n41 ^ n31 ;
  assign n43 = n30 & ~n42 ;
  assign n44 = n43 ^ n30 ;
  assign n45 = n29 & n44 ;
  assign n46 = x5 ^ x2 ;
  assign n47 = ~x8 & x9 ;
  assign n48 = n11 & n47 ;
  assign n49 = x4 & x7 ;
  assign n50 = n15 & n49 ;
  assign n51 = x3 & n50 ;
  assign n52 = ~n48 & ~n51 ;
  assign n53 = n52 ^ x5 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = n54 ^ n46 ;
  assign n56 = ~x4 & ~x7 ;
  assign n57 = ~x9 & n56 ;
  assign n58 = x7 & x9 ;
  assign n59 = x3 & x4 ;
  assign n60 = n58 & n59 ;
  assign n61 = ~n57 & ~n60 ;
  assign n62 = n61 ^ x8 ;
  assign n63 = ~n61 & n62 ;
  assign n64 = n63 ^ n52 ;
  assign n65 = n64 ^ n61 ;
  assign n66 = ~n55 & n65 ;
  assign n67 = n66 ^ n63 ;
  assign n68 = n67 ^ n61 ;
  assign n69 = n46 & ~n68 ;
  assign n70 = ~n45 & ~n69 ;
  assign n71 = n70 ^ x1 ;
  assign n72 = n71 ^ n70 ;
  assign n73 = n72 ^ x0 ;
  assign n74 = x2 & ~x3 ;
  assign n75 = x4 & x9 ;
  assign n76 = n75 ^ x5 ;
  assign n77 = n76 ^ n74 ;
  assign n78 = n75 ^ x9 ;
  assign n79 = n78 ^ x8 ;
  assign n80 = ~x8 & n79 ;
  assign n81 = n80 ^ n75 ;
  assign n82 = n81 ^ x8 ;
  assign n83 = n77 & ~n82 ;
  assign n84 = n83 ^ n80 ;
  assign n85 = n84 ^ x8 ;
  assign n86 = n74 & ~n85 ;
  assign n87 = ~x7 & n86 ;
  assign n88 = x3 & ~x8 ;
  assign n89 = n57 & n88 ;
  assign n90 = n58 ^ x3 ;
  assign n91 = n90 ^ n58 ;
  assign n92 = x9 ^ x7 ;
  assign n93 = n31 & n92 ;
  assign n94 = n93 ^ n58 ;
  assign n95 = n94 ^ n58 ;
  assign n96 = n91 & n95 ;
  assign n97 = n96 ^ n58 ;
  assign n98 = ~x2 & n97 ;
  assign n99 = n98 ^ n58 ;
  assign n100 = x8 & n99 ;
  assign n101 = ~n89 & ~n100 ;
  assign n102 = ~x5 & ~n101 ;
  assign n103 = n102 ^ n87 ;
  assign n104 = ~n87 & n103 ;
  assign n105 = n104 ^ n70 ;
  assign n106 = n105 ^ n87 ;
  assign n107 = n73 & ~n106 ;
  assign n108 = n107 ^ n104 ;
  assign n109 = n108 ^ n87 ;
  assign n110 = x0 & ~n109 ;
  assign n111 = n110 ^ x0 ;
  assign n112 = n28 & ~n111 ;
  assign n113 = ~x6 & ~n112 ;
  assign n114 = ~x8 & ~x9 ;
  assign n115 = ~x3 & ~x4 ;
  assign n116 = n114 & n115 ;
  assign n117 = x5 & x7 ;
  assign n118 = x6 & n117 ;
  assign n119 = n116 & n118 ;
  assign n120 = n24 & n119 ;
  assign n121 = n120 ^ n113 ;
  assign n122 = ~x3 & x9 ;
  assign n123 = n49 & n122 ;
  assign n124 = ~x5 & x8 ;
  assign n125 = n14 & n124 ;
  assign n126 = n123 & n125 ;
  assign n127 = ~x5 & ~x7 ;
  assign n128 = ~x4 & n15 ;
  assign n129 = x3 & n128 ;
  assign n130 = x2 & ~x8 ;
  assign n131 = x2 & x4 ;
  assign n132 = ~x3 & n131 ;
  assign n133 = ~n116 & ~n132 ;
  assign n134 = ~n130 & ~n133 ;
  assign n135 = ~n129 & ~n134 ;
  assign n136 = n127 & ~n135 ;
  assign n137 = ~x7 & n15 ;
  assign n138 = x7 & ~x8 ;
  assign n139 = n122 & n138 ;
  assign n140 = ~n137 & ~n139 ;
  assign n141 = n131 & ~n140 ;
  assign n142 = n48 ^ x2 ;
  assign n143 = n142 ^ n48 ;
  assign n144 = n143 ^ x3 ;
  assign n145 = ~x7 & n75 ;
  assign n146 = n145 ^ n128 ;
  assign n147 = ~n145 & n146 ;
  assign n148 = n147 ^ n48 ;
  assign n149 = n148 ^ n145 ;
  assign n150 = ~n144 & n149 ;
  assign n151 = n150 ^ n147 ;
  assign n152 = n151 ^ n145 ;
  assign n153 = x3 & ~n152 ;
  assign n154 = n153 ^ x3 ;
  assign n155 = ~n141 & ~n154 ;
  assign n156 = x5 & ~n155 ;
  assign n157 = x1 & ~n156 ;
  assign n158 = ~n136 & n157 ;
  assign n159 = n88 & n117 ;
  assign n160 = n75 & n159 ;
  assign n161 = n12 & n93 ;
  assign n162 = ~n20 & ~n127 ;
  assign n163 = ~x5 & ~x9 ;
  assign n164 = ~x3 & ~n11 ;
  assign n165 = ~n163 & n164 ;
  assign n166 = ~n162 & n165 ;
  assign n167 = n166 ^ n13 ;
  assign n168 = n167 ^ x2 ;
  assign n175 = n168 ^ n167 ;
  assign n169 = n168 ^ n19 ;
  assign n170 = n169 ^ n167 ;
  assign n171 = n168 ^ n166 ;
  assign n172 = n171 ^ n19 ;
  assign n173 = n172 ^ n170 ;
  assign n174 = ~n170 & n173 ;
  assign n176 = n175 ^ n174 ;
  assign n177 = n176 ^ n170 ;
  assign n178 = x9 & n22 ;
  assign n179 = n178 ^ n167 ;
  assign n180 = n174 ^ n170 ;
  assign n181 = n179 & ~n180 ;
  assign n182 = n181 ^ n167 ;
  assign n183 = ~n177 & n182 ;
  assign n184 = n183 ^ n167 ;
  assign n185 = n184 ^ n13 ;
  assign n186 = n185 ^ n167 ;
  assign n187 = ~n161 & ~n186 ;
  assign n188 = x8 & ~n187 ;
  assign n189 = ~n160 & ~n188 ;
  assign n192 = x9 ^ x5 ;
  assign n190 = x9 ^ x4 ;
  assign n191 = n190 ^ x3 ;
  assign n193 = n192 ^ n191 ;
  assign n194 = n193 ^ n192 ;
  assign n195 = n194 ^ n190 ;
  assign n196 = n192 ^ n190 ;
  assign n197 = ~n194 & n196 ;
  assign n198 = n197 ^ n195 ;
  assign n199 = n114 & n198 ;
  assign n200 = n199 ^ n197 ;
  assign n201 = n195 & n200 ;
  assign n202 = n201 ^ n197 ;
  assign n203 = ~x7 & n202 ;
  assign n204 = n203 ^ x2 ;
  assign n205 = n20 & n23 ;
  assign n206 = n205 ^ n24 ;
  assign n207 = n204 & n206 ;
  assign n208 = n207 ^ n205 ;
  assign n209 = n24 & n208 ;
  assign n210 = n209 ^ x1 ;
  assign n211 = n189 & ~n210 ;
  assign n212 = x6 & ~n211 ;
  assign n213 = ~n158 & n212 ;
  assign n214 = ~n126 & ~n213 ;
  assign n215 = n214 ^ x0 ;
  assign n216 = n215 ^ n214 ;
  assign n217 = ~x6 & ~x7 ;
  assign n218 = ~x5 & n217 ;
  assign n219 = ~x2 & n218 ;
  assign n220 = x3 & ~n219 ;
  assign n221 = ~n115 & ~n220 ;
  assign n222 = ~n118 & ~n218 ;
  assign n223 = x1 & n15 ;
  assign n224 = ~n222 & n223 ;
  assign n225 = n221 & n224 ;
  assign n227 = x5 & x8 ;
  assign n226 = x6 & ~x8 ;
  assign n228 = n227 ^ n226 ;
  assign n229 = n228 ^ n227 ;
  assign n230 = n227 ^ x5 ;
  assign n231 = n230 ^ n227 ;
  assign n232 = n229 & ~n231 ;
  assign n233 = n232 ^ n227 ;
  assign n234 = ~x3 & n233 ;
  assign n235 = n234 ^ n227 ;
  assign n236 = n18 & n235 ;
  assign n237 = x5 & n139 ;
  assign n238 = ~x6 & n237 ;
  assign n239 = ~n236 & ~n238 ;
  assign n240 = ~x4 & ~n239 ;
  assign n241 = x3 & ~x6 ;
  assign n242 = n137 & n241 ;
  assign n243 = n242 ^ x4 ;
  assign n244 = n242 ^ x5 ;
  assign n245 = n244 ^ x5 ;
  assign n246 = n245 ^ n243 ;
  assign n247 = ~n29 & ~n163 ;
  assign n248 = ~x3 & x6 ;
  assign n249 = n138 & n248 ;
  assign n250 = n249 ^ n247 ;
  assign n251 = ~n247 & ~n250 ;
  assign n252 = n251 ^ x5 ;
  assign n253 = n252 ^ n247 ;
  assign n254 = ~n246 & ~n253 ;
  assign n255 = n254 ^ n251 ;
  assign n256 = n255 ^ n247 ;
  assign n257 = n243 & ~n256 ;
  assign n258 = n257 ^ n242 ;
  assign n259 = ~n240 & ~n258 ;
  assign n260 = n259 ^ x1 ;
  assign n261 = n260 ^ n259 ;
  assign n262 = n261 ^ x2 ;
  assign n263 = ~x6 & x8 ;
  assign n264 = n263 ^ x3 ;
  assign n265 = n264 ^ x9 ;
  assign n266 = n263 ^ n226 ;
  assign n267 = ~n226 & n266 ;
  assign n268 = n267 ^ n226 ;
  assign n269 = n264 ^ n226 ;
  assign n270 = ~n268 & n269 ;
  assign n271 = n270 ^ n267 ;
  assign n272 = n271 ^ n226 ;
  assign n273 = n272 ^ n263 ;
  assign n274 = n265 & n273 ;
  assign n275 = n274 ^ n264 ;
  assign n276 = n127 & n275 ;
  assign n277 = ~n217 & ~n248 ;
  assign n278 = n114 & ~n277 ;
  assign n279 = x5 & n278 ;
  assign n280 = ~n276 & ~n279 ;
  assign n281 = x4 & ~n280 ;
  assign n282 = n11 & n263 ;
  assign n283 = ~n122 & n282 ;
  assign n284 = ~n163 & n283 ;
  assign n285 = n284 ^ n281 ;
  assign n286 = ~n281 & n285 ;
  assign n287 = n286 ^ n259 ;
  assign n288 = n287 ^ n281 ;
  assign n289 = n262 & ~n288 ;
  assign n290 = n289 ^ n286 ;
  assign n291 = n290 ^ n281 ;
  assign n292 = x2 & ~n291 ;
  assign n293 = n292 ^ x2 ;
  assign n294 = ~n225 & ~n293 ;
  assign n295 = ~x3 & ~x5 ;
  assign n296 = n138 & n295 ;
  assign n297 = n296 ^ n159 ;
  assign n302 = n297 ^ n296 ;
  assign n298 = ~x3 & ~n230 ;
  assign n299 = n298 ^ x5 ;
  assign n300 = n299 ^ n297 ;
  assign n301 = n300 ^ n297 ;
  assign n303 = n302 ^ n301 ;
  assign n304 = ~x1 & ~x7 ;
  assign n305 = n304 ^ n297 ;
  assign n306 = n305 ^ n297 ;
  assign n307 = n306 ^ n301 ;
  assign n308 = ~n301 & ~n307 ;
  assign n309 = n308 ^ n301 ;
  assign n310 = n303 & ~n309 ;
  assign n311 = n310 ^ n308 ;
  assign n312 = n311 ^ n297 ;
  assign n313 = n312 ^ n301 ;
  assign n314 = x6 & ~n313 ;
  assign n315 = n314 ^ n296 ;
  assign n316 = ~x9 & n315 ;
  assign n317 = ~x3 & n263 ;
  assign n318 = n29 & n317 ;
  assign n319 = n304 & n318 ;
  assign n320 = ~n316 & ~n319 ;
  assign n321 = n320 ^ x4 ;
  assign n322 = n321 ^ n320 ;
  assign n337 = ~x7 & ~n114 ;
  assign n338 = x3 & ~n337 ;
  assign n339 = x9 ^ x8 ;
  assign n340 = x8 ^ x6 ;
  assign n341 = ~n339 & ~n340 ;
  assign n342 = n341 ^ x6 ;
  assign n343 = ~n338 & n342 ;
  assign n344 = x6 & n58 ;
  assign n345 = n344 ^ n21 ;
  assign n346 = n345 ^ n21 ;
  assign n347 = n217 ^ n21 ;
  assign n348 = n347 ^ n21 ;
  assign n349 = ~n346 & ~n348 ;
  assign n350 = n349 ^ n21 ;
  assign n351 = ~x5 & n350 ;
  assign n352 = n351 ^ n21 ;
  assign n353 = n343 & ~n352 ;
  assign n323 = x7 ^ x5 ;
  assign n324 = n323 ^ x9 ;
  assign n325 = n317 ^ x9 ;
  assign n326 = n325 ^ n324 ;
  assign n327 = x6 & ~n227 ;
  assign n328 = x3 & n327 ;
  assign n329 = n328 ^ x7 ;
  assign n330 = ~x9 & ~n329 ;
  assign n331 = n330 ^ x7 ;
  assign n332 = ~n326 & n331 ;
  assign n333 = n332 ^ n330 ;
  assign n334 = n333 ^ x7 ;
  assign n335 = n334 ^ x9 ;
  assign n336 = n324 & ~n335 ;
  assign n354 = n353 ^ n336 ;
  assign n355 = ~x1 & n354 ;
  assign n356 = n355 ^ n336 ;
  assign n357 = n356 ^ n320 ;
  assign n358 = ~n322 & ~n357 ;
  assign n359 = n358 ^ n320 ;
  assign n360 = ~x2 & ~n359 ;
  assign n361 = n294 & ~n360 ;
  assign n362 = n361 ^ n214 ;
  assign n363 = ~n216 & n362 ;
  assign n364 = n363 ^ n214 ;
  assign n365 = n364 ^ n113 ;
  assign n366 = n121 & ~n365 ;
  assign n367 = n366 ^ n363 ;
  assign n368 = n367 ^ n214 ;
  assign n369 = n368 ^ n120 ;
  assign n370 = ~n113 & ~n369 ;
  assign n371 = n370 ^ n113 ;
  assign y0 = n371 ;
endmodule
