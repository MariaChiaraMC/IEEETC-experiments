module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n11 = x6 & x8 ;
  assign n12 = x5 & ~n11 ;
  assign n13 = x9 & ~n12 ;
  assign n14 = ~x6 & ~x8 ;
  assign n15 = n14 ^ x7 ;
  assign n16 = x0 & x2 ;
  assign n17 = x1 & ~x4 ;
  assign n18 = ~x3 & ~n17 ;
  assign n19 = n16 & n18 ;
  assign n20 = n19 ^ n14 ;
  assign n21 = x7 ^ x5 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = ~n19 & n22 ;
  assign n24 = n23 ^ n19 ;
  assign n25 = ~n20 & ~n24 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n26 ^ n19 ;
  assign n28 = n27 ^ n21 ;
  assign n29 = n15 & n28 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = ~n13 & n30 ;
  assign y0 = n31 ;
endmodule
