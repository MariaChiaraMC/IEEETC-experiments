module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 ;
  assign n9 = ~x1 & x2 ;
  assign n10 = x3 & x4 ;
  assign n11 = n10 ^ x6 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = n10 ^ x3 ;
  assign n14 = ~n12 & ~n13 ;
  assign n15 = n14 ^ n10 ;
  assign n16 = n9 & n15 ;
  assign n17 = ~x6 & ~x7 ;
  assign n18 = x3 ^ x2 ;
  assign n19 = n18 ^ n9 ;
  assign n20 = ~n17 & n19 ;
  assign n21 = n20 ^ n17 ;
  assign n22 = x4 ^ x2 ;
  assign n23 = n22 ^ n20 ;
  assign n24 = ~n18 & n23 ;
  assign n25 = n24 ^ n18 ;
  assign n26 = n25 ^ n9 ;
  assign n27 = ~n21 & n26 ;
  assign n28 = ~n16 & ~n27 ;
  assign n29 = x5 & ~n28 ;
  assign n30 = ~x2 & ~x4 ;
  assign n31 = x6 & x7 ;
  assign n32 = x3 & ~n31 ;
  assign n33 = n30 & n32 ;
  assign n34 = ~x5 & n30 ;
  assign n35 = ~x0 & ~n34 ;
  assign n36 = x2 & ~x3 ;
  assign n37 = x5 ^ x4 ;
  assign n38 = n37 ^ x5 ;
  assign n39 = x6 ^ x5 ;
  assign n40 = ~n38 & ~n39 ;
  assign n41 = n40 ^ x5 ;
  assign n42 = n36 & ~n41 ;
  assign n43 = n35 & ~n42 ;
  assign n44 = ~n33 & n43 ;
  assign n45 = ~x1 & ~n44 ;
  assign n46 = ~n29 & ~n45 ;
  assign n52 = x2 & n10 ;
  assign n47 = x2 & ~n13 ;
  assign n48 = n47 ^ x3 ;
  assign n49 = x1 & ~n48 ;
  assign n50 = ~n31 & n34 ;
  assign n51 = ~n49 & ~n50 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = ~x0 & n53 ;
  assign n55 = n54 ^ n52 ;
  assign n56 = n46 & n55 ;
  assign y0 = ~n56 ;
endmodule
