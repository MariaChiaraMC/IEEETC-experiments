module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 ;
  assign n17 = x4 & ~x6 ;
  assign n18 = x4 & x5 ;
  assign n19 = ~x14 & n18 ;
  assign n20 = x8 ^ x5 ;
  assign n21 = x8 ^ x4 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = x6 ^ x4 ;
  assign n24 = n22 & ~n23 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = ~n20 & n25 ;
  assign n27 = n26 ^ x5 ;
  assign n28 = ~x11 & n27 ;
  assign n29 = ~n19 & ~n28 ;
  assign n30 = ~x10 & ~n29 ;
  assign n31 = ~n17 & ~n30 ;
  assign n32 = x10 & ~x11 ;
  assign n33 = ~x10 & x11 ;
  assign n34 = ~n32 & ~n33 ;
  assign n35 = n34 ^ x4 ;
  assign n36 = n35 ^ n34 ;
  assign n37 = n34 ^ x8 ;
  assign n38 = n37 ^ n34 ;
  assign n39 = ~n36 & ~n38 ;
  assign n40 = n39 ^ n34 ;
  assign n41 = x6 & ~n40 ;
  assign n42 = n41 ^ n34 ;
  assign n43 = n42 ^ x5 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = n44 ^ x7 ;
  assign n46 = x14 & ~x15 ;
  assign n47 = x12 & ~x13 ;
  assign n48 = ~n46 & n47 ;
  assign n49 = x11 ^ x10 ;
  assign n50 = ~x14 & ~n32 ;
  assign n51 = n50 ^ x11 ;
  assign n52 = n49 & ~n51 ;
  assign n53 = n52 ^ x11 ;
  assign n54 = n48 & ~n53 ;
  assign n55 = n54 ^ x4 ;
  assign n56 = ~n54 & ~n55 ;
  assign n57 = n56 ^ n42 ;
  assign n58 = n57 ^ n54 ;
  assign n59 = n45 & n58 ;
  assign n60 = n59 ^ n56 ;
  assign n61 = n60 ^ n54 ;
  assign n62 = x7 & ~n61 ;
  assign n63 = n62 ^ x7 ;
  assign n64 = n31 & n63 ;
  assign n65 = ~x4 & x6 ;
  assign n66 = ~n34 & n65 ;
  assign n67 = ~x4 & ~x5 ;
  assign n68 = x6 ^ x5 ;
  assign n69 = ~n34 & ~n50 ;
  assign n70 = n48 & n69 ;
  assign n71 = x13 ^ x12 ;
  assign n72 = n71 ^ x13 ;
  assign n73 = x14 & x15 ;
  assign n74 = n73 ^ x13 ;
  assign n75 = ~n72 & n74 ;
  assign n76 = n75 ^ x13 ;
  assign n77 = n33 & n76 ;
  assign n78 = ~n70 & ~n77 ;
  assign n79 = n32 & n46 ;
  assign n80 = n78 & ~n79 ;
  assign n81 = n80 ^ n18 ;
  assign n82 = n68 & n81 ;
  assign n83 = n82 ^ n80 ;
  assign n84 = n18 & n83 ;
  assign n85 = ~n67 & ~n84 ;
  assign n86 = ~x7 & ~n85 ;
  assign n87 = ~n66 & n86 ;
  assign n88 = ~x3 & x9 ;
  assign n89 = ~x0 & ~x1 ;
  assign n90 = ~x2 & n89 ;
  assign n91 = n88 & n90 ;
  assign n92 = ~n87 & n91 ;
  assign n93 = ~n64 & n92 ;
  assign y0 = n93 ;
endmodule
