module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 ;
  assign n14 = x0 & ~x2 ;
  assign n9 = ~x5 & ~x7 ;
  assign n10 = ~x4 & x6 ;
  assign n11 = n9 & n10 ;
  assign n12 = n11 ^ x3 ;
  assign n13 = n12 ^ x1 ;
  assign n15 = n14 ^ n13 ;
  assign n16 = n15 ^ n13 ;
  assign n17 = n13 ^ n12 ;
  assign n18 = n17 ^ x3 ;
  assign n19 = n16 & n18 ;
  assign n20 = n19 ^ n12 ;
  assign n21 = x5 & n12 ;
  assign n22 = n21 ^ x3 ;
  assign n23 = n20 & n22 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = x3 & n24 ;
  assign n26 = n25 ^ n19 ;
  assign n27 = n26 ^ n11 ;
  assign n28 = n27 ^ n12 ;
  assign y0 = ~n28 ;
endmodule
