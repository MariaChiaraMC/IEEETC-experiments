module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 ;
  assign n25 = x5 & x6 ;
  assign n26 = ~x4 & ~n25 ;
  assign n9 = x4 ^ x2 ;
  assign n10 = x6 & x7 ;
  assign n11 = n10 ^ x4 ;
  assign n12 = n11 ^ x4 ;
  assign n13 = n12 ^ n9 ;
  assign n15 = ~x5 & ~x7 ;
  assign n14 = ~x6 & ~x7 ;
  assign n16 = n15 ^ n14 ;
  assign n17 = x4 & n16 ;
  assign n18 = n17 ^ n14 ;
  assign n19 = ~n13 & ~n18 ;
  assign n20 = n19 ^ n17 ;
  assign n21 = n20 ^ n14 ;
  assign n22 = n21 ^ x4 ;
  assign n23 = n9 & ~n22 ;
  assign n24 = n23 ^ x2 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = n27 ^ x1 ;
  assign n38 = n28 ^ n27 ;
  assign n29 = ~x2 & ~x4 ;
  assign n30 = x5 & n10 ;
  assign n31 = n29 & ~n30 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = n32 ^ n27 ;
  assign n34 = n31 ^ n24 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = n35 ^ n33 ;
  assign n37 = n33 & ~n36 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = n39 ^ n33 ;
  assign n41 = n27 ^ x6 ;
  assign n42 = n37 ^ n33 ;
  assign n43 = n41 & n42 ;
  assign n44 = n43 ^ n27 ;
  assign n45 = n40 & n44 ;
  assign n46 = n45 ^ n27 ;
  assign n47 = n46 ^ n24 ;
  assign n48 = n47 ^ n27 ;
  assign n49 = ~x3 & ~n48 ;
  assign n52 = x4 & ~x5 ;
  assign n50 = ~x2 & ~x7 ;
  assign n51 = x3 & n50 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = n51 ^ n10 ;
  assign n55 = n54 ^ n10 ;
  assign n56 = n10 ^ x6 ;
  assign n57 = n55 & ~n56 ;
  assign n58 = n57 ^ n10 ;
  assign n59 = n53 & ~n58 ;
  assign n60 = n59 ^ n52 ;
  assign n61 = ~x1 & n60 ;
  assign n62 = ~x1 & ~x6 ;
  assign n63 = x5 ^ x4 ;
  assign n64 = n63 ^ x7 ;
  assign n65 = x7 ^ x5 ;
  assign n66 = n65 ^ x7 ;
  assign n67 = n66 ^ n64 ;
  assign n68 = x3 ^ x2 ;
  assign n69 = x7 & n68 ;
  assign n70 = n69 ^ x2 ;
  assign n71 = n67 & ~n70 ;
  assign n72 = n71 ^ n69 ;
  assign n73 = n72 ^ x2 ;
  assign n74 = n73 ^ x7 ;
  assign n75 = n64 & ~n74 ;
  assign n76 = n62 & n75 ;
  assign n77 = x4 & x5 ;
  assign n78 = n77 ^ x2 ;
  assign n79 = x1 & n10 ;
  assign n80 = n79 ^ n78 ;
  assign n81 = n80 ^ n77 ;
  assign n82 = n81 ^ n80 ;
  assign n83 = x6 & n15 ;
  assign n84 = x4 & ~x7 ;
  assign n85 = x3 & ~x5 ;
  assign n86 = ~n84 & n85 ;
  assign n87 = ~n83 & ~n86 ;
  assign n88 = ~x1 & n87 ;
  assign n89 = n88 ^ n80 ;
  assign n90 = n89 ^ n78 ;
  assign n91 = n82 & n90 ;
  assign n92 = n91 ^ n88 ;
  assign n93 = ~n14 & n88 ;
  assign n94 = n93 ^ n78 ;
  assign n95 = n92 & ~n94 ;
  assign n96 = n95 ^ n93 ;
  assign n97 = ~n78 & n96 ;
  assign n98 = n97 ^ n91 ;
  assign n99 = n98 ^ x2 ;
  assign n100 = n99 ^ n88 ;
  assign n101 = ~n76 & ~n100 ;
  assign n102 = ~n61 & n101 ;
  assign n103 = ~n49 & n102 ;
  assign n104 = ~x0 & ~n103 ;
  assign y0 = n104 ;
endmodule
