module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 ;
  assign n10 = x7 & x8 ;
  assign n16 = ~x2 & ~x5 ;
  assign n66 = n10 & n16 ;
  assign n67 = x6 & x7 ;
  assign n80 = n16 & n67 ;
  assign n35 = ~x7 & ~x8 ;
  assign n72 = x2 & ~x6 ;
  assign n81 = n35 & n72 ;
  assign n82 = x5 & n81 ;
  assign n83 = ~n80 & ~n82 ;
  assign n22 = ~x2 & ~x8 ;
  assign n68 = ~n22 & n67 ;
  assign n69 = n68 ^ x5 ;
  assign n70 = n68 ^ x8 ;
  assign n71 = n70 ^ x8 ;
  assign n73 = ~x7 & x8 ;
  assign n74 = n72 & n73 ;
  assign n75 = n74 ^ x8 ;
  assign n76 = ~n71 & n75 ;
  assign n77 = n76 ^ x8 ;
  assign n78 = ~n69 & ~n77 ;
  assign n79 = n78 ^ x5 ;
  assign n84 = n83 ^ n79 ;
  assign n85 = x1 & n84 ;
  assign n86 = n85 ^ n79 ;
  assign n87 = ~n66 & n86 ;
  assign n11 = x1 & x2 ;
  assign n12 = n10 & n11 ;
  assign n13 = x5 & n10 ;
  assign n14 = ~x4 & n13 ;
  assign n15 = ~x2 & n14 ;
  assign n17 = ~x4 & ~n16 ;
  assign n18 = x1 & x7 ;
  assign n19 = ~x8 & n18 ;
  assign n20 = ~n17 & n19 ;
  assign n21 = x5 & ~x7 ;
  assign n23 = ~x4 & n22 ;
  assign n24 = x4 & x8 ;
  assign n25 = ~n23 & ~n24 ;
  assign n26 = n21 & ~n25 ;
  assign n27 = ~n20 & ~n26 ;
  assign n28 = ~n15 & n27 ;
  assign n29 = n28 ^ x6 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = x2 & n13 ;
  assign n32 = x5 & n18 ;
  assign n33 = n23 & n32 ;
  assign n34 = ~n31 & ~n33 ;
  assign n37 = ~x5 & x8 ;
  assign n38 = x1 & n37 ;
  assign n36 = ~x5 & n35 ;
  assign n39 = n38 ^ n36 ;
  assign n40 = n39 ^ x4 ;
  assign n48 = n40 ^ n39 ;
  assign n41 = x5 & ~n11 ;
  assign n42 = n41 ^ n40 ;
  assign n43 = n42 ^ n39 ;
  assign n44 = n40 ^ n36 ;
  assign n45 = n44 ^ n41 ;
  assign n46 = n45 ^ n43 ;
  assign n47 = ~n43 & n46 ;
  assign n49 = n48 ^ n47 ;
  assign n50 = n49 ^ n43 ;
  assign n51 = ~x1 & ~x2 ;
  assign n52 = ~x7 & ~n51 ;
  assign n53 = n52 ^ n39 ;
  assign n54 = n47 ^ n43 ;
  assign n55 = n53 & ~n54 ;
  assign n56 = n55 ^ n39 ;
  assign n57 = ~n50 & n56 ;
  assign n58 = n57 ^ n39 ;
  assign n59 = n58 ^ n38 ;
  assign n60 = n59 ^ n39 ;
  assign n61 = n34 & ~n60 ;
  assign n62 = n61 ^ n28 ;
  assign n63 = n30 & n62 ;
  assign n64 = n63 ^ n28 ;
  assign n65 = ~n12 & n64 ;
  assign n88 = n87 ^ n65 ;
  assign n89 = n88 ^ n87 ;
  assign n90 = ~x5 & ~x6 ;
  assign n91 = x8 & n90 ;
  assign n92 = ~x2 & n91 ;
  assign n93 = ~n80 & ~n92 ;
  assign n94 = ~n81 & n93 ;
  assign n95 = ~x4 & ~n94 ;
  assign n97 = x4 & x6 ;
  assign n98 = ~n24 & ~n97 ;
  assign n99 = x2 & ~n98 ;
  assign n96 = ~n10 & n72 ;
  assign n100 = n99 ^ n96 ;
  assign n101 = n100 ^ x5 ;
  assign n108 = n101 ^ n100 ;
  assign n102 = n101 ^ n35 ;
  assign n103 = n102 ^ n100 ;
  assign n104 = n101 ^ n96 ;
  assign n105 = n104 ^ n35 ;
  assign n106 = n105 ^ n103 ;
  assign n107 = ~n103 & ~n106 ;
  assign n109 = n108 ^ n107 ;
  assign n110 = n109 ^ n103 ;
  assign n111 = n100 ^ x6 ;
  assign n112 = n107 ^ n103 ;
  assign n113 = n111 & ~n112 ;
  assign n114 = n113 ^ n100 ;
  assign n115 = ~n110 & n114 ;
  assign n116 = n115 ^ n100 ;
  assign n117 = n116 ^ n99 ;
  assign n118 = n117 ^ n100 ;
  assign n119 = ~n95 & ~n118 ;
  assign n120 = ~x1 & ~n119 ;
  assign n121 = n120 ^ n87 ;
  assign n122 = n121 ^ n87 ;
  assign n123 = n89 & ~n122 ;
  assign n124 = n123 ^ n87 ;
  assign n125 = ~x3 & n124 ;
  assign n126 = n125 ^ n87 ;
  assign n127 = x3 & x5 ;
  assign n128 = n72 & n127 ;
  assign n129 = n10 & n128 ;
  assign n130 = x7 & ~x8 ;
  assign n131 = x1 & ~x2 ;
  assign n132 = n130 & n131 ;
  assign n133 = x3 & ~x6 ;
  assign n134 = ~x1 & ~x7 ;
  assign n135 = n133 & n134 ;
  assign n136 = x6 & ~x8 ;
  assign n137 = n136 ^ x3 ;
  assign n138 = n137 ^ n136 ;
  assign n139 = n136 ^ n73 ;
  assign n140 = n139 ^ n136 ;
  assign n141 = n138 & n140 ;
  assign n142 = n141 ^ n136 ;
  assign n143 = x1 & n142 ;
  assign n144 = n143 ^ n136 ;
  assign n145 = x2 & n144 ;
  assign n146 = ~n135 & ~n145 ;
  assign n147 = ~n132 & n146 ;
  assign n148 = ~x5 & ~n147 ;
  assign n149 = x3 ^ x2 ;
  assign n150 = x5 & x8 ;
  assign n151 = n150 ^ x3 ;
  assign n152 = n151 ^ n150 ;
  assign n153 = n152 ^ n149 ;
  assign n154 = n35 ^ x5 ;
  assign n155 = x5 & n154 ;
  assign n156 = n155 ^ n150 ;
  assign n157 = n156 ^ x5 ;
  assign n158 = ~n153 & ~n157 ;
  assign n159 = n158 ^ n155 ;
  assign n160 = n159 ^ x5 ;
  assign n161 = ~n149 & n160 ;
  assign n162 = n161 ^ x2 ;
  assign n163 = x6 & ~n162 ;
  assign n164 = x5 & ~x8 ;
  assign n165 = ~n67 & ~n164 ;
  assign n166 = x2 & ~n165 ;
  assign n167 = ~n136 & n166 ;
  assign n168 = ~n13 & ~n167 ;
  assign n169 = ~n163 & n168 ;
  assign n170 = x1 & ~n169 ;
  assign n171 = ~n148 & ~n170 ;
  assign n172 = ~n129 & n171 ;
  assign n173 = n172 ^ x4 ;
  assign n174 = n173 ^ n172 ;
  assign n175 = n51 & n150 ;
  assign n176 = ~x7 & n175 ;
  assign n177 = ~x5 & ~n10 ;
  assign n178 = ~n134 & n177 ;
  assign n179 = n178 ^ x2 ;
  assign n180 = n179 ^ x3 ;
  assign n181 = n180 ^ n178 ;
  assign n187 = n181 ^ n179 ;
  assign n188 = n187 ^ n178 ;
  assign n189 = n188 ^ n178 ;
  assign n190 = ~x1 & x5 ;
  assign n191 = x2 & ~n130 ;
  assign n192 = ~n190 & n191 ;
  assign n193 = n192 ^ n179 ;
  assign n194 = n193 ^ n179 ;
  assign n195 = n194 ^ n178 ;
  assign n196 = n189 & ~n195 ;
  assign n182 = ~n10 & ~n21 ;
  assign n183 = n182 ^ n179 ;
  assign n184 = n183 ^ n181 ;
  assign n185 = n184 ^ n178 ;
  assign n186 = n181 & ~n185 ;
  assign n197 = n196 ^ n186 ;
  assign n198 = n197 ^ n181 ;
  assign n199 = n186 ^ n178 ;
  assign n200 = n199 ^ n188 ;
  assign n201 = n178 & n200 ;
  assign n202 = n201 ^ n186 ;
  assign n203 = n198 & n202 ;
  assign n204 = n203 ^ n196 ;
  assign n205 = n204 ^ n201 ;
  assign n206 = n205 ^ n181 ;
  assign n207 = n206 ^ n178 ;
  assign n208 = n207 ^ n188 ;
  assign n209 = n208 ^ x2 ;
  assign n210 = ~n176 & ~n209 ;
  assign n211 = n210 ^ x3 ;
  assign n212 = n211 ^ n210 ;
  assign n216 = x5 ^ x2 ;
  assign n217 = n216 ^ x7 ;
  assign n218 = n217 ^ x8 ;
  assign n213 = x2 ^ x1 ;
  assign n214 = n213 ^ x8 ;
  assign n227 = n218 ^ n214 ;
  assign n215 = n214 ^ x7 ;
  assign n219 = n218 ^ n215 ;
  assign n220 = n219 ^ n218 ;
  assign n221 = n220 ^ n214 ;
  assign n222 = n218 ^ x5 ;
  assign n223 = n222 ^ x8 ;
  assign n224 = n223 ^ n219 ;
  assign n225 = n224 ^ n221 ;
  assign n226 = ~n221 & ~n225 ;
  assign n228 = n227 ^ n226 ;
  assign n229 = n228 ^ n221 ;
  assign n230 = n214 ^ x8 ;
  assign n231 = n230 ^ n214 ;
  assign n232 = n226 ^ n221 ;
  assign n233 = ~n231 & ~n232 ;
  assign n234 = n233 ^ n214 ;
  assign n235 = n229 & n234 ;
  assign n236 = n235 ^ n214 ;
  assign n237 = n236 ^ x2 ;
  assign n238 = n237 ^ n214 ;
  assign n239 = n238 ^ n210 ;
  assign n240 = n239 ^ n210 ;
  assign n241 = n212 & ~n240 ;
  assign n242 = n241 ^ n210 ;
  assign n243 = ~x6 & ~n242 ;
  assign n244 = n243 ^ n210 ;
  assign n245 = n244 ^ n172 ;
  assign n246 = ~n174 & n245 ;
  assign n247 = n246 ^ n172 ;
  assign n248 = n126 & n247 ;
  assign n249 = ~x0 & ~n248 ;
  assign n250 = n97 ^ x0 ;
  assign n251 = n250 ^ n37 ;
  assign n252 = n251 ^ n97 ;
  assign n253 = n252 ^ n251 ;
  assign n261 = n67 ^ x8 ;
  assign n262 = n261 ^ n67 ;
  assign n263 = n262 ^ x4 ;
  assign n254 = x8 ^ x7 ;
  assign n255 = n254 ^ x5 ;
  assign n264 = n255 ^ n67 ;
  assign n265 = n264 ^ x4 ;
  assign n266 = n265 ^ x4 ;
  assign n267 = n263 & ~n266 ;
  assign n256 = n67 ^ x5 ;
  assign n257 = n256 ^ n67 ;
  assign n258 = n257 ^ n255 ;
  assign n259 = n258 ^ x4 ;
  assign n260 = n255 & n259 ;
  assign n268 = n267 ^ n260 ;
  assign n269 = n268 ^ n255 ;
  assign n270 = n260 ^ x4 ;
  assign n271 = n270 ^ n265 ;
  assign n272 = x4 & ~n271 ;
  assign n273 = n272 ^ n260 ;
  assign n274 = n269 & n273 ;
  assign n275 = n274 ^ n267 ;
  assign n276 = n275 ^ n272 ;
  assign n277 = n276 ^ n255 ;
  assign n278 = n277 ^ x4 ;
  assign n279 = n278 ^ n265 ;
  assign n280 = n279 ^ n251 ;
  assign n281 = n280 ^ n250 ;
  assign n282 = n253 & n281 ;
  assign n283 = n282 ^ n279 ;
  assign n284 = ~n130 & n279 ;
  assign n285 = n284 ^ n250 ;
  assign n286 = n283 & ~n285 ;
  assign n287 = n286 ^ n284 ;
  assign n288 = ~n250 & n287 ;
  assign n289 = n288 ^ n282 ;
  assign n290 = n289 ^ x0 ;
  assign n291 = n290 ^ n279 ;
  assign n292 = n51 & n291 ;
  assign n293 = ~x3 & n292 ;
  assign n294 = ~n249 & ~n293 ;
  assign y0 = ~n294 ;
endmodule
