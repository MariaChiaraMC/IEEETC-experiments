module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n11 = ~x3 & ~x6 ;
  assign n12 = ~x4 & n11 ;
  assign n13 = ~x2 & x3 ;
  assign n14 = ~x5 & n13 ;
  assign n15 = ~n12 & ~n14 ;
  assign n16 = ~x0 & ~n15 ;
  assign n17 = x8 & ~n16 ;
  assign n18 = x2 & x5 ;
  assign n19 = n18 ^ x1 ;
  assign n20 = n19 ^ n18 ;
  assign n21 = x6 ^ x3 ;
  assign n22 = x7 ^ x6 ;
  assign n23 = n22 ^ x7 ;
  assign n24 = ~x4 & x5 ;
  assign n25 = n24 ^ x7 ;
  assign n26 = n23 & n25 ;
  assign n27 = n26 ^ x7 ;
  assign n28 = ~n21 & n27 ;
  assign n29 = n28 ^ n18 ;
  assign n30 = n20 & n29 ;
  assign n31 = n30 ^ n18 ;
  assign n32 = n17 & ~n31 ;
  assign y0 = ~n32 ;
endmodule
