module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 ;
  assign n17 = ~x9 & ~x10 ;
  assign n18 = x4 & x5 ;
  assign n19 = ~x6 & n18 ;
  assign n20 = x15 ^ x14 ;
  assign n21 = ~x13 & ~n20 ;
  assign n22 = n19 & ~n21 ;
  assign n23 = ~n17 & n22 ;
  assign n24 = ~x8 & ~n23 ;
  assign n25 = ~x3 & ~x7 ;
  assign n26 = ~x0 & ~x2 ;
  assign n27 = x1 & ~x12 ;
  assign n28 = n26 & n27 ;
  assign n29 = ~x11 & n28 ;
  assign n30 = n25 & n29 ;
  assign n31 = x13 ^ x8 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = ~x4 & ~x5 ;
  assign n34 = ~x14 & ~x15 ;
  assign n35 = n17 & n34 ;
  assign n36 = n33 & n35 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = ~x13 & ~n37 ;
  assign n39 = n38 ^ n34 ;
  assign n40 = n32 & n39 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n41 ^ n34 ;
  assign n43 = n42 ^ x13 ;
  assign n44 = n30 & ~n43 ;
  assign n45 = ~n24 & n44 ;
  assign y0 = n45 ;
endmodule
