module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 ;
  assign n17 = ~x0 & ~x2 ;
  assign n18 = ~x3 & n17 ;
  assign n19 = x10 & n18 ;
  assign n20 = ~x1 & n19 ;
  assign n23 = x11 ^ x6 ;
  assign n21 = x9 ^ x5 ;
  assign n22 = n21 ^ x8 ;
  assign n24 = n23 ^ n22 ;
  assign n25 = n23 ^ x11 ;
  assign n26 = n25 ^ x5 ;
  assign n27 = n24 & n26 ;
  assign n28 = n27 ^ x11 ;
  assign n29 = ~x8 & ~x11 ;
  assign n30 = n29 ^ x5 ;
  assign n31 = ~n28 & n30 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = x5 & n32 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = n34 ^ x11 ;
  assign n36 = n35 ^ x5 ;
  assign n37 = n36 ^ n35 ;
  assign n38 = x6 & ~x11 ;
  assign n39 = n38 ^ n35 ;
  assign n40 = n39 ^ n35 ;
  assign n41 = ~n37 & ~n40 ;
  assign n42 = n41 ^ n35 ;
  assign n43 = ~x7 & n42 ;
  assign n44 = n43 ^ n35 ;
  assign n45 = n44 ^ x4 ;
  assign n46 = n45 ^ n44 ;
  assign n47 = n46 ^ n20 ;
  assign n48 = ~x5 & x6 ;
  assign n49 = x14 & ~x15 ;
  assign n50 = x12 & ~x13 ;
  assign n51 = ~n49 & ~n50 ;
  assign n52 = n38 & ~n51 ;
  assign n53 = ~x7 & ~n52 ;
  assign n54 = ~n48 & ~n53 ;
  assign n55 = ~x5 & ~x7 ;
  assign n56 = n55 ^ n54 ;
  assign n57 = ~n54 & n56 ;
  assign n58 = n57 ^ n44 ;
  assign n59 = n58 ^ n54 ;
  assign n60 = n47 & ~n59 ;
  assign n61 = n60 ^ n57 ;
  assign n62 = n61 ^ n54 ;
  assign n63 = n20 & ~n62 ;
  assign n64 = n63 ^ n20 ;
  assign y0 = n64 ;
endmodule
