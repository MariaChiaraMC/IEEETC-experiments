module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 ;
  assign n11 = x7 & x8 ;
  assign n12 = ~x7 & ~x8 ;
  assign n13 = ~n11 & ~n12 ;
  assign n14 = x3 & x9 ;
  assign n15 = ~x1 & ~x2 ;
  assign n16 = ~x4 & x6 ;
  assign n17 = n15 & n16 ;
  assign n18 = n14 & n17 ;
  assign n19 = ~n13 & n18 ;
  assign n20 = ~x0 & ~n19 ;
  assign n79 = ~x3 & ~x6 ;
  assign n120 = x8 ^ x1 ;
  assign n65 = ~x2 & ~x7 ;
  assign n80 = ~x4 & ~x9 ;
  assign n81 = n65 & n80 ;
  assign n121 = ~x2 & ~x4 ;
  assign n122 = x7 & n121 ;
  assign n123 = n122 ^ x9 ;
  assign n124 = n123 ^ n122 ;
  assign n125 = x2 & x4 ;
  assign n126 = n125 ^ n122 ;
  assign n127 = ~n124 & n126 ;
  assign n128 = n127 ^ n122 ;
  assign n129 = x1 & n128 ;
  assign n130 = ~n81 & ~n129 ;
  assign n131 = n130 ^ n120 ;
  assign n132 = n131 ^ x8 ;
  assign n133 = n132 ^ n131 ;
  assign n134 = ~x8 & x9 ;
  assign n135 = n121 & n134 ;
  assign n136 = n135 ^ n131 ;
  assign n137 = n136 ^ n120 ;
  assign n138 = n133 & n137 ;
  assign n139 = n138 ^ n135 ;
  assign n33 = ~x2 & x4 ;
  assign n140 = x7 & ~x9 ;
  assign n141 = n33 & n140 ;
  assign n24 = x2 & ~x4 ;
  assign n71 = ~x7 & x9 ;
  assign n142 = n24 & n71 ;
  assign n143 = ~n141 & ~n142 ;
  assign n144 = ~n135 & n143 ;
  assign n145 = n144 ^ n120 ;
  assign n146 = ~n139 & n145 ;
  assign n147 = n146 ^ n144 ;
  assign n148 = n120 & n147 ;
  assign n149 = n148 ^ n138 ;
  assign n150 = n149 ^ x1 ;
  assign n151 = n150 ^ n135 ;
  assign n152 = n79 & n151 ;
  assign n48 = x3 & ~x9 ;
  assign n153 = ~n12 & ~n48 ;
  assign n154 = ~x1 & ~n153 ;
  assign n155 = ~x8 & ~x9 ;
  assign n156 = ~x1 & x2 ;
  assign n157 = ~n155 & ~n156 ;
  assign n158 = x4 & x7 ;
  assign n51 = ~x3 & x4 ;
  assign n159 = x6 & ~n51 ;
  assign n160 = ~n158 & n159 ;
  assign n161 = x8 ^ x4 ;
  assign n162 = n161 ^ x8 ;
  assign n50 = x8 & x9 ;
  assign n163 = x3 & ~x7 ;
  assign n164 = ~n50 & ~n163 ;
  assign n165 = n164 ^ x8 ;
  assign n166 = ~n162 & n165 ;
  assign n167 = n166 ^ x8 ;
  assign n168 = x2 & ~x3 ;
  assign n169 = ~x8 & n168 ;
  assign n170 = n169 ^ n160 ;
  assign n171 = ~n167 & n170 ;
  assign n172 = n171 ^ n169 ;
  assign n173 = n160 & n172 ;
  assign n174 = n173 ^ n160 ;
  assign n175 = ~n157 & n174 ;
  assign n176 = ~n154 & n175 ;
  assign n177 = x3 & ~x6 ;
  assign n178 = ~x9 & ~n15 ;
  assign n179 = x7 ^ x4 ;
  assign n180 = ~x9 & n179 ;
  assign n181 = ~n178 & ~n180 ;
  assign n182 = ~n24 & ~n33 ;
  assign n183 = n182 ^ x1 ;
  assign n184 = n183 ^ n182 ;
  assign n185 = n184 ^ x9 ;
  assign n186 = n158 ^ x2 ;
  assign n187 = x2 & n186 ;
  assign n188 = n187 ^ n182 ;
  assign n189 = n188 ^ x2 ;
  assign n190 = ~n185 & ~n189 ;
  assign n191 = n190 ^ n187 ;
  assign n192 = n191 ^ x2 ;
  assign n193 = x9 & n192 ;
  assign n194 = n193 ^ x9 ;
  assign n195 = n181 & ~n194 ;
  assign n196 = n195 ^ x8 ;
  assign n197 = n196 ^ n195 ;
  assign n198 = n197 ^ n177 ;
  assign n199 = x7 ^ x2 ;
  assign n200 = x1 & x4 ;
  assign n201 = n200 ^ x7 ;
  assign n202 = n199 & n201 ;
  assign n203 = n202 ^ x7 ;
  assign n204 = n178 & ~n203 ;
  assign n205 = n71 & n121 ;
  assign n206 = n205 ^ n204 ;
  assign n207 = ~n204 & n206 ;
  assign n208 = n207 ^ n195 ;
  assign n209 = n208 ^ n204 ;
  assign n210 = n198 & n209 ;
  assign n211 = n210 ^ n207 ;
  assign n212 = n211 ^ n204 ;
  assign n213 = n177 & ~n212 ;
  assign n214 = n213 ^ n177 ;
  assign n215 = ~n176 & ~n214 ;
  assign n216 = ~n152 & n215 ;
  assign n64 = x4 & x6 ;
  assign n66 = n50 & n65 ;
  assign n67 = x3 & n66 ;
  assign n68 = ~n64 & n67 ;
  assign n49 = ~x4 & n48 ;
  assign n69 = n49 ^ x3 ;
  assign n70 = n69 ^ n49 ;
  assign n72 = n71 ^ n49 ;
  assign n73 = n72 ^ n49 ;
  assign n74 = ~n70 & n73 ;
  assign n75 = n74 ^ n49 ;
  assign n76 = x6 & n75 ;
  assign n77 = n76 ^ n49 ;
  assign n78 = x2 & n77 ;
  assign n82 = n79 & n81 ;
  assign n83 = x2 & x7 ;
  assign n84 = n14 & n64 ;
  assign n85 = ~n49 & ~n84 ;
  assign n86 = n83 & ~n85 ;
  assign n87 = ~n82 & ~n86 ;
  assign n88 = ~n78 & n87 ;
  assign n89 = ~x8 & ~n88 ;
  assign n97 = x9 ^ x2 ;
  assign n90 = x9 ^ x4 ;
  assign n91 = n90 ^ x3 ;
  assign n98 = n97 ^ n91 ;
  assign n92 = x9 ^ x6 ;
  assign n93 = n92 ^ n91 ;
  assign n94 = n93 ^ n90 ;
  assign n95 = n94 ^ x9 ;
  assign n96 = n95 ^ n91 ;
  assign n99 = n98 ^ n96 ;
  assign n102 = n95 ^ x9 ;
  assign n100 = n90 ^ x9 ;
  assign n101 = n100 ^ n96 ;
  assign n103 = n102 ^ n101 ;
  assign n104 = n99 & n103 ;
  assign n105 = n104 ^ n95 ;
  assign n106 = n105 ^ n100 ;
  assign n107 = n106 ^ n102 ;
  assign n108 = n101 ^ n98 ;
  assign n109 = ~n105 & n108 ;
  assign n110 = n109 ^ n95 ;
  assign n111 = n110 ^ n96 ;
  assign n112 = n111 ^ n98 ;
  assign n113 = ~n107 & ~n112 ;
  assign n114 = n11 & n113 ;
  assign n115 = ~n89 & ~n114 ;
  assign n116 = ~n68 & n115 ;
  assign n21 = x7 & ~x8 ;
  assign n22 = ~x3 & n21 ;
  assign n23 = x4 & ~x6 ;
  assign n25 = x6 & n24 ;
  assign n26 = ~n23 & ~n25 ;
  assign n27 = n26 ^ x9 ;
  assign n28 = n26 & ~n27 ;
  assign n29 = ~x2 & n28 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n22 & ~n30 ;
  assign n32 = ~x6 & ~x9 ;
  assign n34 = n32 & n33 ;
  assign n35 = n13 & n34 ;
  assign n36 = ~n31 & ~n35 ;
  assign n37 = ~x2 & x7 ;
  assign n38 = ~x6 & x8 ;
  assign n39 = n38 ^ x4 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = x6 & ~x8 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = n40 & n42 ;
  assign n44 = n43 ^ n38 ;
  assign n45 = n37 & n44 ;
  assign n46 = n14 & n45 ;
  assign n47 = x6 & ~x7 ;
  assign n52 = n50 & n51 ;
  assign n53 = ~n49 & ~n52 ;
  assign n54 = n47 & ~n53 ;
  assign n55 = x4 & ~n32 ;
  assign n56 = ~x4 & ~x6 ;
  assign n57 = n11 & ~n56 ;
  assign n58 = ~n55 & n57 ;
  assign n59 = x3 & n58 ;
  assign n60 = ~n54 & ~n59 ;
  assign n61 = x2 & ~n60 ;
  assign n62 = ~n46 & ~n61 ;
  assign n63 = n36 & n62 ;
  assign n117 = n116 ^ n63 ;
  assign n118 = x1 & n117 ;
  assign n119 = n118 ^ n116 ;
  assign n217 = n216 ^ n119 ;
  assign n218 = n217 ^ n216 ;
  assign n219 = ~x3 & n155 ;
  assign n220 = n23 & n219 ;
  assign n221 = n37 & n220 ;
  assign n222 = n221 ^ n216 ;
  assign n223 = n222 ^ n216 ;
  assign n224 = n218 & ~n223 ;
  assign n225 = n224 ^ n216 ;
  assign n226 = x5 & n225 ;
  assign n227 = n226 ^ n216 ;
  assign n228 = n20 & n227 ;
  assign n259 = x5 & x6 ;
  assign n260 = n122 & n259 ;
  assign n261 = x5 & ~x7 ;
  assign n262 = ~x4 & ~x7 ;
  assign n263 = x4 & n259 ;
  assign n264 = ~n262 & ~n263 ;
  assign n265 = x2 & ~n264 ;
  assign n266 = ~n261 & n265 ;
  assign n267 = ~n260 & ~n266 ;
  assign n268 = n134 & ~n267 ;
  assign n229 = x8 & ~x9 ;
  assign n230 = x4 & n229 ;
  assign n231 = n56 & n134 ;
  assign n232 = ~n230 & ~n231 ;
  assign n233 = n65 & ~n232 ;
  assign n235 = x9 & n64 ;
  assign n234 = ~x4 & ~n38 ;
  assign n236 = n235 ^ n234 ;
  assign n237 = n234 ^ n32 ;
  assign n238 = n234 ^ x8 ;
  assign n239 = n234 & ~n238 ;
  assign n240 = n239 ^ n234 ;
  assign n241 = n237 & n240 ;
  assign n242 = n241 ^ n239 ;
  assign n243 = n242 ^ n234 ;
  assign n244 = n243 ^ x8 ;
  assign n245 = n236 & ~n244 ;
  assign n246 = n245 ^ n234 ;
  assign n247 = n83 & n246 ;
  assign n248 = ~n233 & ~n247 ;
  assign n249 = n248 ^ x9 ;
  assign n250 = n249 ^ n248 ;
  assign n251 = x8 & n25 ;
  assign n252 = ~n45 & ~n251 ;
  assign n253 = n252 ^ n248 ;
  assign n254 = n253 ^ n248 ;
  assign n255 = ~n250 & ~n254 ;
  assign n256 = n255 ^ n248 ;
  assign n257 = x5 & ~n256 ;
  assign n258 = n257 ^ n248 ;
  assign n269 = n268 ^ n258 ;
  assign n270 = n269 ^ n258 ;
  assign n271 = ~x5 & n56 ;
  assign n272 = ~n263 & ~n271 ;
  assign n273 = n37 & n50 ;
  assign n274 = ~n272 & n273 ;
  assign n275 = n33 & n38 ;
  assign n276 = n140 ^ x7 ;
  assign n277 = ~x5 & ~n276 ;
  assign n278 = n277 ^ x7 ;
  assign n279 = n275 & ~n278 ;
  assign n280 = ~n274 & ~n279 ;
  assign n281 = n280 ^ n258 ;
  assign n282 = n281 ^ n258 ;
  assign n283 = ~n270 & n282 ;
  assign n284 = n283 ^ n258 ;
  assign n285 = x1 & n284 ;
  assign n286 = n285 ^ n258 ;
  assign n287 = n286 ^ x3 ;
  assign n288 = n287 ^ n286 ;
  assign n289 = n288 ^ x0 ;
  assign n290 = ~x1 & n21 ;
  assign n291 = n125 & n290 ;
  assign n292 = n259 & ~n291 ;
  assign n293 = x2 ^ x1 ;
  assign n294 = n293 ^ x4 ;
  assign n295 = n294 ^ x8 ;
  assign n296 = x4 ^ x2 ;
  assign n297 = n296 ^ x6 ;
  assign n298 = n297 ^ x4 ;
  assign n299 = n298 ^ x8 ;
  assign n300 = n299 ^ n297 ;
  assign n301 = n300 ^ n295 ;
  assign n302 = n297 ^ x6 ;
  assign n303 = n302 ^ x8 ;
  assign n304 = x8 & n303 ;
  assign n305 = n304 ^ n297 ;
  assign n306 = n305 ^ x8 ;
  assign n307 = n301 & n306 ;
  assign n308 = n307 ^ n304 ;
  assign n309 = n308 ^ x8 ;
  assign n310 = n295 & n309 ;
  assign n311 = x9 & ~n310 ;
  assign n312 = ~x4 & x8 ;
  assign n313 = ~x9 & ~n312 ;
  assign n314 = ~n178 & ~n313 ;
  assign n315 = x8 ^ x2 ;
  assign n316 = n200 & ~n315 ;
  assign n317 = ~n314 & ~n316 ;
  assign n318 = x7 & ~n32 ;
  assign n319 = ~n317 & n318 ;
  assign n320 = ~n311 & n319 ;
  assign n321 = n121 ^ x4 ;
  assign n322 = ~n229 & n321 ;
  assign n323 = n322 ^ x4 ;
  assign n324 = n47 & n323 ;
  assign n325 = ~x1 & n324 ;
  assign n326 = ~x5 & ~n325 ;
  assign n327 = ~n320 & n326 ;
  assign n328 = ~n292 & ~n327 ;
  assign n329 = x8 ^ x7 ;
  assign n330 = x7 ^ x1 ;
  assign n331 = n329 & n330 ;
  assign n332 = n121 & n331 ;
  assign n333 = ~x9 & n332 ;
  assign n334 = n65 & n134 ;
  assign n335 = n200 & n334 ;
  assign n336 = ~x6 & ~n335 ;
  assign n338 = x1 & ~x7 ;
  assign n339 = n125 & n338 ;
  assign n337 = x9 ^ x8 ;
  assign n340 = n339 ^ n337 ;
  assign n351 = n340 ^ n339 ;
  assign n341 = x4 & n15 ;
  assign n342 = n341 ^ n339 ;
  assign n343 = n342 ^ n340 ;
  assign n344 = n343 ^ n340 ;
  assign n345 = n344 ^ n339 ;
  assign n346 = n343 ^ x9 ;
  assign n347 = n346 ^ x7 ;
  assign n348 = n347 ^ n343 ;
  assign n349 = n348 ^ n345 ;
  assign n350 = n345 & ~n349 ;
  assign n352 = n351 ^ n350 ;
  assign n353 = n352 ^ n345 ;
  assign n354 = n339 ^ x7 ;
  assign n355 = n350 ^ n345 ;
  assign n356 = ~n354 & n355 ;
  assign n357 = n356 ^ n339 ;
  assign n358 = ~n353 & ~n357 ;
  assign n359 = n358 ^ n339 ;
  assign n360 = n359 ^ n337 ;
  assign n361 = n360 ^ n339 ;
  assign n362 = n336 & n361 ;
  assign n363 = ~n333 & n362 ;
  assign n364 = x5 & n363 ;
  assign n365 = n364 ^ n328 ;
  assign n366 = n328 & ~n365 ;
  assign n367 = n366 ^ n286 ;
  assign n368 = n367 ^ n328 ;
  assign n369 = ~n289 & ~n368 ;
  assign n370 = n369 ^ n366 ;
  assign n371 = n370 ^ n328 ;
  assign n372 = x0 & n371 ;
  assign n373 = n372 ^ x0 ;
  assign n374 = ~n228 & ~n373 ;
  assign n375 = x5 & ~x9 ;
  assign n376 = n121 & n375 ;
  assign n377 = ~x3 & x6 ;
  assign n378 = n377 ^ x8 ;
  assign n379 = n378 ^ n377 ;
  assign n380 = n377 ^ n177 ;
  assign n381 = ~n379 & n380 ;
  assign n382 = n381 ^ n377 ;
  assign n383 = ~n329 & n382 ;
  assign n384 = n376 & n383 ;
  assign n385 = x1 & n384 ;
  assign n386 = ~n374 & ~n385 ;
  assign y0 = ~n386 ;
endmodule
