module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 ;
  assign n8 = ~x4 & ~x5 ;
  assign n9 = x1 & ~n8 ;
  assign n10 = x0 & x2 ;
  assign n11 = ~x1 & ~x4 ;
  assign n12 = ~n10 & ~n11 ;
  assign n13 = ~n9 & ~n12 ;
  assign n14 = ~x5 & ~x6 ;
  assign n15 = x0 & n14 ;
  assign n16 = ~x2 & ~n15 ;
  assign n17 = n13 & ~n16 ;
  assign n18 = ~x3 & ~n17 ;
  assign n19 = x2 ^ x0 ;
  assign n20 = x4 & ~n14 ;
  assign n21 = n20 ^ x0 ;
  assign n22 = n19 & ~n21 ;
  assign n23 = n22 ^ x0 ;
  assign n24 = x1 & ~n23 ;
  assign n25 = n18 & ~n24 ;
  assign n26 = x2 ^ x1 ;
  assign n27 = n26 ^ n11 ;
  assign n28 = n27 ^ x2 ;
  assign n29 = n28 ^ n27 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n26 ^ x6 ;
  assign n32 = n26 ^ x5 ;
  assign n33 = ~n31 & ~n32 ;
  assign n34 = n27 ^ n26 ;
  assign n35 = n29 & n34 ;
  assign n36 = n35 ^ n30 ;
  assign n37 = n33 & ~n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = ~n30 & n38 ;
  assign n40 = n39 ^ n35 ;
  assign n41 = n40 ^ n26 ;
  assign n42 = ~x0 & ~n41 ;
  assign n43 = ~x0 & n9 ;
  assign n44 = ~n11 & ~n43 ;
  assign n45 = ~x2 & n44 ;
  assign n46 = x3 & ~n45 ;
  assign n47 = ~n42 & n46 ;
  assign n48 = ~n25 & ~n47 ;
  assign y0 = n48 ;
endmodule
