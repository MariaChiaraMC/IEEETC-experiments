module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 ;
  assign n13 = x4 & x8 ;
  assign n14 = ~x9 & x10 ;
  assign n15 = x2 & x7 ;
  assign n16 = n14 & ~n15 ;
  assign n17 = ~n13 & n16 ;
  assign n18 = x6 & ~n17 ;
  assign n19 = x7 ^ x4 ;
  assign n20 = n19 ^ x7 ;
  assign n21 = x6 & x8 ;
  assign n22 = n21 ^ x7 ;
  assign n23 = ~n20 & n22 ;
  assign n24 = n23 ^ x7 ;
  assign n25 = ~x3 & ~x7 ;
  assign n26 = n25 ^ x0 ;
  assign n27 = ~n24 & ~n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = ~x0 & n28 ;
  assign n30 = n29 ^ x0 ;
  assign n31 = x11 ^ x6 ;
  assign n32 = n14 ^ x11 ;
  assign n33 = x11 ^ x5 ;
  assign n34 = n33 ^ n14 ;
  assign n35 = ~n14 & ~n34 ;
  assign n36 = n35 ^ n14 ;
  assign n37 = ~n32 & ~n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = n38 ^ n14 ;
  assign n40 = n39 ^ n33 ;
  assign n41 = n31 & ~n40 ;
  assign n42 = n41 ^ n33 ;
  assign n43 = ~n30 & n42 ;
  assign n44 = ~n18 & n43 ;
  assign y0 = n44 ;
endmodule
