module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 ;
  output y0 ;
  wire n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 ;
  assign n26 = ~x19 & ~x21 ;
  assign n27 = ~x14 & ~x24 ;
  assign n28 = ~x15 & ~x22 ;
  assign n29 = n27 & n28 ;
  assign n30 = ~x18 & ~x23 ;
  assign n31 = n29 & n30 ;
  assign n32 = n26 & n31 ;
  assign n33 = ~x13 & ~x16 ;
  assign n34 = ~x11 & ~x17 ;
  assign n35 = ~x20 & n34 ;
  assign n36 = ~x12 & n35 ;
  assign n37 = n33 & n36 ;
  assign n38 = n32 & n37 ;
  assign n39 = x9 & n38 ;
  assign n40 = x18 & x23 ;
  assign n41 = x14 & x24 ;
  assign n42 = x15 & x22 ;
  assign n43 = n41 & n42 ;
  assign n44 = x19 & x21 ;
  assign n45 = n43 & n44 ;
  assign n46 = n40 & n45 ;
  assign n47 = x11 & x17 ;
  assign n48 = x20 & n47 ;
  assign n49 = x13 & x16 ;
  assign n50 = n48 & n49 ;
  assign n51 = x12 & n50 ;
  assign n52 = n46 & n51 ;
  assign n53 = x6 & n52 ;
  assign n54 = ~n39 & ~n53 ;
  assign n55 = ~x4 & ~x5 ;
  assign n56 = ~n54 & n55 ;
  assign n57 = ~x2 & n56 ;
  assign n61 = x3 & n52 ;
  assign n62 = x8 & n38 ;
  assign n63 = ~n61 & ~n62 ;
  assign n58 = x10 & n38 ;
  assign n59 = x7 & n52 ;
  assign n60 = ~n58 & ~n59 ;
  assign n64 = n63 ^ n60 ;
  assign n65 = n64 ^ x0 ;
  assign n66 = n65 ^ x1 ;
  assign n67 = n66 ^ n64 ;
  assign n68 = n64 ^ n60 ;
  assign n69 = n67 ^ x2 ;
  assign n70 = n69 ^ n67 ;
  assign n71 = ~n68 & ~n70 ;
  assign n72 = n71 ^ n64 ;
  assign n73 = n64 ^ x1 ;
  assign n74 = n69 & n73 ;
  assign n75 = n74 ^ n67 ;
  assign n76 = n75 ^ n69 ;
  assign n77 = n72 & ~n76 ;
  assign n78 = ~n67 & n77 ;
  assign n79 = n78 ^ n71 ;
  assign n80 = n79 ^ n63 ;
  assign n81 = ~n57 & n80 ;
  assign y0 = ~n81 ;
endmodule
