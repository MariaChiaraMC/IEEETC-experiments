module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 ;
  assign n17 = x3 & ~x7 ;
  assign n18 = ~x0 & ~x6 ;
  assign n19 = x5 & n18 ;
  assign n20 = n17 & n19 ;
  assign n21 = x1 ^ x0 ;
  assign n22 = n21 ^ x0 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n23 ^ n21 ;
  assign n25 = n21 & n24 ;
  assign n26 = n25 ^ n21 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = n27 ^ x3 ;
  assign n29 = n24 ^ x3 ;
  assign n30 = x9 & x10 ;
  assign n31 = x6 & ~n30 ;
  assign n32 = x7 & ~n31 ;
  assign n33 = ~x9 & ~x10 ;
  assign n34 = ~x8 & ~x11 ;
  assign n35 = ~x12 & n34 ;
  assign n36 = ~n33 & n35 ;
  assign n37 = x14 ^ x13 ;
  assign n38 = n37 ^ x15 ;
  assign n39 = x14 & x15 ;
  assign n40 = n38 & n39 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n36 & n41 ;
  assign n43 = ~n32 & n42 ;
  assign n44 = n43 ^ x7 ;
  assign n45 = n44 ^ n21 ;
  assign n46 = n29 & n45 ;
  assign n47 = n46 ^ x7 ;
  assign n48 = n47 ^ n23 ;
  assign n49 = n21 ^ x5 ;
  assign n50 = n49 ^ x7 ;
  assign n51 = n49 & n50 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = n52 ^ n21 ;
  assign n54 = n53 ^ n23 ;
  assign n55 = n54 ^ x3 ;
  assign n56 = n48 & n55 ;
  assign n57 = n56 ^ n21 ;
  assign n58 = n28 & n57 ;
  assign n59 = n58 ^ n56 ;
  assign n60 = n59 ^ n21 ;
  assign n61 = ~n20 & ~n60 ;
  assign y0 = ~n61 ;
endmodule
