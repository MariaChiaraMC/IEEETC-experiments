module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 ;
  assign n11 = x7 & ~x9 ;
  assign n12 = n11 ^ x3 ;
  assign n13 = ~x8 & ~n12 ;
  assign n14 = n13 ^ x3 ;
  assign n15 = x2 & ~n14 ;
  assign n16 = ~x3 & x8 ;
  assign n17 = ~x3 & ~x5 ;
  assign n18 = ~x7 & ~n17 ;
  assign n19 = ~n16 & n18 ;
  assign n20 = x3 & x9 ;
  assign n21 = ~x4 & ~n20 ;
  assign n22 = ~x8 & ~n21 ;
  assign n23 = ~n19 & ~n22 ;
  assign n24 = ~n15 & n23 ;
  assign y0 = n24 ;
endmodule
