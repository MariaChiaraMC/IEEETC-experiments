module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 ;
  output y0 ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 ;
  assign n18 = ~x1 & x10 ;
  assign n19 = x0 & x12 ;
  assign n20 = x15 & n19 ;
  assign n21 = n18 & n20 ;
  assign n22 = ~x8 & ~x9 ;
  assign n23 = x13 & n22 ;
  assign n24 = x14 & x16 ;
  assign n25 = x11 & n24 ;
  assign n26 = n23 & n25 ;
  assign n27 = n26 ^ n21 ;
  assign n28 = x3 & x7 ;
  assign n29 = x2 & n28 ;
  assign n30 = ~x6 & n29 ;
  assign n31 = n30 ^ x4 ;
  assign n32 = n31 ^ n30 ;
  assign n33 = x5 & ~x7 ;
  assign n34 = ~x3 & x6 ;
  assign n35 = n33 & n34 ;
  assign n36 = ~x2 & n35 ;
  assign n37 = n36 ^ n30 ;
  assign n38 = ~n32 & n37 ;
  assign n39 = n38 ^ n30 ;
  assign n40 = n39 ^ n21 ;
  assign n41 = n27 & n40 ;
  assign n42 = n41 ^ n38 ;
  assign n43 = n42 ^ n30 ;
  assign n44 = n43 ^ n26 ;
  assign n45 = n21 & n44 ;
  assign n46 = n45 ^ n21 ;
  assign y0 = n46 ;
endmodule
