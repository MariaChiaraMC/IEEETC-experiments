module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n13 = ~x8 & ~x10 ;
  assign n14 = ~x4 & ~n13 ;
  assign n15 = ~x5 & x7 ;
  assign n16 = ~x11 & ~n15 ;
  assign n17 = ~n14 & n16 ;
  assign n18 = ~x0 & ~x9 ;
  assign n19 = ~x6 & n18 ;
  assign n20 = x5 ^ x4 ;
  assign n21 = n20 ^ x5 ;
  assign n22 = x10 ^ x5 ;
  assign n23 = n21 & ~n22 ;
  assign n24 = n23 ^ x5 ;
  assign n25 = x5 & ~x7 ;
  assign n26 = n25 ^ n19 ;
  assign n27 = n24 & n26 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n19 & n28 ;
  assign n30 = n29 ^ n19 ;
  assign n31 = n17 & n30 ;
  assign y0 = n31 ;
endmodule
