module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 ;
  assign n15 = x12 & x13 ;
  assign n16 = ~x6 & ~x11 ;
  assign n17 = x3 & ~x5 ;
  assign n18 = x1 & ~x7 ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = n16 & ~n19 ;
  assign n21 = x7 & ~x10 ;
  assign n22 = x1 & x6 ;
  assign n23 = n21 & n22 ;
  assign n24 = x3 & ~x10 ;
  assign n25 = x5 & x6 ;
  assign n26 = n24 & n25 ;
  assign n27 = ~n23 & ~n26 ;
  assign n28 = ~n20 & n27 ;
  assign n29 = n15 & ~n28 ;
  assign n30 = x1 & ~x5 ;
  assign n31 = ~x1 & x5 ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = n32 ^ x6 ;
  assign n34 = x6 ^ x4 ;
  assign n35 = n34 ^ n33 ;
  assign n36 = ~x7 & ~x11 ;
  assign n37 = x13 & n36 ;
  assign n38 = ~x3 & n37 ;
  assign n39 = x7 & x13 ;
  assign n40 = ~x11 & n39 ;
  assign n41 = x3 & n40 ;
  assign n42 = ~n38 & ~n41 ;
  assign n43 = n42 ^ n32 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = ~x3 & n21 ;
  assign n46 = x12 & n45 ;
  assign n47 = ~x7 & x12 ;
  assign n48 = n24 & n47 ;
  assign n49 = ~n46 & ~n48 ;
  assign n50 = n49 ^ n42 ;
  assign n51 = ~n44 & n50 ;
  assign n52 = n51 ^ n42 ;
  assign n53 = n52 ^ n33 ;
  assign n54 = n35 & ~n53 ;
  assign n55 = n54 ^ n51 ;
  assign n56 = n55 ^ n42 ;
  assign n57 = n56 ^ n34 ;
  assign n58 = n33 & ~n57 ;
  assign n59 = n58 ^ n33 ;
  assign n60 = n59 ^ x2 ;
  assign n61 = n60 ^ n59 ;
  assign n62 = x7 ^ x5 ;
  assign n63 = n62 ^ n15 ;
  assign n64 = x10 ^ x5 ;
  assign n65 = n64 ^ x10 ;
  assign n66 = x11 ^ x10 ;
  assign n67 = ~n65 & n66 ;
  assign n68 = n67 ^ x10 ;
  assign n69 = n68 ^ n62 ;
  assign n70 = ~n63 & n69 ;
  assign n71 = n70 ^ n67 ;
  assign n72 = n71 ^ x10 ;
  assign n73 = n72 ^ n15 ;
  assign n74 = ~n62 & ~n73 ;
  assign n75 = n74 ^ n62 ;
  assign n76 = x4 & x5 ;
  assign n77 = x6 & n76 ;
  assign n78 = n38 & n77 ;
  assign n79 = ~x4 & ~x12 ;
  assign n80 = x3 & x13 ;
  assign n81 = ~n79 & n80 ;
  assign n82 = n81 ^ x12 ;
  assign n83 = x7 & n25 ;
  assign n84 = n83 ^ n81 ;
  assign n85 = n84 ^ n83 ;
  assign n86 = n85 ^ n82 ;
  assign n87 = ~x4 & ~x5 ;
  assign n88 = ~x6 & n87 ;
  assign n89 = n88 ^ n45 ;
  assign n90 = n45 & n89 ;
  assign n91 = n90 ^ n83 ;
  assign n92 = n91 ^ n45 ;
  assign n93 = ~n86 & ~n92 ;
  assign n94 = n93 ^ n90 ;
  assign n95 = n94 ^ n45 ;
  assign n96 = n82 & n95 ;
  assign n97 = n96 ^ n81 ;
  assign n98 = ~n78 & ~n97 ;
  assign n99 = ~x6 & x12 ;
  assign n100 = ~x7 & n99 ;
  assign n101 = n87 & n100 ;
  assign n102 = x3 & n101 ;
  assign n103 = n98 & ~n102 ;
  assign n104 = n103 ^ x1 ;
  assign n105 = n104 ^ n103 ;
  assign n106 = x4 & ~x5 ;
  assign n107 = x6 & n106 ;
  assign n114 = n40 & n107 ;
  assign n108 = n37 & n107 ;
  assign n109 = x5 & ~x6 ;
  assign n110 = ~x4 & n109 ;
  assign n111 = x12 & n21 ;
  assign n112 = n110 & n111 ;
  assign n113 = ~n108 & ~n112 ;
  assign n115 = n114 ^ n113 ;
  assign n116 = n115 ^ n113 ;
  assign n117 = ~x10 & n110 ;
  assign n118 = n47 & n117 ;
  assign n119 = n118 ^ n113 ;
  assign n120 = n119 ^ n113 ;
  assign n121 = ~n116 & ~n120 ;
  assign n122 = n121 ^ n113 ;
  assign n123 = x3 & n122 ;
  assign n124 = n123 ^ n113 ;
  assign n125 = n124 ^ n103 ;
  assign n126 = ~n105 & n125 ;
  assign n127 = n126 ^ n103 ;
  assign n128 = n75 & n127 ;
  assign n129 = n128 ^ n59 ;
  assign n130 = n61 & ~n129 ;
  assign n131 = n130 ^ n59 ;
  assign n132 = ~n29 & ~n131 ;
  assign n133 = x9 & ~n132 ;
  assign n134 = ~x3 & x11 ;
  assign n135 = n101 & ~n134 ;
  assign n136 = ~x12 & ~n76 ;
  assign n137 = n21 & ~n136 ;
  assign n138 = n137 ^ x12 ;
  assign n139 = n138 ^ x13 ;
  assign n140 = n36 ^ x6 ;
  assign n141 = n140 ^ n138 ;
  assign n142 = ~n137 & ~n141 ;
  assign n143 = n142 ^ x6 ;
  assign n144 = n143 ^ n137 ;
  assign n145 = n144 ^ n138 ;
  assign n146 = n145 ^ x13 ;
  assign n147 = n139 & n146 ;
  assign n148 = n147 ^ n142 ;
  assign n149 = n148 ^ x6 ;
  assign n150 = n149 ^ n138 ;
  assign n151 = x13 & ~n150 ;
  assign n152 = n151 ^ x13 ;
  assign n153 = n152 ^ x13 ;
  assign n154 = n98 & ~n153 ;
  assign n155 = ~n135 & n154 ;
  assign n156 = x1 & x2 ;
  assign n157 = ~x8 & n156 ;
  assign n158 = ~n155 & n157 ;
  assign n159 = ~n133 & ~n158 ;
  assign n160 = x0 & ~n159 ;
  assign n274 = x8 & n87 ;
  assign n275 = ~x0 & ~x1 ;
  assign n276 = x8 & x10 ;
  assign n277 = n275 & n276 ;
  assign n278 = ~n274 & ~n277 ;
  assign n279 = ~x8 & ~x10 ;
  assign n280 = n106 ^ x0 ;
  assign n281 = n280 ^ n106 ;
  assign n282 = n281 ^ n279 ;
  assign n198 = x5 & x13 ;
  assign n283 = ~x1 & x4 ;
  assign n284 = n283 ^ n279 ;
  assign n285 = n198 & ~n284 ;
  assign n286 = n285 ^ n106 ;
  assign n287 = n282 & n286 ;
  assign n288 = n287 ^ n285 ;
  assign n289 = ~n279 & n288 ;
  assign n290 = n289 ^ n285 ;
  assign n291 = n290 ^ n287 ;
  assign n292 = n278 & ~n291 ;
  assign n293 = x11 & ~n292 ;
  assign n294 = ~n274 & ~n276 ;
  assign n295 = ~x0 & x4 ;
  assign n296 = x0 & ~x4 ;
  assign n297 = ~n295 & ~n296 ;
  assign n298 = ~n32 & ~n297 ;
  assign n299 = ~n294 & n298 ;
  assign n300 = ~x8 & ~x11 ;
  assign n312 = ~x0 & ~x5 ;
  assign n301 = x5 & x10 ;
  assign n303 = ~x0 & ~x4 ;
  assign n302 = x0 & x4 ;
  assign n304 = n303 ^ n302 ;
  assign n305 = n304 ^ n303 ;
  assign n306 = n303 ^ x13 ;
  assign n307 = n306 ^ n303 ;
  assign n308 = n305 & n307 ;
  assign n309 = n308 ^ n303 ;
  assign n310 = ~n301 & n309 ;
  assign n311 = n310 ^ n303 ;
  assign n313 = n312 ^ n311 ;
  assign n314 = n313 ^ n311 ;
  assign n315 = x4 & x10 ;
  assign n316 = n315 ^ n311 ;
  assign n317 = n316 ^ n311 ;
  assign n318 = n314 & ~n317 ;
  assign n319 = n318 ^ n311 ;
  assign n320 = x1 & n319 ;
  assign n321 = n320 ^ n311 ;
  assign n322 = n300 & n321 ;
  assign n323 = ~n299 & ~n322 ;
  assign n324 = x3 & ~n323 ;
  assign n325 = x2 & n324 ;
  assign n326 = ~n293 & ~n325 ;
  assign n327 = ~x6 & ~x12 ;
  assign n328 = ~x7 & n327 ;
  assign n329 = ~n326 & n328 ;
  assign n330 = ~x3 & x10 ;
  assign n228 = ~x2 & ~x5 ;
  assign n229 = ~x1 & ~x6 ;
  assign n230 = ~n228 & ~n229 ;
  assign n331 = n79 & ~n230 ;
  assign n266 = ~x5 & ~x6 ;
  assign n332 = ~x0 & ~x12 ;
  assign n333 = n266 & n332 ;
  assign n334 = ~x2 & n275 ;
  assign n335 = ~n333 & ~n334 ;
  assign n336 = ~n331 & n335 ;
  assign n337 = x11 & ~n336 ;
  assign n338 = x8 & n337 ;
  assign n339 = n338 ^ x7 ;
  assign n340 = x6 & ~x12 ;
  assign n341 = ~x4 & ~n32 ;
  assign n342 = x8 & n341 ;
  assign n343 = x0 & n342 ;
  assign n344 = n340 & n343 ;
  assign n345 = n303 ^ n295 ;
  assign n346 = n345 ^ n295 ;
  assign n347 = n295 ^ x11 ;
  assign n348 = n347 ^ n295 ;
  assign n349 = n346 & ~n348 ;
  assign n350 = n349 ^ n295 ;
  assign n351 = ~x8 & n350 ;
  assign n352 = n351 ^ n295 ;
  assign n353 = ~n32 & n352 ;
  assign n233 = x1 & x12 ;
  assign n354 = x6 & ~n233 ;
  assign n355 = n353 & n354 ;
  assign n356 = x13 & n300 ;
  assign n262 = x1 & ~x6 ;
  assign n357 = ~n136 & n262 ;
  assign n238 = ~x1 & x6 ;
  assign n358 = ~x5 & n238 ;
  assign n359 = ~n79 & n358 ;
  assign n360 = ~n357 & ~n359 ;
  assign n361 = n356 & ~n360 ;
  assign n362 = x0 & n361 ;
  assign n363 = ~n355 & ~n362 ;
  assign n364 = ~n344 & n363 ;
  assign n365 = n364 ^ x2 ;
  assign n366 = n365 ^ n364 ;
  assign n367 = x0 & ~x1 ;
  assign n368 = n106 & n356 ;
  assign n369 = n367 & n368 ;
  assign n370 = ~n353 & ~n369 ;
  assign n371 = ~n343 & n370 ;
  assign n372 = n327 & ~n371 ;
  assign n373 = n372 ^ n364 ;
  assign n374 = n366 & ~n373 ;
  assign n375 = n374 ^ n364 ;
  assign n376 = n375 ^ n338 ;
  assign n377 = ~n339 & n376 ;
  assign n378 = n377 ^ n374 ;
  assign n379 = n378 ^ n364 ;
  assign n380 = n379 ^ x7 ;
  assign n381 = ~n338 & ~n380 ;
  assign n382 = n381 ^ n338 ;
  assign n383 = n382 ^ n338 ;
  assign n384 = n330 & ~n383 ;
  assign n385 = ~n329 & ~n384 ;
  assign n209 = x6 ^ x2 ;
  assign n386 = n32 & ~n209 ;
  assign n387 = ~n275 & n386 ;
  assign n388 = x2 & n358 ;
  assign n389 = ~x4 & n388 ;
  assign n390 = ~n387 & ~n389 ;
  assign n391 = ~x7 & x8 ;
  assign n392 = n297 & n391 ;
  assign n393 = ~n390 & n392 ;
  assign n394 = x10 ^ x8 ;
  assign n395 = ~x0 & n25 ;
  assign n239 = ~x2 & x5 ;
  assign n240 = ~n238 & ~n239 ;
  assign n396 = x4 & ~n240 ;
  assign n397 = ~n395 & ~n396 ;
  assign n398 = n397 ^ x10 ;
  assign n399 = n398 ^ n397 ;
  assign n400 = n399 ^ n394 ;
  assign n401 = x1 & ~n209 ;
  assign n402 = x5 & n401 ;
  assign n403 = ~n388 & ~n402 ;
  assign n404 = n295 & ~n403 ;
  assign n161 = x2 & x6 ;
  assign n405 = x12 & n296 ;
  assign n406 = n161 & n405 ;
  assign n407 = n31 & n406 ;
  assign n408 = ~n404 & ~n407 ;
  assign n409 = n408 ^ x7 ;
  assign n410 = ~x7 & n409 ;
  assign n411 = n410 ^ n397 ;
  assign n412 = n411 ^ x7 ;
  assign n413 = n400 & n412 ;
  assign n414 = n413 ^ n410 ;
  assign n415 = n414 ^ x7 ;
  assign n416 = ~n394 & ~n415 ;
  assign n417 = ~n393 & ~n416 ;
  assign n418 = n134 & ~n417 ;
  assign n419 = x3 & ~x12 ;
  assign n244 = x2 & x5 ;
  assign n245 = ~n22 & ~n244 ;
  assign n436 = ~n245 & n315 ;
  assign n437 = ~x6 & x11 ;
  assign n438 = ~n301 & ~n437 ;
  assign n439 = ~n109 & ~n438 ;
  assign n440 = ~n156 & ~n439 ;
  assign n441 = x0 & ~n440 ;
  assign n263 = x2 & ~x5 ;
  assign n264 = ~n262 & ~n263 ;
  assign n442 = ~x4 & x11 ;
  assign n443 = ~n264 & n442 ;
  assign n444 = ~n441 & ~n443 ;
  assign n445 = ~n436 & n444 ;
  assign n420 = x10 & ~x11 ;
  assign n421 = ~x4 & n420 ;
  assign n422 = ~n245 & n421 ;
  assign n423 = ~x5 & x11 ;
  assign n424 = x2 & x4 ;
  assign n425 = n423 & n424 ;
  assign n426 = x11 ^ x2 ;
  assign n427 = n426 ^ x2 ;
  assign n428 = x4 & ~x6 ;
  assign n429 = n428 ^ x2 ;
  assign n430 = n427 & n429 ;
  assign n431 = n430 ^ x2 ;
  assign n432 = x1 & n431 ;
  assign n433 = ~n425 & ~n432 ;
  assign n434 = ~x10 & ~n433 ;
  assign n435 = ~n422 & ~n434 ;
  assign n446 = n445 ^ n435 ;
  assign n447 = n446 ^ n445 ;
  assign n448 = n445 ^ x0 ;
  assign n449 = n448 ^ n445 ;
  assign n450 = ~n447 & ~n449 ;
  assign n451 = n450 ^ n445 ;
  assign n452 = ~x8 & ~n451 ;
  assign n453 = n452 ^ n445 ;
  assign n454 = n419 & ~n453 ;
  assign n455 = x8 ^ x0 ;
  assign n456 = n455 ^ x8 ;
  assign n457 = n279 ^ x8 ;
  assign n458 = n457 ^ x8 ;
  assign n459 = ~n456 & n458 ;
  assign n460 = n459 ^ x8 ;
  assign n461 = x4 & n460 ;
  assign n462 = n461 ^ x8 ;
  assign n463 = n156 & n462 ;
  assign n464 = x0 & x8 ;
  assign n465 = ~n264 & n464 ;
  assign n466 = ~n463 & ~n465 ;
  assign n467 = ~x7 & ~n466 ;
  assign n468 = ~n276 & ~n467 ;
  assign n469 = x11 & ~x12 ;
  assign n470 = ~n468 & n469 ;
  assign n471 = ~n454 & ~n470 ;
  assign n472 = n332 ^ n156 ;
  assign n473 = n472 ^ n332 ;
  assign n474 = n473 ^ n395 ;
  assign n475 = x0 & x12 ;
  assign n476 = x6 ^ x1 ;
  assign n477 = n475 & n476 ;
  assign n478 = n477 ^ x5 ;
  assign n479 = ~x5 & ~n478 ;
  assign n480 = n479 ^ n332 ;
  assign n481 = n480 ^ x5 ;
  assign n482 = n474 & ~n481 ;
  assign n483 = n482 ^ n479 ;
  assign n484 = n483 ^ x5 ;
  assign n485 = ~n395 & ~n484 ;
  assign n486 = n485 ^ n395 ;
  assign n487 = n421 & n486 ;
  assign n488 = n423 ^ x1 ;
  assign n489 = n488 ^ n423 ;
  assign n490 = n489 ^ n209 ;
  assign n491 = n16 ^ x5 ;
  assign n492 = ~n16 & ~n491 ;
  assign n493 = n492 ^ n423 ;
  assign n494 = n493 ^ n16 ;
  assign n495 = ~n490 & ~n494 ;
  assign n496 = n495 ^ n492 ;
  assign n497 = n496 ^ n16 ;
  assign n498 = ~n209 & ~n497 ;
  assign n499 = n295 & n498 ;
  assign n500 = n156 & n395 ;
  assign n501 = ~x11 & n500 ;
  assign n502 = n238 & ~n423 ;
  assign n503 = x2 & ~n502 ;
  assign n504 = n405 & ~n503 ;
  assign n505 = x5 ^ x1 ;
  assign n506 = n437 ^ x5 ;
  assign n507 = n505 & ~n506 ;
  assign n508 = ~x2 & n507 ;
  assign n509 = n508 ^ x2 ;
  assign n510 = n504 & n509 ;
  assign n511 = ~n501 & ~n510 ;
  assign n512 = ~n499 & n511 ;
  assign n513 = n24 & ~n512 ;
  assign n514 = ~n487 & ~n513 ;
  assign n515 = n514 ^ x8 ;
  assign n516 = n515 ^ n514 ;
  assign n517 = x4 ^ x0 ;
  assign n518 = n498 ^ x4 ;
  assign n519 = n518 ^ n498 ;
  assign n520 = n519 ^ n517 ;
  assign n521 = n386 ^ x11 ;
  assign n522 = n386 & n521 ;
  assign n523 = n522 ^ n498 ;
  assign n524 = n523 ^ n386 ;
  assign n525 = n520 & n524 ;
  assign n526 = n525 ^ n522 ;
  assign n527 = n526 ^ n386 ;
  assign n528 = ~n517 & n527 ;
  assign n529 = x3 & n528 ;
  assign n530 = ~x0 & ~n240 ;
  assign n531 = ~x2 & n283 ;
  assign n532 = ~n530 & ~n531 ;
  assign n533 = x11 & ~n532 ;
  assign n534 = ~n77 & ~n533 ;
  assign n535 = x10 & ~n534 ;
  assign n536 = x10 & ~x12 ;
  assign n537 = x0 & ~n245 ;
  assign n538 = x1 & n424 ;
  assign n539 = ~n537 & ~n538 ;
  assign n540 = n536 & ~n539 ;
  assign n541 = ~n535 & ~n540 ;
  assign n542 = ~n529 & n541 ;
  assign n543 = n542 ^ n514 ;
  assign n544 = n516 & n543 ;
  assign n545 = n544 ^ n514 ;
  assign n546 = x7 & ~n545 ;
  assign n547 = n471 & ~n546 ;
  assign n548 = ~n418 & n547 ;
  assign n549 = ~x13 & ~n548 ;
  assign n550 = n385 & ~n549 ;
  assign n162 = ~n42 & n87 ;
  assign n163 = n161 & n162 ;
  assign n164 = ~x10 & ~x11 ;
  assign n165 = n39 ^ x6 ;
  assign n166 = n165 ^ n39 ;
  assign n167 = n166 ^ n164 ;
  assign n168 = n47 ^ n39 ;
  assign n169 = ~n167 & n168 ;
  assign n170 = n169 ^ n47 ;
  assign n171 = n164 & n170 ;
  assign n172 = ~n163 & ~n171 ;
  assign n173 = x4 & n109 ;
  assign n174 = ~n49 & n173 ;
  assign n175 = n174 ^ x2 ;
  assign n176 = n175 ^ n174 ;
  assign n177 = ~n45 & ~n48 ;
  assign n178 = n77 & ~n177 ;
  assign n179 = n36 & n88 ;
  assign n180 = ~n164 & ~n179 ;
  assign n181 = n180 ^ x3 ;
  assign n182 = n181 ^ n180 ;
  assign n183 = n182 ^ n178 ;
  assign n184 = n88 ^ n40 ;
  assign n185 = n88 & n184 ;
  assign n186 = n185 ^ n180 ;
  assign n187 = n186 ^ n88 ;
  assign n188 = ~n183 & ~n187 ;
  assign n189 = n188 ^ n185 ;
  assign n190 = n189 ^ n88 ;
  assign n191 = ~n178 & n190 ;
  assign n192 = n191 ^ n178 ;
  assign n193 = n192 ^ n174 ;
  assign n194 = ~n176 & n193 ;
  assign n195 = n194 ^ n174 ;
  assign n196 = n172 & ~n195 ;
  assign n197 = ~x1 & ~n196 ;
  assign n199 = ~n99 & ~n198 ;
  assign n200 = ~x3 & ~n109 ;
  assign n201 = ~n199 & n200 ;
  assign n202 = n39 ^ x5 ;
  assign n203 = n202 ^ n39 ;
  assign n204 = n168 & ~n203 ;
  assign n205 = n204 ^ n39 ;
  assign n206 = ~x2 & n205 ;
  assign n207 = ~n201 & ~n206 ;
  assign n208 = n164 & ~n207 ;
  assign n210 = ~n49 & n106 ;
  assign n211 = n210 ^ n209 ;
  assign n212 = n211 ^ n210 ;
  assign n213 = ~x4 & x5 ;
  assign n214 = ~n42 & n213 ;
  assign n215 = n214 ^ n210 ;
  assign n216 = ~n212 & n215 ;
  assign n217 = n216 ^ n210 ;
  assign n218 = x1 & n217 ;
  assign n219 = ~n208 & ~n218 ;
  assign n220 = ~n197 & n219 ;
  assign n221 = ~x0 & ~n220 ;
  assign n222 = ~x11 & x12 ;
  assign n223 = n222 ^ x13 ;
  assign n224 = n222 ^ x4 ;
  assign n225 = n224 ^ n223 ;
  assign n234 = x2 & x7 ;
  assign n235 = n233 & n234 ;
  assign n236 = ~x2 & x7 ;
  assign n237 = ~x1 & n236 ;
  assign n241 = ~x3 & ~n240 ;
  assign n242 = ~n237 & ~n241 ;
  assign n243 = ~x11 & ~n242 ;
  assign n246 = x3 & x12 ;
  assign n247 = ~n245 & n246 ;
  assign n248 = ~n83 & ~n247 ;
  assign n249 = ~n243 & n248 ;
  assign n250 = ~n235 & n249 ;
  assign n226 = ~x2 & ~x7 ;
  assign n227 = ~x1 & n226 ;
  assign n231 = ~x3 & ~n230 ;
  assign n232 = ~n227 & ~n231 ;
  assign n251 = n250 ^ n232 ;
  assign n252 = ~x4 & n251 ;
  assign n253 = n252 ^ n250 ;
  assign n254 = n225 & n253 ;
  assign n255 = n254 ^ n252 ;
  assign n256 = n255 ^ n250 ;
  assign n257 = n256 ^ x4 ;
  assign n258 = n223 & ~n257 ;
  assign n259 = n258 ^ x13 ;
  assign n260 = ~x10 & n259 ;
  assign n261 = ~x4 & n222 ;
  assign n265 = n80 & ~n264 ;
  assign n267 = x13 & n156 ;
  assign n268 = ~n266 & ~n267 ;
  assign n269 = ~x7 & ~n268 ;
  assign n270 = ~n265 & ~n269 ;
  assign n271 = n261 & ~n270 ;
  assign n272 = ~n260 & ~n271 ;
  assign n273 = ~n221 & n272 ;
  assign n551 = n550 ^ n273 ;
  assign n552 = n551 ^ n273 ;
  assign n553 = n340 & n420 ;
  assign n554 = n303 & n553 ;
  assign n555 = n17 & n554 ;
  assign n556 = ~n134 & ~n419 ;
  assign n557 = x6 & x10 ;
  assign n558 = x0 & ~n557 ;
  assign n559 = ~n556 & n558 ;
  assign n560 = ~x13 & ~n87 ;
  assign n561 = ~n136 & ~n560 ;
  assign n562 = n559 & n561 ;
  assign n563 = ~n437 & n562 ;
  assign n564 = ~n555 & ~n563 ;
  assign n565 = x1 & ~n564 ;
  assign n566 = x4 & ~x13 ;
  assign n567 = n367 & ~n566 ;
  assign n570 = n80 & n536 ;
  assign n571 = n107 & n570 ;
  assign n568 = x5 & ~x10 ;
  assign n569 = n99 & n568 ;
  assign n572 = n571 ^ n569 ;
  assign n573 = n572 ^ n571 ;
  assign n574 = n571 ^ x3 ;
  assign n575 = n574 ^ n571 ;
  assign n576 = n573 & ~n575 ;
  assign n577 = n576 ^ n571 ;
  assign n578 = x11 & n577 ;
  assign n579 = n578 ^ n571 ;
  assign n580 = n567 & n579 ;
  assign n581 = n275 & ~n315 ;
  assign n582 = n134 & n266 ;
  assign n585 = n582 ^ n553 ;
  assign n586 = n585 ^ n582 ;
  assign n583 = n582 ^ x5 ;
  assign n584 = n583 ^ n582 ;
  assign n587 = n586 ^ n584 ;
  assign n588 = n582 ^ x3 ;
  assign n589 = n588 ^ n582 ;
  assign n590 = n589 ^ n586 ;
  assign n591 = n586 & n590 ;
  assign n592 = n591 ^ n586 ;
  assign n593 = n587 & n592 ;
  assign n594 = n593 ^ n591 ;
  assign n595 = n594 ^ n582 ;
  assign n596 = n595 ^ n586 ;
  assign n597 = ~x4 & n596 ;
  assign n598 = n597 ^ n582 ;
  assign n599 = n581 & n598 ;
  assign n600 = ~x8 & ~n599 ;
  assign n601 = ~n580 & n600 ;
  assign n602 = ~n565 & n601 ;
  assign n603 = x11 & n312 ;
  assign n604 = ~x1 & n442 ;
  assign n605 = ~n603 & ~n604 ;
  assign n606 = x3 & x6 ;
  assign n607 = n298 & n606 ;
  assign n608 = n605 & ~n607 ;
  assign n609 = n536 & ~n608 ;
  assign n610 = n229 & n442 ;
  assign n611 = n312 & n610 ;
  assign n612 = ~x3 & n611 ;
  assign n613 = x8 & ~n612 ;
  assign n614 = ~n609 & n613 ;
  assign n615 = n226 & ~n614 ;
  assign n616 = ~n602 & n615 ;
  assign n617 = n616 ^ n273 ;
  assign n618 = n617 ^ n273 ;
  assign n619 = n552 & ~n618 ;
  assign n620 = n619 ^ n273 ;
  assign n621 = ~x9 & n620 ;
  assign n622 = n621 ^ n273 ;
  assign n623 = ~n160 & n622 ;
  assign y0 = ~n623 ;
endmodule
