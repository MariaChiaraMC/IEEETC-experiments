module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 ;
  assign n17 = ~x2 & ~x3 ;
  assign n18 = ~x0 & n17 ;
  assign n19 = ~x8 & n18 ;
  assign n20 = x1 & n19 ;
  assign n21 = ~x9 & ~x10 ;
  assign n22 = n21 ^ x7 ;
  assign n23 = n22 ^ n21 ;
  assign n24 = n23 ^ x6 ;
  assign n25 = n21 ^ x4 ;
  assign n26 = n21 ^ x5 ;
  assign n27 = n26 ^ n25 ;
  assign n28 = ~n25 & ~n27 ;
  assign n29 = n28 ^ n21 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = n24 & n30 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = n32 ^ n25 ;
  assign n34 = ~x6 & ~n33 ;
  assign n35 = n34 ^ n21 ;
  assign n36 = n20 & ~n35 ;
  assign n37 = x10 ^ x9 ;
  assign n38 = x13 & ~x15 ;
  assign n39 = ~x11 & ~x12 ;
  assign n40 = n38 & n39 ;
  assign n41 = ~x14 & n40 ;
  assign n42 = n41 ^ x7 ;
  assign n44 = n42 ^ n41 ;
  assign n43 = n42 ^ x9 ;
  assign n45 = n44 ^ n43 ;
  assign n46 = n45 ^ n37 ;
  assign n47 = ~n37 & n46 ;
  assign n48 = n47 ^ n42 ;
  assign n49 = n48 ^ n37 ;
  assign n50 = n42 ^ x5 ;
  assign n51 = n44 & ~n50 ;
  assign n52 = n51 ^ n42 ;
  assign n53 = n49 & ~n52 ;
  assign n54 = n53 ^ n42 ;
  assign n55 = n54 ^ n41 ;
  assign n56 = n36 & ~n55 ;
  assign y0 = n56 ;
endmodule
