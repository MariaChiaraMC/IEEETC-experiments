module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 ;
  assign n15 = ~x4 & x8 ;
  assign n16 = x0 & x2 ;
  assign n17 = x1 & n16 ;
  assign n18 = n15 & n17 ;
  assign n19 = ~x7 & n18 ;
  assign n20 = ~x5 & ~x11 ;
  assign n21 = x5 & ~x10 ;
  assign n22 = ~n20 & ~n21 ;
  assign n23 = ~x12 & ~n22 ;
  assign n24 = x2 & ~x6 ;
  assign n25 = x6 & n20 ;
  assign n26 = x4 & x8 ;
  assign n27 = ~n21 & ~n26 ;
  assign n28 = ~n25 & n27 ;
  assign n29 = x7 & ~n28 ;
  assign n30 = ~n24 & n29 ;
  assign n31 = ~n23 & ~n30 ;
  assign n32 = ~x1 & ~n31 ;
  assign n33 = ~x4 & ~x11 ;
  assign n34 = x5 & x6 ;
  assign n35 = n33 & n34 ;
  assign n36 = x4 & ~x10 ;
  assign n37 = ~x8 & ~n36 ;
  assign n38 = x1 & ~x5 ;
  assign n39 = ~n24 & ~n38 ;
  assign n40 = ~n37 & n39 ;
  assign n41 = ~n35 & ~n40 ;
  assign n42 = x7 & ~n41 ;
  assign n43 = ~n33 & ~n36 ;
  assign n44 = ~x12 & ~n43 ;
  assign n45 = ~n42 & ~n44 ;
  assign n46 = ~x0 & ~n45 ;
  assign n47 = ~x6 & x11 ;
  assign n48 = ~x2 & ~n47 ;
  assign n49 = x6 & x10 ;
  assign n50 = n48 & ~n49 ;
  assign n51 = ~n24 & n26 ;
  assign n52 = x5 & n51 ;
  assign n53 = ~n50 & ~n52 ;
  assign n54 = x7 & ~n53 ;
  assign n55 = x8 & ~x12 ;
  assign n56 = ~n54 & ~n55 ;
  assign n57 = ~n46 & n56 ;
  assign n58 = ~n32 & n57 ;
  assign n59 = ~n19 & n58 ;
  assign n60 = ~x13 & ~n59 ;
  assign n61 = ~x1 & ~x6 ;
  assign n62 = x2 & ~n61 ;
  assign n63 = x4 & ~x8 ;
  assign n64 = x1 & x5 ;
  assign n65 = ~x8 & x11 ;
  assign n66 = ~n64 & ~n65 ;
  assign n67 = ~n63 & n66 ;
  assign n68 = ~n62 & n67 ;
  assign n69 = ~x5 & ~x6 ;
  assign n70 = ~n37 & n69 ;
  assign n71 = ~n68 & ~n70 ;
  assign n72 = ~x7 & ~n71 ;
  assign n73 = ~x7 & ~x11 ;
  assign n74 = ~x4 & ~x5 ;
  assign n75 = ~x6 & n74 ;
  assign n76 = n73 & n75 ;
  assign n77 = ~n72 & ~n76 ;
  assign n78 = ~x0 & ~n77 ;
  assign n79 = ~x12 & n78 ;
  assign n80 = ~x2 & ~x6 ;
  assign n81 = ~x11 & n80 ;
  assign n82 = x2 & x6 ;
  assign n83 = ~x1 & n20 ;
  assign n84 = n15 & ~n64 ;
  assign n85 = ~n83 & ~n84 ;
  assign n86 = ~x2 & x6 ;
  assign n87 = ~x5 & ~n86 ;
  assign n88 = x1 & ~x6 ;
  assign n89 = ~n87 & ~n88 ;
  assign n90 = ~x10 & n89 ;
  assign n91 = n85 & ~n90 ;
  assign n92 = ~n82 & ~n91 ;
  assign n93 = ~n81 & ~n92 ;
  assign n94 = ~x7 & ~x12 ;
  assign n95 = ~n93 & n94 ;
  assign n96 = ~n79 & ~n95 ;
  assign n97 = ~n60 & n96 ;
  assign n98 = x3 & ~n97 ;
  assign n99 = ~x0 & x4 ;
  assign n100 = ~x10 & n99 ;
  assign n101 = n69 & n100 ;
  assign n102 = x13 & ~n101 ;
  assign n103 = ~x8 & ~n99 ;
  assign n104 = ~x8 & x10 ;
  assign n105 = ~n103 & ~n104 ;
  assign n106 = ~n102 & n105 ;
  assign n107 = ~x0 & ~x5 ;
  assign n108 = x8 & n107 ;
  assign n109 = ~n84 & ~n108 ;
  assign n110 = ~n82 & ~n109 ;
  assign n111 = ~x0 & x8 ;
  assign n112 = ~n21 & ~n111 ;
  assign n113 = n61 & ~n112 ;
  assign n114 = ~n110 & ~n113 ;
  assign n115 = ~n106 & n114 ;
  assign n116 = x11 & n94 ;
  assign n117 = ~n115 & n116 ;
  assign n118 = x0 & ~x4 ;
  assign n119 = x8 & ~n118 ;
  assign n120 = n119 ^ x1 ;
  assign n121 = n119 ^ x5 ;
  assign n122 = n121 ^ x5 ;
  assign n123 = n25 ^ x5 ;
  assign n124 = ~n122 & ~n123 ;
  assign n125 = n124 ^ x5 ;
  assign n126 = ~n120 & n125 ;
  assign n127 = n126 ^ x1 ;
  assign n128 = ~n24 & ~n127 ;
  assign n129 = ~n75 & n128 ;
  assign n130 = ~x0 & n33 ;
  assign n131 = n130 ^ x12 ;
  assign n132 = n130 ^ x8 ;
  assign n133 = n132 ^ x8 ;
  assign n134 = n34 ^ x8 ;
  assign n135 = n133 & ~n134 ;
  assign n136 = n135 ^ x8 ;
  assign n137 = ~n131 & ~n136 ;
  assign n138 = n137 ^ x12 ;
  assign n139 = ~n129 & n138 ;
  assign n140 = x7 & ~x13 ;
  assign n141 = x10 & n140 ;
  assign n142 = ~n139 & n141 ;
  assign n143 = ~n117 & ~n142 ;
  assign n144 = ~n98 & n143 ;
  assign n145 = ~x9 & ~n144 ;
  assign n146 = x12 ^ x3 ;
  assign n147 = x5 & n49 ;
  assign n148 = ~n63 & ~n118 ;
  assign n149 = n147 & ~n148 ;
  assign n150 = ~x2 & ~n49 ;
  assign n151 = n38 & ~n150 ;
  assign n152 = ~n149 & ~n151 ;
  assign n153 = ~x4 & n17 ;
  assign n154 = ~n24 & ~n153 ;
  assign n155 = n152 & n154 ;
  assign n156 = n73 & ~n155 ;
  assign n157 = n156 ^ n146 ;
  assign n158 = n157 ^ x12 ;
  assign n159 = n158 ^ n157 ;
  assign n167 = ~x4 & x12 ;
  assign n160 = x4 & x10 ;
  assign n161 = x5 & ~n80 ;
  assign n162 = x1 & x6 ;
  assign n163 = ~n161 & ~n162 ;
  assign n164 = n160 & ~n163 ;
  assign n168 = n167 ^ n164 ;
  assign n169 = n168 ^ n164 ;
  assign n165 = n164 ^ n89 ;
  assign n166 = n165 ^ n164 ;
  assign n170 = n169 ^ n166 ;
  assign n171 = n164 ^ x11 ;
  assign n172 = n171 ^ n164 ;
  assign n173 = n172 ^ n169 ;
  assign n174 = n169 & n173 ;
  assign n175 = n174 ^ n169 ;
  assign n176 = ~n170 & n175 ;
  assign n177 = n176 ^ n174 ;
  assign n178 = n177 ^ n164 ;
  assign n179 = n178 ^ n169 ;
  assign n180 = ~x7 & n179 ;
  assign n181 = n180 ^ n164 ;
  assign n182 = ~n111 & n181 ;
  assign n183 = ~x8 & n17 ;
  assign n184 = ~x9 & ~n183 ;
  assign n185 = x10 & n65 ;
  assign n186 = n184 & ~n185 ;
  assign n187 = n186 ^ x7 ;
  assign n188 = n187 ^ n182 ;
  assign n189 = ~n74 & ~n107 ;
  assign n190 = x2 & n189 ;
  assign n191 = x5 & n47 ;
  assign n192 = ~n147 & ~n191 ;
  assign n193 = n104 & n192 ;
  assign n194 = x0 & x6 ;
  assign n195 = n194 ^ n192 ;
  assign n196 = x2 & ~n74 ;
  assign n197 = n196 ^ n193 ;
  assign n198 = ~n195 & n197 ;
  assign n199 = n198 ^ n196 ;
  assign n200 = n193 & n199 ;
  assign n201 = n200 ^ n192 ;
  assign n202 = ~n190 & n201 ;
  assign n203 = x1 & ~n202 ;
  assign n204 = n104 & n161 ;
  assign n205 = x11 & n160 ;
  assign n206 = ~n204 & ~n205 ;
  assign n207 = x0 & ~n206 ;
  assign n208 = ~n82 & ~n207 ;
  assign n209 = ~n203 & n208 ;
  assign n210 = n209 ^ x12 ;
  assign n211 = n186 & n210 ;
  assign n212 = n211 ^ x12 ;
  assign n213 = n188 & ~n212 ;
  assign n214 = n213 ^ n211 ;
  assign n215 = n214 ^ x12 ;
  assign n216 = n215 ^ n186 ;
  assign n217 = ~n182 & ~n216 ;
  assign n218 = ~n140 & ~n217 ;
  assign n219 = n218 ^ n157 ;
  assign n220 = n219 ^ n146 ;
  assign n221 = n159 & ~n220 ;
  assign n222 = n221 ^ n218 ;
  assign n223 = ~x7 & x11 ;
  assign n224 = x0 & ~x6 ;
  assign n225 = x2 & ~x4 ;
  assign n226 = ~n224 & ~n225 ;
  assign n227 = ~x8 & ~n226 ;
  assign n228 = ~n69 & ~n227 ;
  assign n229 = x1 & ~n228 ;
  assign n230 = x0 & ~x8 ;
  assign n231 = n87 & n230 ;
  assign n232 = x10 & n118 ;
  assign n233 = ~n231 & ~n232 ;
  assign n234 = ~n229 & n233 ;
  assign n235 = n223 & ~n234 ;
  assign n236 = ~x1 & ~x2 ;
  assign n237 = ~n50 & ~n236 ;
  assign n238 = x11 ^ x10 ;
  assign n239 = n238 ^ x0 ;
  assign n240 = x10 ^ x5 ;
  assign n241 = x10 ^ x6 ;
  assign n242 = n241 ^ n240 ;
  assign n243 = ~n240 & n242 ;
  assign n244 = n243 ^ x10 ;
  assign n245 = n244 ^ n240 ;
  assign n246 = n239 & ~n245 ;
  assign n247 = n246 ^ n243 ;
  assign n248 = n247 ^ n240 ;
  assign n249 = x0 & ~n248 ;
  assign n250 = ~n237 & ~n249 ;
  assign n251 = x13 & ~n250 ;
  assign n252 = x6 & ~n38 ;
  assign n253 = ~n150 & ~n252 ;
  assign n254 = ~x7 & n253 ;
  assign n255 = ~n251 & ~n254 ;
  assign n256 = ~n235 & n255 ;
  assign n257 = ~n218 & n256 ;
  assign n258 = n257 ^ n146 ;
  assign n259 = ~n222 & ~n258 ;
  assign n260 = n259 ^ n257 ;
  assign n261 = ~n146 & n260 ;
  assign n262 = n261 ^ n221 ;
  assign n263 = n262 ^ x3 ;
  assign n264 = n263 ^ n218 ;
  assign n265 = ~n145 & n264 ;
  assign n266 = ~x10 & n86 ;
  assign n267 = x5 & ~n118 ;
  assign n268 = n105 & n267 ;
  assign n269 = ~n100 & n112 ;
  assign n270 = ~n26 & n269 ;
  assign n271 = ~x1 & ~n270 ;
  assign n272 = ~n268 & ~n271 ;
  assign n273 = n236 & ~n269 ;
  assign n274 = x13 & ~n273 ;
  assign n275 = ~n24 & ~n274 ;
  assign n276 = ~n272 & n275 ;
  assign n277 = ~n266 & ~n276 ;
  assign n278 = n223 & ~n277 ;
  assign n279 = ~x9 & n278 ;
  assign n290 = x4 & ~n224 ;
  assign n291 = n65 & ~n290 ;
  assign n292 = ~n86 & n291 ;
  assign n293 = x12 & ~n267 ;
  assign n294 = ~n48 & n293 ;
  assign n295 = ~n292 & ~n294 ;
  assign n296 = x1 & ~n295 ;
  assign n297 = x12 & n24 ;
  assign n298 = n184 & ~n297 ;
  assign n299 = x12 & n118 ;
  assign n300 = ~n103 & ~n299 ;
  assign n301 = n87 & ~n300 ;
  assign n302 = x11 & n301 ;
  assign n303 = n298 & ~n302 ;
  assign n304 = ~n296 & n303 ;
  assign n280 = ~x12 & ~n82 ;
  assign n281 = ~x0 & ~n63 ;
  assign n282 = ~n65 & n281 ;
  assign n283 = ~n20 & ~n282 ;
  assign n284 = n236 & ~n283 ;
  assign n285 = ~n280 & ~n284 ;
  assign n286 = ~x0 & n67 ;
  assign n287 = n85 & ~n286 ;
  assign n288 = ~n285 & ~n287 ;
  assign n289 = ~n81 & ~n288 ;
  assign n305 = n304 ^ n289 ;
  assign n306 = n305 ^ n304 ;
  assign n307 = n304 ^ x9 ;
  assign n308 = n307 ^ n304 ;
  assign n309 = ~n306 & ~n308 ;
  assign n310 = n309 ^ n304 ;
  assign n311 = x10 & ~n310 ;
  assign n312 = n311 ^ n304 ;
  assign n313 = n312 ^ x7 ;
  assign n314 = n313 ^ n312 ;
  assign n315 = n314 ^ n279 ;
  assign n316 = x4 & x13 ;
  assign n317 = x8 & ~n316 ;
  assign n318 = x10 & ~n317 ;
  assign n319 = n161 & n318 ;
  assign n320 = ~n281 & n319 ;
  assign n321 = x13 & ~n150 ;
  assign n322 = n189 & n321 ;
  assign n323 = ~x4 & ~n194 ;
  assign n324 = n104 & ~n323 ;
  assign n325 = ~n80 & n324 ;
  assign n326 = ~n322 & ~n325 ;
  assign n327 = x1 & ~n326 ;
  assign n328 = x13 & n82 ;
  assign n329 = n184 & ~n328 ;
  assign n330 = ~n327 & n329 ;
  assign n331 = ~n320 & n330 ;
  assign n332 = n331 ^ x11 ;
  assign n333 = ~x11 & n332 ;
  assign n334 = n333 ^ n312 ;
  assign n335 = n334 ^ x11 ;
  assign n336 = n315 & n335 ;
  assign n337 = n336 ^ n333 ;
  assign n338 = n337 ^ x11 ;
  assign n339 = ~n279 & ~n338 ;
  assign n340 = n339 ^ n279 ;
  assign n341 = ~x3 & n340 ;
  assign n342 = ~n190 & ~n191 ;
  assign n343 = x1 & ~n342 ;
  assign n344 = ~n15 & ~n99 ;
  assign n345 = x11 & n69 ;
  assign n346 = n344 & n345 ;
  assign n347 = ~n82 & ~n346 ;
  assign n348 = ~n343 & n347 ;
  assign n349 = ~x10 & x13 ;
  assign n350 = x7 & n349 ;
  assign n351 = ~n348 & n350 ;
  assign n352 = ~n341 & ~n351 ;
  assign n353 = n265 & n352 ;
  assign y0 = ~n353 ;
endmodule
