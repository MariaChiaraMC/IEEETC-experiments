module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 ;
  assign n16 = x7 & x13 ;
  assign n17 = ~x5 & n16 ;
  assign n18 = x1 & n17 ;
  assign n19 = x5 & ~x9 ;
  assign n20 = ~x1 & ~x6 ;
  assign n21 = x8 & ~x13 ;
  assign n22 = ~n20 & n21 ;
  assign n23 = n19 & n22 ;
  assign n24 = x14 & n23 ;
  assign n25 = x5 & ~x7 ;
  assign n26 = x14 ^ x13 ;
  assign n27 = x14 ^ x10 ;
  assign n28 = n27 ^ x10 ;
  assign n29 = x10 ^ x9 ;
  assign n30 = n28 & ~n29 ;
  assign n31 = n30 ^ x10 ;
  assign n32 = ~n26 & n31 ;
  assign n33 = ~n25 & n32 ;
  assign n34 = ~n24 & ~n33 ;
  assign n35 = ~n18 & n34 ;
  assign n36 = x3 & ~n35 ;
  assign n37 = x10 & ~x14 ;
  assign n38 = x10 & ~x13 ;
  assign n39 = x7 & n38 ;
  assign n40 = ~n37 & ~n39 ;
  assign n41 = ~x5 & n38 ;
  assign n42 = ~n17 & ~n41 ;
  assign n43 = n40 & n42 ;
  assign n44 = x9 & ~n43 ;
  assign n45 = ~n36 & ~n44 ;
  assign n46 = x4 & ~n45 ;
  assign n47 = x9 & n37 ;
  assign n50 = ~x13 & n47 ;
  assign n51 = ~x7 & n50 ;
  assign n48 = ~x7 & ~x8 ;
  assign n49 = n47 & ~n48 ;
  assign n52 = n51 ^ n49 ;
  assign n53 = n52 ^ n49 ;
  assign n54 = ~x4 & ~x10 ;
  assign n55 = x3 & n54 ;
  assign n56 = x8 ^ x7 ;
  assign n57 = n55 & n56 ;
  assign n58 = n57 ^ n49 ;
  assign n59 = n58 ^ n49 ;
  assign n60 = ~n53 & ~n59 ;
  assign n61 = n60 ^ n49 ;
  assign n62 = x6 & ~n61 ;
  assign n63 = n62 ^ n49 ;
  assign n64 = ~x5 & n63 ;
  assign n65 = ~n46 & ~n64 ;
  assign n66 = ~x0 & ~n65 ;
  assign n67 = ~x9 & ~x10 ;
  assign n68 = x1 & x13 ;
  assign n69 = n67 & ~n68 ;
  assign n70 = ~x11 & ~n69 ;
  assign n71 = x4 & x5 ;
  assign n72 = n71 ^ x3 ;
  assign n73 = x9 & ~n40 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = n74 ^ n71 ;
  assign n76 = n75 ^ n74 ;
  assign n77 = ~x4 & ~x5 ;
  assign n78 = n56 & n77 ;
  assign n79 = ~x13 & ~x14 ;
  assign n80 = ~x10 & n79 ;
  assign n81 = n78 & n80 ;
  assign n82 = n81 ^ n74 ;
  assign n83 = n82 ^ n72 ;
  assign n84 = n76 & ~n83 ;
  assign n85 = n84 ^ n81 ;
  assign n86 = x7 & n32 ;
  assign n87 = ~n81 & ~n86 ;
  assign n88 = n87 ^ n72 ;
  assign n89 = ~n85 & ~n88 ;
  assign n90 = n89 ^ n87 ;
  assign n91 = ~n72 & n90 ;
  assign n92 = n91 ^ n84 ;
  assign n93 = n92 ^ x3 ;
  assign n94 = n93 ^ n81 ;
  assign n95 = x6 & ~n94 ;
  assign n96 = n70 & ~n95 ;
  assign n97 = ~n66 & n96 ;
  assign n98 = x3 & x8 ;
  assign n99 = ~x0 & x10 ;
  assign n100 = n98 & n99 ;
  assign n101 = x4 & n100 ;
  assign n102 = ~x13 & n19 ;
  assign n103 = n101 & n102 ;
  assign n104 = x9 & ~x10 ;
  assign n105 = x0 & n104 ;
  assign n106 = ~x1 & n105 ;
  assign n107 = ~n103 & ~n106 ;
  assign n108 = x14 & ~n107 ;
  assign n109 = ~x7 & n77 ;
  assign n110 = n21 & n99 ;
  assign n111 = x9 & n110 ;
  assign n112 = n109 & n111 ;
  assign n113 = n112 ^ x3 ;
  assign n114 = n113 ^ x11 ;
  assign n115 = n67 ^ x6 ;
  assign n116 = x3 & ~n115 ;
  assign n117 = n116 ^ n67 ;
  assign n118 = ~n114 & ~n117 ;
  assign n119 = n118 ^ n116 ;
  assign n120 = n119 ^ n67 ;
  assign n121 = n120 ^ x3 ;
  assign n122 = x11 & ~n121 ;
  assign n123 = ~n108 & n122 ;
  assign n124 = ~n97 & ~n123 ;
  assign n125 = x13 & n104 ;
  assign n126 = ~x0 & n125 ;
  assign n127 = x13 & x14 ;
  assign n128 = ~x5 & x14 ;
  assign n129 = ~x13 & ~n128 ;
  assign n130 = ~n127 & ~n129 ;
  assign n131 = n67 & n130 ;
  assign n132 = ~n126 & ~n131 ;
  assign n133 = ~x12 & n132 ;
  assign n134 = ~n124 & n133 ;
  assign n135 = ~x3 & x14 ;
  assign n136 = x11 & n135 ;
  assign n137 = x7 & ~x8 ;
  assign n138 = n137 ^ x6 ;
  assign n139 = n136 & ~n138 ;
  assign n140 = n104 & ~n139 ;
  assign n141 = ~x13 & n140 ;
  assign n142 = x14 & n38 ;
  assign n143 = n142 ^ n100 ;
  assign n144 = n143 ^ n142 ;
  assign n145 = ~x14 & n18 ;
  assign n146 = ~x2 & x5 ;
  assign n147 = ~x13 & n146 ;
  assign n148 = ~n20 & n147 ;
  assign n149 = ~n145 & ~n148 ;
  assign n150 = n149 ^ n142 ;
  assign n151 = n150 ^ n142 ;
  assign n152 = n144 & ~n151 ;
  assign n153 = n152 ^ n142 ;
  assign n154 = x4 & n153 ;
  assign n155 = n154 ^ n142 ;
  assign n156 = n155 ^ x11 ;
  assign n157 = n156 ^ n155 ;
  assign n158 = x4 & ~x10 ;
  assign n159 = ~x6 & x13 ;
  assign n160 = n109 & n159 ;
  assign n161 = n98 & n160 ;
  assign n162 = ~n158 & ~n161 ;
  assign n163 = x14 & ~n162 ;
  assign n164 = n163 ^ n155 ;
  assign n165 = ~n157 & n164 ;
  assign n166 = n165 ^ n155 ;
  assign n167 = ~x9 & n166 ;
  assign n168 = x12 & ~n167 ;
  assign n169 = ~n141 & n168 ;
  assign n170 = ~n134 & ~n169 ;
  assign n171 = x11 ^ x9 ;
  assign n172 = n171 ^ x10 ;
  assign n173 = x13 ^ x11 ;
  assign n174 = n173 ^ x13 ;
  assign n175 = n127 ^ x14 ;
  assign n176 = x3 & ~n175 ;
  assign n177 = n176 ^ x14 ;
  assign n178 = n177 ^ x13 ;
  assign n179 = ~n174 & ~n178 ;
  assign n180 = n179 ^ x13 ;
  assign n181 = n180 ^ n171 ;
  assign n182 = n172 & ~n181 ;
  assign n183 = n182 ^ n179 ;
  assign n184 = n183 ^ x13 ;
  assign n185 = n184 ^ x10 ;
  assign n186 = ~n171 & ~n185 ;
  assign n187 = n186 ^ n171 ;
  assign n188 = ~n170 & n187 ;
  assign y0 = ~n188 ;
endmodule
