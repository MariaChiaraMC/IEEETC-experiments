module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 ;
  assign n135 = x9 & x12 ;
  assign n93 = ~x4 & ~x5 ;
  assign n116 = x6 & n93 ;
  assign n37 = ~x11 & ~x14 ;
  assign n115 = ~x7 & ~x8 ;
  assign n136 = n37 & ~n115 ;
  assign n137 = n116 & n136 ;
  assign n138 = ~n135 & ~n137 ;
  assign n139 = ~x6 & x11 ;
  assign n140 = ~n138 & n139 ;
  assign n141 = x8 ^ x7 ;
  assign n142 = n141 ^ n139 ;
  assign n19 = x5 & ~x7 ;
  assign n143 = n140 ^ n19 ;
  assign n144 = n142 & n143 ;
  assign n145 = n144 ^ n19 ;
  assign n146 = n140 & n145 ;
  assign n147 = n146 ^ n138 ;
  assign n148 = ~x13 & ~n147 ;
  assign n128 = ~x9 & ~x11 ;
  assign n149 = x9 & ~x13 ;
  assign n150 = x12 & n149 ;
  assign n151 = ~n128 & ~n150 ;
  assign n152 = ~x3 & x14 ;
  assign n153 = ~n151 & ~n152 ;
  assign n70 = x4 & ~x9 ;
  assign n154 = ~x11 & n70 ;
  assign n155 = x7 & n37 ;
  assign n156 = ~n154 & ~n155 ;
  assign n157 = ~x10 & n156 ;
  assign n158 = x12 & ~n157 ;
  assign n159 = x11 & x13 ;
  assign n160 = ~x7 & x8 ;
  assign n161 = x6 & n160 ;
  assign n162 = ~n159 & ~n161 ;
  assign n163 = n135 & ~n162 ;
  assign n164 = ~n158 & ~n163 ;
  assign n165 = ~n153 & n164 ;
  assign n166 = ~n148 & n165 ;
  assign n16 = ~x5 & x7 ;
  assign n17 = x13 & n16 ;
  assign n18 = x9 & n17 ;
  assign n20 = x10 & ~n19 ;
  assign n21 = x9 ^ x3 ;
  assign n22 = n21 ^ x13 ;
  assign n23 = x13 ^ x9 ;
  assign n24 = x14 ^ x9 ;
  assign n25 = ~n23 & n24 ;
  assign n26 = n25 ^ x9 ;
  assign n27 = ~n22 & n26 ;
  assign n28 = n27 ^ x3 ;
  assign n29 = n20 & ~n28 ;
  assign n30 = x9 & x10 ;
  assign n31 = ~x14 & n30 ;
  assign n32 = ~n29 & ~n31 ;
  assign n33 = ~n18 & n32 ;
  assign n34 = x4 & ~x11 ;
  assign n35 = ~n33 & n34 ;
  assign n36 = ~x5 & n30 ;
  assign n38 = n37 ^ x6 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = x13 ^ x8 ;
  assign n41 = n40 ^ n37 ;
  assign n42 = n41 ^ n39 ;
  assign n43 = n39 & n42 ;
  assign n44 = n43 ^ n41 ;
  assign n45 = n44 ^ x13 ;
  assign n46 = n45 ^ n37 ;
  assign n48 = x7 ^ x6 ;
  assign n49 = n48 ^ n39 ;
  assign n47 = n39 ^ n37 ;
  assign n50 = n49 ^ n47 ;
  assign n51 = ~n37 & ~n50 ;
  assign n52 = n51 ^ n39 ;
  assign n53 = ~x4 & x11 ;
  assign n54 = ~x13 & n53 ;
  assign n55 = n54 ^ n37 ;
  assign n56 = n52 & ~n55 ;
  assign n57 = n56 ^ n49 ;
  assign n58 = n46 & n57 ;
  assign n59 = n58 ^ n51 ;
  assign n60 = n59 ^ n43 ;
  assign n61 = n60 ^ n41 ;
  assign n62 = n61 ^ x13 ;
  assign n63 = n62 ^ n49 ;
  assign n64 = n63 ^ n39 ;
  assign n65 = n36 & ~n64 ;
  assign n66 = ~x1 & ~x6 ;
  assign n67 = ~x11 & n66 ;
  assign n68 = x3 & ~x8 ;
  assign n69 = x5 & ~n68 ;
  assign n71 = ~x13 & x14 ;
  assign n72 = n70 & n71 ;
  assign n73 = n69 & n72 ;
  assign n74 = ~n67 & n73 ;
  assign n75 = ~n65 & ~n74 ;
  assign n76 = ~n35 & n75 ;
  assign n77 = ~x0 & ~n76 ;
  assign n78 = x1 & n16 ;
  assign n79 = x4 & n78 ;
  assign n80 = x3 & n79 ;
  assign n81 = ~x9 & x13 ;
  assign n82 = x4 & x5 ;
  assign n83 = x6 & n82 ;
  assign n84 = n30 & n83 ;
  assign n85 = ~n81 & ~n84 ;
  assign n86 = ~n80 & ~n85 ;
  assign n87 = n37 & n86 ;
  assign n88 = x7 & x10 ;
  assign n89 = n83 & n88 ;
  assign n90 = ~n28 & n89 ;
  assign n91 = n90 ^ x14 ;
  assign n92 = n91 ^ n90 ;
  assign n94 = ~x6 & n93 ;
  assign n95 = ~x9 & ~x13 ;
  assign n96 = x7 & x8 ;
  assign n97 = n95 & n96 ;
  assign n98 = n94 & n97 ;
  assign n99 = n98 ^ n90 ;
  assign n100 = n99 ^ n90 ;
  assign n101 = ~n92 & n100 ;
  assign n102 = n101 ^ n90 ;
  assign n103 = x11 & n102 ;
  assign n104 = n103 ^ n90 ;
  assign n105 = ~n87 & ~n104 ;
  assign n106 = x14 ^ x1 ;
  assign n107 = n106 ^ x1 ;
  assign n108 = x13 ^ x1 ;
  assign n109 = ~n107 & n108 ;
  assign n110 = n109 ^ x1 ;
  assign n111 = x0 & n110 ;
  assign n112 = x11 ^ x0 ;
  assign n113 = n112 ^ x11 ;
  assign n114 = n113 ^ n111 ;
  assign n117 = ~n115 & n116 ;
  assign n118 = ~x13 & ~n117 ;
  assign n119 = n118 ^ n71 ;
  assign n120 = x11 & n119 ;
  assign n121 = n120 ^ n118 ;
  assign n122 = n114 & ~n121 ;
  assign n123 = n122 ^ n120 ;
  assign n124 = n123 ^ n118 ;
  assign n125 = n124 ^ x11 ;
  assign n126 = ~n111 & ~n125 ;
  assign n127 = x9 & ~n126 ;
  assign n129 = x13 & n128 ;
  assign n130 = x1 & n129 ;
  assign n131 = ~x10 & ~n130 ;
  assign n132 = ~n127 & n131 ;
  assign n133 = n105 & ~n132 ;
  assign n134 = ~n77 & n133 ;
  assign n167 = n166 ^ n134 ;
  assign n168 = n167 ^ x12 ;
  assign n175 = n168 ^ n167 ;
  assign n169 = n168 ^ x10 ;
  assign n170 = n169 ^ n167 ;
  assign n171 = n168 ^ n134 ;
  assign n172 = n171 ^ x10 ;
  assign n173 = n172 ^ n170 ;
  assign n174 = ~n170 & n173 ;
  assign n176 = n175 ^ n174 ;
  assign n177 = n176 ^ n170 ;
  assign n178 = ~x0 & x11 ;
  assign n179 = ~x3 & ~x14 ;
  assign n180 = x13 & n179 ;
  assign n181 = n79 & n180 ;
  assign n182 = ~x2 & ~x13 ;
  assign n183 = n69 & n182 ;
  assign n184 = ~n66 & n183 ;
  assign n185 = ~n181 & ~n184 ;
  assign n186 = n178 & ~n185 ;
  assign n187 = x7 & ~x8 ;
  assign n188 = x14 & n94 ;
  assign n189 = n187 & n188 ;
  assign n190 = ~n53 & ~n189 ;
  assign n191 = ~x13 & ~n190 ;
  assign n192 = ~n186 & ~n191 ;
  assign n193 = ~x9 & ~n192 ;
  assign n194 = x13 & n160 ;
  assign n195 = n188 & n194 ;
  assign n196 = ~x11 & n195 ;
  assign n197 = ~n193 & ~n196 ;
  assign n198 = n197 ^ n167 ;
  assign n199 = n174 ^ n170 ;
  assign n200 = n198 & ~n199 ;
  assign n201 = n200 ^ n167 ;
  assign n202 = n177 & n201 ;
  assign n203 = n202 ^ n167 ;
  assign n204 = n203 ^ n166 ;
  assign n205 = n204 ^ n167 ;
  assign y0 = ~n205 ;
endmodule
