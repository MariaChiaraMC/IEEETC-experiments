module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 ;
  assign n69 = x5 & x7 ;
  assign n70 = ~x2 & n69 ;
  assign n71 = ~x0 & ~n70 ;
  assign n72 = ~x3 & ~n71 ;
  assign n17 = x3 & ~x6 ;
  assign n18 = x9 ^ x8 ;
  assign n19 = n18 ^ x10 ;
  assign n20 = x10 ^ x9 ;
  assign n21 = x10 ^ x5 ;
  assign n22 = x10 & ~n21 ;
  assign n23 = n22 ^ x10 ;
  assign n24 = n20 & n23 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = n25 ^ x10 ;
  assign n27 = n26 ^ x5 ;
  assign n28 = n19 & ~n27 ;
  assign n29 = n28 ^ x5 ;
  assign n30 = n17 & n29 ;
  assign n31 = n30 ^ x3 ;
  assign n32 = n31 ^ x7 ;
  assign n58 = n32 ^ n31 ;
  assign n33 = x15 ^ x14 ;
  assign n34 = n33 ^ x13 ;
  assign n35 = x15 ^ x13 ;
  assign n36 = x9 & x10 ;
  assign n37 = x6 & ~n36 ;
  assign n38 = x7 & ~n37 ;
  assign n39 = ~x9 & ~x10 ;
  assign n40 = ~x8 & ~n39 ;
  assign n41 = ~x11 & ~x12 ;
  assign n42 = n40 & n41 ;
  assign n43 = ~n38 & n42 ;
  assign n44 = n43 ^ x13 ;
  assign n45 = x13 & n44 ;
  assign n46 = n45 ^ x13 ;
  assign n47 = n35 & n46 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = n48 ^ x13 ;
  assign n50 = n49 ^ n43 ;
  assign n51 = n34 & n50 ;
  assign n52 = n51 ^ n32 ;
  assign n53 = n52 ^ n31 ;
  assign n54 = n32 ^ n30 ;
  assign n55 = n54 ^ n51 ;
  assign n56 = n55 ^ n53 ;
  assign n57 = n53 & n56 ;
  assign n59 = n58 ^ n57 ;
  assign n60 = n59 ^ n53 ;
  assign n61 = n31 ^ x5 ;
  assign n62 = n57 ^ n53 ;
  assign n63 = ~n61 & n62 ;
  assign n64 = n63 ^ n31 ;
  assign n65 = ~n60 & ~n64 ;
  assign n66 = n65 ^ n31 ;
  assign n67 = n66 ^ x3 ;
  assign n68 = n67 ^ n31 ;
  assign n73 = n72 ^ n68 ;
  assign n74 = n73 ^ n72 ;
  assign n75 = ~x0 & ~x2 ;
  assign n76 = n75 ^ n72 ;
  assign n77 = n76 ^ n72 ;
  assign n78 = ~n74 & n77 ;
  assign n79 = n78 ^ n72 ;
  assign n80 = x1 & n79 ;
  assign n81 = n80 ^ n72 ;
  assign n82 = x4 & n81 ;
  assign y0 = n82 ;
endmodule
