module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 ;
  assign n11 = ~x6 & ~x8 ;
  assign n10 = x5 ^ x4 ;
  assign n12 = n11 ^ n10 ;
  assign n13 = n12 ^ x5 ;
  assign n14 = n11 ^ x7 ;
  assign n15 = n14 ^ x7 ;
  assign n16 = x0 & x3 ;
  assign n17 = ~x1 & x2 ;
  assign n18 = n16 & n17 ;
  assign n19 = ~x7 & n18 ;
  assign n20 = n19 ^ x7 ;
  assign n21 = n15 & n20 ;
  assign n22 = n21 ^ x7 ;
  assign n23 = n22 ^ n12 ;
  assign n24 = ~n13 & n23 ;
  assign n25 = n24 ^ n21 ;
  assign n26 = n25 ^ x7 ;
  assign n27 = n26 ^ x5 ;
  assign n28 = n12 & ~n27 ;
  assign n29 = n28 ^ n12 ;
  assign n30 = n29 ^ n10 ;
  assign y0 = n30 ;
endmodule
