module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n13 = x8 & x9 ;
  assign n14 = x5 & ~x11 ;
  assign n15 = ~x1 & n14 ;
  assign n16 = x0 & n15 ;
  assign n17 = n16 ^ n13 ;
  assign n20 = x2 & x4 ;
  assign n21 = x3 & n20 ;
  assign n18 = x7 & x10 ;
  assign n19 = x6 & n18 ;
  assign n22 = n21 ^ n19 ;
  assign n23 = n22 ^ n19 ;
  assign n24 = ~x6 & ~x7 ;
  assign n25 = n24 ^ n19 ;
  assign n26 = ~n23 & n25 ;
  assign n27 = n26 ^ n19 ;
  assign n28 = n27 ^ n13 ;
  assign n29 = n17 & n28 ;
  assign n30 = n29 ^ n26 ;
  assign n31 = n30 ^ n19 ;
  assign n32 = n31 ^ n16 ;
  assign n33 = n13 & n32 ;
  assign n34 = n33 ^ n13 ;
  assign y0 = n34 ;
endmodule
