module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 ;
  assign n15 = x6 ^ x1 ;
  assign n13 = x7 ^ x6 ;
  assign n12 = x6 ^ x4 ;
  assign n14 = n13 ^ n12 ;
  assign n16 = n15 ^ n14 ;
  assign n10 = x6 ^ x3 ;
  assign n17 = n16 ^ n10 ;
  assign n18 = n17 ^ x6 ;
  assign n20 = n18 ^ n13 ;
  assign n21 = n20 ^ n15 ;
  assign n22 = n21 ^ n10 ;
  assign n23 = n22 ^ x6 ;
  assign n11 = n10 ^ x6 ;
  assign n19 = n18 ^ n11 ;
  assign n24 = n23 ^ n19 ;
  assign n28 = x8 ^ x6 ;
  assign n29 = n28 ^ n15 ;
  assign n25 = n15 ^ n10 ;
  assign n26 = n25 ^ x6 ;
  assign n27 = n26 ^ x6 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n30 ^ n18 ;
  assign n32 = ~n11 & n31 ;
  assign n33 = n32 ^ n26 ;
  assign n34 = n24 & n33 ;
  assign n35 = n34 ^ n26 ;
  assign n36 = n35 ^ n29 ;
  assign n37 = n36 ^ n18 ;
  assign n38 = n33 ^ n29 ;
  assign n39 = n38 ^ n18 ;
  assign n40 = ~n23 & n39 ;
  assign n41 = n40 ^ n11 ;
  assign n42 = n37 & ~n41 ;
  assign n43 = n42 ^ n32 ;
  assign n44 = n43 ^ n34 ;
  assign n45 = n44 ^ n40 ;
  assign n46 = n45 ^ n26 ;
  assign n47 = n46 ^ x6 ;
  assign n48 = n47 ^ n26 ;
  assign n49 = x2 & n48 ;
  assign n50 = x4 ^ x3 ;
  assign n51 = ~x7 & ~x8 ;
  assign n52 = n51 ^ x4 ;
  assign n53 = n52 ^ n51 ;
  assign n54 = x7 & x8 ;
  assign n55 = n54 ^ n51 ;
  assign n56 = n53 & n55 ;
  assign n57 = n56 ^ n51 ;
  assign n58 = n50 & n57 ;
  assign n59 = n58 ^ x3 ;
  assign n60 = ~x2 & ~n59 ;
  assign n61 = x6 & ~n60 ;
  assign n62 = x1 & ~n61 ;
  assign n63 = x2 & x7 ;
  assign n64 = n63 ^ x3 ;
  assign n65 = ~x4 & ~x8 ;
  assign n66 = n65 ^ n63 ;
  assign n67 = n66 ^ n65 ;
  assign n68 = n67 ^ n64 ;
  assign n69 = x2 & x8 ;
  assign n70 = n69 ^ x4 ;
  assign n71 = x4 & n70 ;
  assign n72 = n71 ^ n65 ;
  assign n73 = n72 ^ x4 ;
  assign n74 = ~n68 & n73 ;
  assign n75 = n74 ^ n71 ;
  assign n76 = n75 ^ x4 ;
  assign n77 = n64 & n76 ;
  assign n78 = n77 ^ n63 ;
  assign n79 = n62 & ~n78 ;
  assign n80 = ~n49 & ~n79 ;
  assign n83 = n80 ^ x1 ;
  assign n84 = n83 ^ n80 ;
  assign n81 = n80 ^ x6 ;
  assign n82 = n81 ^ n80 ;
  assign n85 = n84 ^ n82 ;
  assign n86 = x3 & x4 ;
  assign n87 = n63 & ~n86 ;
  assign n88 = x3 & ~n65 ;
  assign n89 = x7 & n88 ;
  assign n90 = n89 ^ n69 ;
  assign n91 = n90 ^ n89 ;
  assign n92 = ~x3 & ~x4 ;
  assign n93 = n92 ^ n89 ;
  assign n94 = n91 & ~n93 ;
  assign n95 = n94 ^ n89 ;
  assign n96 = ~n87 & ~n95 ;
  assign n97 = n96 ^ n80 ;
  assign n98 = n97 ^ n80 ;
  assign n99 = n98 ^ n84 ;
  assign n100 = n84 & ~n99 ;
  assign n101 = n100 ^ n84 ;
  assign n102 = n85 & n101 ;
  assign n103 = n102 ^ n100 ;
  assign n104 = n103 ^ n80 ;
  assign n105 = n104 ^ n84 ;
  assign n106 = ~x5 & ~n105 ;
  assign n107 = n106 ^ n80 ;
  assign n108 = x0 & ~n107 ;
  assign y0 = n108 ;
endmodule
