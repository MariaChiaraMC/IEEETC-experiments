module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 ;
  assign n15 = ~x0 & x3 ;
  assign n16 = x1 & x6 ;
  assign n21 = x5 & ~x11 ;
  assign n22 = ~x10 & ~x12 ;
  assign n23 = x4 & ~x13 ;
  assign n24 = n22 & n23 ;
  assign n25 = n21 & n24 ;
  assign n17 = ~x2 & ~x4 ;
  assign n18 = ~x5 & n17 ;
  assign n26 = n25 ^ n18 ;
  assign n27 = n26 ^ n18 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = n19 ^ n18 ;
  assign n28 = n27 ^ n20 ;
  assign n29 = x7 & ~x8 ;
  assign n30 = ~x9 & n29 ;
  assign n31 = n30 ^ n18 ;
  assign n32 = n31 ^ n18 ;
  assign n33 = n32 ^ n27 ;
  assign n34 = n27 & n33 ;
  assign n35 = n34 ^ n27 ;
  assign n36 = n28 & n35 ;
  assign n37 = n36 ^ n34 ;
  assign n38 = n37 ^ n18 ;
  assign n39 = n38 ^ n27 ;
  assign n40 = n16 & n39 ;
  assign n41 = n40 ^ n18 ;
  assign n42 = n15 & n41 ;
  assign y0 = n42 ;
endmodule
