module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 ;
  assign n8 = x5 ^ x2 ;
  assign n9 = n8 ^ x1 ;
  assign n10 = n9 ^ x0 ;
  assign n11 = ~x3 & ~x4 ;
  assign n12 = ~x2 & ~n11 ;
  assign n13 = ~x6 & ~n12 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = n14 ^ n9 ;
  assign n16 = x1 & n15 ;
  assign n17 = n16 ^ x5 ;
  assign n18 = n17 ^ x1 ;
  assign n19 = n18 ^ n9 ;
  assign n20 = n19 ^ x0 ;
  assign n21 = ~n10 & ~n20 ;
  assign n22 = n21 ^ n16 ;
  assign n23 = n22 ^ x5 ;
  assign n24 = n23 ^ n9 ;
  assign n25 = ~x0 & n24 ;
  assign n26 = n25 ^ x0 ;
  assign n27 = n26 ^ x0 ;
  assign n28 = x3 & x4 ;
  assign n29 = n28 ^ x1 ;
  assign n30 = x6 ^ x2 ;
  assign n31 = n28 ^ x2 ;
  assign n32 = n31 ^ x2 ;
  assign n33 = n30 & n32 ;
  assign n34 = n33 ^ x2 ;
  assign n35 = n29 & n34 ;
  assign n36 = n35 ^ x1 ;
  assign n37 = n27 & n36 ;
  assign y0 = n37 ;
endmodule
