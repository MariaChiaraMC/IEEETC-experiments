module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 ;
  assign n7 = x1 & ~x5 ;
  assign n8 = x0 & x4 ;
  assign n9 = n7 & n8 ;
  assign n10 = ~x3 & n9 ;
  assign n11 = x3 ^ x0 ;
  assign n12 = n11 ^ x1 ;
  assign n13 = n12 ^ x0 ;
  assign n14 = n13 ^ x5 ;
  assign n15 = x4 ^ x1 ;
  assign n16 = ~x4 & n15 ;
  assign n17 = n16 ^ x0 ;
  assign n18 = n17 ^ x4 ;
  assign n19 = ~n14 & n18 ;
  assign n20 = n19 ^ n16 ;
  assign n21 = n20 ^ x4 ;
  assign n22 = x5 & ~n21 ;
  assign n23 = ~n10 & ~n22 ;
  assign n24 = ~x0 & ~x4 ;
  assign n25 = x3 & ~n7 ;
  assign n26 = n24 & ~n25 ;
  assign n27 = ~x2 & ~n26 ;
  assign n28 = n23 & n27 ;
  assign n29 = x4 ^ x0 ;
  assign n30 = n29 ^ x1 ;
  assign n31 = n30 ^ n29 ;
  assign n32 = n29 ^ x4 ;
  assign n33 = n32 ^ n29 ;
  assign n34 = n31 & n33 ;
  assign n35 = n34 ^ n29 ;
  assign n36 = ~x5 & ~n35 ;
  assign n37 = n36 ^ n29 ;
  assign n38 = x3 & ~n37 ;
  assign n39 = x2 & ~n38 ;
  assign n40 = x0 & x5 ;
  assign n41 = ~n24 & ~n40 ;
  assign n42 = n41 ^ x3 ;
  assign n43 = n41 ^ n8 ;
  assign n44 = n41 ^ x1 ;
  assign n45 = n41 & ~n44 ;
  assign n46 = n45 ^ n41 ;
  assign n47 = n43 & n46 ;
  assign n48 = n47 ^ n45 ;
  assign n49 = n48 ^ n41 ;
  assign n50 = n49 ^ x1 ;
  assign n51 = n42 & ~n50 ;
  assign n52 = n39 & ~n51 ;
  assign n53 = ~n28 & ~n52 ;
  assign y0 = n53 ;
endmodule
