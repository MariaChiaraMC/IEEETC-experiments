module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 ;
  output y0 ;
  wire n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 ;
  assign n14 = x8 ^ x7 ;
  assign n15 = n14 ^ x7 ;
  assign n16 = x11 & x12 ;
  assign n17 = ~x9 & ~n16 ;
  assign n18 = n17 ^ x10 ;
  assign n19 = x4 & x5 ;
  assign n20 = x3 & x6 ;
  assign n21 = x2 & ~n20 ;
  assign n22 = ~n19 & n21 ;
  assign n23 = x1 & ~n22 ;
  assign n24 = ~x12 & ~n23 ;
  assign n25 = ~x11 & n24 ;
  assign n26 = n25 ^ n17 ;
  assign n27 = x10 ^ x7 ;
  assign n28 = n27 ^ n25 ;
  assign n29 = n25 & ~n28 ;
  assign n30 = n29 ^ n25 ;
  assign n31 = n26 & n30 ;
  assign n32 = n31 ^ n29 ;
  assign n33 = n32 ^ n25 ;
  assign n34 = n33 ^ n27 ;
  assign n35 = n18 & ~n34 ;
  assign n36 = n35 ^ x7 ;
  assign n37 = n36 ^ x7 ;
  assign n38 = ~n15 & ~n37 ;
  assign n39 = n38 ^ x7 ;
  assign n40 = ~x0 & ~n39 ;
  assign y0 = n40 ;
endmodule
