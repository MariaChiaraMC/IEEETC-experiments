module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 ;
  assign n8 = x5 ^ x0 ;
  assign n9 = x5 ^ x1 ;
  assign n10 = x6 ^ x1 ;
  assign n11 = n10 ^ x1 ;
  assign n12 = n9 & n11 ;
  assign n13 = n12 ^ x1 ;
  assign n14 = ~n8 & n13 ;
  assign n15 = n14 ^ x0 ;
  assign n16 = x4 & ~n15 ;
  assign n17 = ~x4 & ~x6 ;
  assign n18 = ~x5 & n17 ;
  assign n19 = ~x3 & ~n18 ;
  assign n20 = ~x2 & n19 ;
  assign n21 = ~n16 & n20 ;
  assign y0 = n21 ;
endmodule
