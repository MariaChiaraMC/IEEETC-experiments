module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 ;
  assign n9 = x2 & ~x4 ;
  assign n18 = n9 ^ x3 ;
  assign n19 = n9 ^ x7 ;
  assign n20 = n19 ^ x7 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = x5 ^ x4 ;
  assign n23 = x4 & n22 ;
  assign n24 = n23 ^ x7 ;
  assign n25 = n24 ^ x4 ;
  assign n26 = n21 & n25 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = n27 ^ x4 ;
  assign n29 = ~n18 & n28 ;
  assign n30 = n29 ^ n9 ;
  assign n10 = n9 ^ x5 ;
  assign n11 = x4 ^ x3 ;
  assign n12 = n9 ^ x4 ;
  assign n13 = n12 ^ x4 ;
  assign n14 = n11 & n13 ;
  assign n15 = n14 ^ x4 ;
  assign n16 = n10 & n15 ;
  assign n17 = n16 ^ x5 ;
  assign n31 = n30 ^ n17 ;
  assign n32 = ~x6 & n31 ;
  assign n33 = n32 ^ n30 ;
  assign n34 = ~x1 & n33 ;
  assign n41 = x4 ^ x1 ;
  assign n42 = ~x3 & ~x5 ;
  assign n43 = n42 ^ x4 ;
  assign n44 = n43 ^ n42 ;
  assign n36 = x3 & ~x5 ;
  assign n37 = x6 & n36 ;
  assign n45 = n42 ^ n37 ;
  assign n46 = n44 & n45 ;
  assign n47 = n46 ^ n42 ;
  assign n48 = n41 & n47 ;
  assign n49 = n48 ^ x1 ;
  assign n50 = x5 ^ x3 ;
  assign n51 = ~x1 & ~x7 ;
  assign n52 = n51 ^ x3 ;
  assign n53 = n51 ^ x6 ;
  assign n54 = ~n51 & n53 ;
  assign n55 = n54 ^ n51 ;
  assign n56 = n52 & ~n55 ;
  assign n57 = n56 ^ n54 ;
  assign n58 = n57 ^ n51 ;
  assign n59 = n58 ^ x6 ;
  assign n60 = ~n50 & n59 ;
  assign n61 = ~n49 & ~n60 ;
  assign n38 = ~x1 & ~x4 ;
  assign n39 = n37 & n38 ;
  assign n35 = x7 ^ x2 ;
  assign n40 = n39 ^ n35 ;
  assign n62 = n61 ^ n40 ;
  assign n63 = n62 ^ n35 ;
  assign n64 = n40 ^ x7 ;
  assign n65 = n64 ^ n40 ;
  assign n66 = n65 ^ n63 ;
  assign n67 = n63 & n66 ;
  assign n68 = n67 ^ n61 ;
  assign n69 = n68 ^ n63 ;
  assign n70 = n61 ^ x6 ;
  assign n71 = n70 ^ n35 ;
  assign n72 = ~x6 & ~n71 ;
  assign n73 = n72 ^ x6 ;
  assign n74 = n73 ^ n61 ;
  assign n75 = ~x3 & x4 ;
  assign n76 = n75 ^ x6 ;
  assign n77 = ~n70 & ~n76 ;
  assign n78 = n77 ^ n75 ;
  assign n79 = n78 ^ n35 ;
  assign n80 = ~n74 & n79 ;
  assign n81 = n80 ^ n35 ;
  assign n82 = n69 & n81 ;
  assign n83 = n82 ^ n67 ;
  assign n84 = n83 ^ n80 ;
  assign n85 = n84 ^ n63 ;
  assign n86 = n85 ^ x2 ;
  assign n87 = n86 ^ n61 ;
  assign n88 = ~n34 & n87 ;
  assign n89 = ~x0 & ~n88 ;
  assign y0 = n89 ;
endmodule
