module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 ;
  assign n16 = ~x10 & ~x14 ;
  assign n17 = ~x0 & ~x6 ;
  assign n18 = ~x1 & n17 ;
  assign n19 = ~x2 & n18 ;
  assign n20 = x13 ^ x7 ;
  assign n21 = x7 ^ x5 ;
  assign n22 = n21 ^ n20 ;
  assign n23 = x13 ^ x8 ;
  assign n24 = n23 ^ x8 ;
  assign n25 = ~x8 & ~x9 ;
  assign n26 = n25 ^ x8 ;
  assign n27 = n24 & n26 ;
  assign n28 = n27 ^ x8 ;
  assign n29 = n28 ^ n20 ;
  assign n30 = ~n22 & n29 ;
  assign n31 = n30 ^ n27 ;
  assign n32 = n31 ^ x8 ;
  assign n33 = n32 ^ n21 ;
  assign n34 = n20 & ~n33 ;
  assign n35 = n34 ^ n20 ;
  assign n36 = n19 & n35 ;
  assign n37 = x0 & x6 ;
  assign n38 = x1 & n37 ;
  assign n39 = x7 & ~x13 ;
  assign n40 = n39 ^ n38 ;
  assign n41 = x8 & x9 ;
  assign n42 = x2 & n41 ;
  assign n43 = n42 ^ x5 ;
  assign n44 = n43 ^ n42 ;
  assign n45 = n42 ^ x9 ;
  assign n46 = ~n44 & ~n45 ;
  assign n47 = n46 ^ n42 ;
  assign n48 = n47 ^ n38 ;
  assign n49 = n40 & n48 ;
  assign n50 = n49 ^ n46 ;
  assign n51 = n50 ^ n42 ;
  assign n52 = n51 ^ n39 ;
  assign n53 = n38 & n52 ;
  assign n54 = n53 ^ n38 ;
  assign n55 = ~n36 & ~n54 ;
  assign n56 = ~x3 & ~n55 ;
  assign n57 = ~x5 & n38 ;
  assign n58 = ~x2 & x3 ;
  assign n59 = n58 ^ x13 ;
  assign n60 = x2 & x7 ;
  assign n61 = n60 ^ n41 ;
  assign n62 = n61 ^ n41 ;
  assign n63 = n41 ^ x9 ;
  assign n64 = n62 & ~n63 ;
  assign n65 = n64 ^ n41 ;
  assign n66 = n65 ^ n58 ;
  assign n67 = n59 & ~n66 ;
  assign n68 = n67 ^ n64 ;
  assign n69 = n68 ^ n41 ;
  assign n70 = n69 ^ x13 ;
  assign n71 = ~n58 & ~n70 ;
  assign n72 = n71 ^ n58 ;
  assign n73 = n57 & ~n72 ;
  assign n74 = ~n56 & ~n73 ;
  assign n75 = n74 ^ x4 ;
  assign n76 = n75 ^ n74 ;
  assign n77 = ~x5 & n39 ;
  assign n78 = x2 & x6 ;
  assign n79 = x0 & n78 ;
  assign n80 = n77 & n79 ;
  assign n81 = ~x1 & x3 ;
  assign n82 = x9 ^ x8 ;
  assign n83 = n81 & ~n82 ;
  assign n84 = n80 & n83 ;
  assign n85 = n84 ^ n74 ;
  assign n86 = n76 & ~n85 ;
  assign n87 = n86 ^ n74 ;
  assign n88 = n16 & ~n87 ;
  assign n89 = x2 & x10 ;
  assign n90 = ~x8 & n18 ;
  assign n91 = n89 & n90 ;
  assign n92 = ~x4 & n77 ;
  assign n93 = n92 ^ x3 ;
  assign n94 = n93 ^ n92 ;
  assign n95 = x5 & x13 ;
  assign n96 = x4 & x14 ;
  assign n97 = n95 & n96 ;
  assign n98 = x9 & n97 ;
  assign n99 = n98 ^ n92 ;
  assign n100 = ~n94 & n99 ;
  assign n101 = n100 ^ n92 ;
  assign n102 = n91 & n101 ;
  assign n103 = ~n88 & ~n102 ;
  assign n104 = ~x11 & ~x12 ;
  assign n105 = ~n103 & n104 ;
  assign y0 = n105 ;
endmodule
