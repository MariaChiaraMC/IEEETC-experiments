module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 ;
  assign n9 = x4 ^ x1 ;
  assign n10 = n9 ^ x3 ;
  assign n11 = n10 ^ x4 ;
  assign n14 = n11 ^ x4 ;
  assign n12 = n11 ^ x5 ;
  assign n15 = n14 ^ n12 ;
  assign n16 = n15 ^ n12 ;
  assign n17 = n16 ^ n11 ;
  assign n18 = n17 ^ n9 ;
  assign n13 = n12 ^ n11 ;
  assign n19 = n18 ^ n13 ;
  assign n20 = n11 ^ n9 ;
  assign n21 = n20 ^ n13 ;
  assign n22 = n21 ^ n18 ;
  assign n23 = n19 & n22 ;
  assign n24 = n23 ^ n11 ;
  assign n25 = n24 ^ n13 ;
  assign n26 = n25 ^ n18 ;
  assign n27 = n9 ^ x2 ;
  assign n28 = n27 ^ n11 ;
  assign n29 = ~x2 & ~x6 ;
  assign n30 = ~x7 & n29 ;
  assign n31 = n30 ^ n9 ;
  assign n32 = n31 ^ x2 ;
  assign n33 = n32 ^ n11 ;
  assign n34 = ~n28 & ~n33 ;
  assign n35 = n34 ^ n31 ;
  assign n36 = n35 ^ x2 ;
  assign n37 = n36 ^ n11 ;
  assign n38 = n37 ^ n18 ;
  assign n39 = n33 ^ n13 ;
  assign n40 = n32 ^ n9 ;
  assign n41 = n40 ^ n11 ;
  assign n42 = n41 ^ n13 ;
  assign n43 = n42 ^ n18 ;
  assign n44 = n39 & ~n43 ;
  assign n45 = n44 ^ n31 ;
  assign n46 = n45 ^ n18 ;
  assign n47 = n38 & ~n46 ;
  assign n48 = n47 ^ n11 ;
  assign n49 = n48 ^ n13 ;
  assign n50 = n26 & ~n49 ;
  assign n51 = n50 ^ n23 ;
  assign n52 = n51 ^ n11 ;
  assign n53 = n52 ^ n13 ;
  assign n54 = n53 ^ n18 ;
  assign n55 = n54 ^ x1 ;
  assign n56 = ~x0 & ~n55 ;
  assign n57 = ~x1 & x7 ;
  assign n58 = ~x6 & ~n57 ;
  assign n59 = ~x5 & ~n58 ;
  assign n60 = x6 ^ x2 ;
  assign n61 = ~n59 & ~n60 ;
  assign n62 = ~x4 & ~n61 ;
  assign n63 = ~x3 & n62 ;
  assign n64 = n56 & ~n63 ;
  assign y0 = n64 ;
endmodule
