module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n13 = x3 ^ x2 ;
  assign n14 = n13 ^ x2 ;
  assign n15 = x4 ^ x2 ;
  assign n16 = ~n14 & ~n15 ;
  assign n17 = n16 ^ x2 ;
  assign n18 = ~x2 & x10 ;
  assign n19 = n18 ^ x7 ;
  assign n20 = ~n17 & n19 ;
  assign n21 = n20 ^ n18 ;
  assign n22 = x7 & n21 ;
  assign n23 = n22 ^ x7 ;
  assign n24 = n23 ^ x9 ;
  assign n25 = n23 ^ x4 ;
  assign n26 = n25 ^ x4 ;
  assign n27 = x4 & ~x7 ;
  assign n28 = x2 & x3 ;
  assign n29 = n27 & ~n28 ;
  assign n30 = n29 ^ x4 ;
  assign n31 = ~n26 & ~n30 ;
  assign n32 = n31 ^ x4 ;
  assign n33 = n24 & n32 ;
  assign n34 = n33 ^ x9 ;
  assign y0 = n34 ;
endmodule
