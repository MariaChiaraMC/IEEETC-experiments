module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 ;
  output y0 ;
  wire n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 ;
  assign n24 = ~x3 & ~x4 ;
  assign n25 = x1 ^ x0 ;
  assign n26 = n25 ^ x5 ;
  assign n27 = n24 & n26 ;
  assign n28 = n27 ^ n24 ;
  assign n29 = x2 ^ x0 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n25 & ~n30 ;
  assign n32 = n31 ^ n25 ;
  assign n33 = n32 ^ x5 ;
  assign n34 = n28 & n33 ;
  assign n35 = x14 & ~n34 ;
  assign n36 = ~x18 & ~x19 ;
  assign n37 = x1 & x4 ;
  assign n38 = x2 & ~x3 ;
  assign n39 = n37 & n38 ;
  assign n40 = ~x6 & ~x7 ;
  assign n41 = ~x12 & n40 ;
  assign n42 = ~x11 & ~x13 ;
  assign n43 = n41 & n42 ;
  assign n44 = ~x8 & x10 ;
  assign n45 = ~x1 & x3 ;
  assign n46 = n44 & n45 ;
  assign n47 = ~x2 & ~x4 ;
  assign n48 = n46 & n47 ;
  assign n49 = n43 & n48 ;
  assign n50 = ~n39 & ~n49 ;
  assign n51 = ~x0 & ~n50 ;
  assign n52 = ~x3 & x4 ;
  assign n53 = ~x8 & x9 ;
  assign n54 = x11 & ~x12 ;
  assign n55 = x6 & x7 ;
  assign n56 = ~x15 & ~n55 ;
  assign n57 = n54 & ~n56 ;
  assign n58 = n53 & n57 ;
  assign n59 = ~x1 & ~n58 ;
  assign n60 = x8 & ~x10 ;
  assign n61 = x15 & n60 ;
  assign n62 = x10 ^ x8 ;
  assign n63 = ~x10 & x11 ;
  assign n64 = n63 ^ x9 ;
  assign n65 = n62 & ~n64 ;
  assign n66 = ~x13 & n65 ;
  assign n67 = ~n61 & ~n66 ;
  assign n68 = n41 & ~n67 ;
  assign n69 = ~x8 & ~x9 ;
  assign n70 = n63 & n69 ;
  assign n71 = n70 ^ x6 ;
  assign n72 = x13 & ~n71 ;
  assign n73 = n72 ^ x6 ;
  assign n74 = x12 & ~n73 ;
  assign n75 = x11 & n40 ;
  assign n76 = ~x13 & n69 ;
  assign n77 = ~x15 & ~n76 ;
  assign n78 = n75 & ~n77 ;
  assign n79 = ~n74 & ~n78 ;
  assign n80 = ~x16 & ~n79 ;
  assign n81 = x9 & x10 ;
  assign n82 = x8 & n42 ;
  assign n83 = ~x15 & ~n82 ;
  assign n84 = n81 & ~n83 ;
  assign n85 = ~x12 & n84 ;
  assign n86 = ~x12 & ~x13 ;
  assign n87 = ~n81 & n86 ;
  assign n88 = ~x11 & n86 ;
  assign n89 = x6 & ~n88 ;
  assign n90 = ~n87 & n89 ;
  assign n91 = n90 ^ x13 ;
  assign n92 = n91 ^ x17 ;
  assign n93 = x15 ^ x7 ;
  assign n94 = ~x13 & ~n93 ;
  assign n95 = n94 ^ x15 ;
  assign n96 = ~n92 & ~n95 ;
  assign n97 = n96 ^ n94 ;
  assign n98 = n97 ^ x15 ;
  assign n99 = n98 ^ x13 ;
  assign n100 = ~x17 & n99 ;
  assign n101 = ~n85 & n100 ;
  assign n102 = ~n80 & n101 ;
  assign n103 = ~n68 & n102 ;
  assign n104 = n103 ^ x2 ;
  assign n105 = n104 ^ n103 ;
  assign n106 = n60 ^ x13 ;
  assign n107 = n106 ^ x13 ;
  assign n110 = x13 ^ x12 ;
  assign n108 = x13 ^ x9 ;
  assign n109 = n108 ^ x13 ;
  assign n111 = n110 ^ n109 ;
  assign n112 = ~n107 & ~n111 ;
  assign n113 = n112 ^ n107 ;
  assign n114 = n113 ^ n110 ;
  assign n115 = x13 ^ x10 ;
  assign n116 = x13 ^ x11 ;
  assign n117 = n116 ^ n109 ;
  assign n118 = n115 & n117 ;
  assign n119 = n118 ^ x10 ;
  assign n120 = n119 ^ x13 ;
  assign n121 = n120 ^ n109 ;
  assign n122 = n121 ^ n116 ;
  assign n123 = n122 ^ n110 ;
  assign n124 = n109 ^ x13 ;
  assign n125 = ~n110 & n124 ;
  assign n126 = n125 ^ n109 ;
  assign n127 = n126 ^ n116 ;
  assign n128 = n127 ^ n110 ;
  assign n129 = ~n123 & ~n128 ;
  assign n130 = n129 ^ n116 ;
  assign n131 = n114 & n130 ;
  assign n132 = n131 ^ n125 ;
  assign n133 = n132 ^ n129 ;
  assign n134 = n133 ^ n109 ;
  assign n135 = n134 ^ n116 ;
  assign n136 = n135 ^ x12 ;
  assign n137 = n136 ^ n110 ;
  assign n138 = n137 ^ n103 ;
  assign n139 = ~n105 & ~n138 ;
  assign n140 = n139 ^ n103 ;
  assign n141 = n59 & n140 ;
  assign n142 = n52 & ~n141 ;
  assign n143 = x4 ^ x2 ;
  assign n144 = n143 ^ n45 ;
  assign n145 = ~x9 & n63 ;
  assign n146 = ~x13 & ~n41 ;
  assign n147 = n145 & ~n146 ;
  assign n148 = x9 & n43 ;
  assign n149 = ~n147 & ~n148 ;
  assign n150 = ~x8 & ~n149 ;
  assign n151 = n150 ^ x15 ;
  assign n152 = n151 ^ n143 ;
  assign n153 = x2 & ~n152 ;
  assign n154 = n153 ^ x15 ;
  assign n155 = n154 ^ x2 ;
  assign n156 = n155 ^ n143 ;
  assign n157 = n156 ^ n45 ;
  assign n158 = n144 & ~n157 ;
  assign n159 = n158 ^ n153 ;
  assign n160 = n159 ^ x15 ;
  assign n161 = n160 ^ n143 ;
  assign n162 = n45 & ~n161 ;
  assign n163 = n162 ^ n45 ;
  assign n164 = n163 ^ n45 ;
  assign n165 = ~n142 & ~n164 ;
  assign n166 = ~x0 & ~n165 ;
  assign n167 = x16 & n39 ;
  assign n168 = x4 ^ x1 ;
  assign n169 = n168 ^ x3 ;
  assign n170 = x20 ^ x4 ;
  assign n171 = n170 ^ x20 ;
  assign n172 = x13 & n70 ;
  assign n173 = x9 & n86 ;
  assign n174 = ~n172 & ~n173 ;
  assign n175 = ~x8 & n40 ;
  assign n176 = n86 & n175 ;
  assign n177 = x11 ^ x10 ;
  assign n178 = n176 & n177 ;
  assign n179 = n174 & ~n178 ;
  assign n180 = n179 ^ x20 ;
  assign n181 = ~n171 & ~n180 ;
  assign n182 = n181 ^ x20 ;
  assign n183 = n182 ^ n168 ;
  assign n184 = n169 & n183 ;
  assign n185 = n184 ^ n181 ;
  assign n186 = n185 ^ x20 ;
  assign n187 = n186 ^ x3 ;
  assign n188 = n168 & n187 ;
  assign n189 = n188 ^ n168 ;
  assign n190 = x0 & n189 ;
  assign n191 = n54 & n81 ;
  assign n192 = x13 ^ x0 ;
  assign n193 = x1 & n192 ;
  assign n194 = n193 ^ x0 ;
  assign n195 = ~n191 & ~n194 ;
  assign n196 = x15 & n52 ;
  assign n197 = ~n195 & n196 ;
  assign n198 = ~n190 & ~n197 ;
  assign n199 = ~x2 & ~n198 ;
  assign n200 = ~n167 & ~n199 ;
  assign n201 = ~n166 & n200 ;
  assign n202 = n201 ^ x5 ;
  assign n203 = n202 ^ n201 ;
  assign n204 = ~x1 & x2 ;
  assign n205 = n40 & n63 ;
  assign n206 = ~x4 & n205 ;
  assign n207 = n204 & n206 ;
  assign n208 = x8 & n173 ;
  assign n209 = x3 & n208 ;
  assign n210 = n207 & n209 ;
  assign n211 = x10 & ~x11 ;
  assign n212 = n47 & n211 ;
  assign n213 = ~n206 & ~n212 ;
  assign n214 = n208 & ~n213 ;
  assign n215 = n45 & n214 ;
  assign n216 = x2 & ~x22 ;
  assign n217 = n37 & ~n216 ;
  assign n218 = n217 ^ x3 ;
  assign n219 = n218 ^ n217 ;
  assign n220 = n219 ^ n215 ;
  assign n221 = n40 & n44 ;
  assign n222 = ~n81 & ~n221 ;
  assign n223 = ~x4 & ~n53 ;
  assign n224 = n88 & n223 ;
  assign n225 = ~n222 & n224 ;
  assign n226 = ~x8 & n148 ;
  assign n227 = ~n70 & ~n226 ;
  assign n228 = ~x4 & n227 ;
  assign n229 = ~x1 & ~n228 ;
  assign n230 = ~n225 & ~n229 ;
  assign n231 = n230 ^ x2 ;
  assign n232 = ~n230 & ~n231 ;
  assign n233 = n232 ^ n217 ;
  assign n234 = n233 ^ n230 ;
  assign n235 = n220 & ~n234 ;
  assign n236 = n235 ^ n232 ;
  assign n237 = n236 ^ n230 ;
  assign n238 = ~n215 & ~n237 ;
  assign n239 = n238 ^ n215 ;
  assign n240 = n239 ^ x0 ;
  assign n241 = n240 ^ n239 ;
  assign n242 = n241 ^ n210 ;
  assign n243 = x2 ^ x1 ;
  assign n244 = n61 ^ x11 ;
  assign n245 = n244 ^ n61 ;
  assign n246 = n61 ^ n44 ;
  assign n247 = ~n245 & n246 ;
  assign n248 = n247 ^ n61 ;
  assign n249 = n248 ^ x2 ;
  assign n250 = n243 & n249 ;
  assign n251 = n250 ^ n247 ;
  assign n252 = n251 ^ n61 ;
  assign n253 = n252 ^ x1 ;
  assign n254 = x2 & n253 ;
  assign n255 = n254 ^ x2 ;
  assign n256 = n173 & n255 ;
  assign n257 = ~x3 & ~n256 ;
  assign n258 = n40 & ~n257 ;
  assign n259 = ~x1 & x15 ;
  assign n260 = x22 & n259 ;
  assign n261 = n47 & n260 ;
  assign n262 = x21 & n261 ;
  assign n263 = ~n258 & ~n262 ;
  assign n264 = n47 & n226 ;
  assign n265 = x3 & ~n264 ;
  assign n266 = n265 ^ n263 ;
  assign n267 = ~n263 & n266 ;
  assign n268 = n267 ^ n239 ;
  assign n269 = n268 ^ n263 ;
  assign n270 = n242 & ~n269 ;
  assign n271 = n270 ^ n267 ;
  assign n272 = n271 ^ n263 ;
  assign n273 = ~n210 & ~n272 ;
  assign n274 = n273 ^ n210 ;
  assign n275 = n274 ^ n201 ;
  assign n276 = ~n203 & ~n275 ;
  assign n277 = n276 ^ n201 ;
  assign n278 = ~n51 & n277 ;
  assign n279 = n36 & ~n278 ;
  assign n280 = n35 & ~n279 ;
  assign y0 = ~n280 ;
endmodule
