module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 ;
  output y0 ;
  wire n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 ;
  assign n14 = ~x10 & x11 ;
  assign n15 = ~x7 & ~x9 ;
  assign n16 = x8 & ~x12 ;
  assign n17 = n15 & n16 ;
  assign n18 = n14 & n17 ;
  assign n19 = ~x6 & ~n18 ;
  assign n20 = ~x2 & x5 ;
  assign n21 = ~x3 & x4 ;
  assign n22 = x6 & ~x7 ;
  assign n23 = ~x0 & ~x1 ;
  assign n24 = ~n22 & n23 ;
  assign n25 = n21 & n24 ;
  assign n26 = n20 & n25 ;
  assign n27 = ~n19 & n26 ;
  assign y0 = n27 ;
endmodule
