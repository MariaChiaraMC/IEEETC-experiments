module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 ;
  assign n16 = ~x3 & x4 ;
  assign n17 = x1 ^ x0 ;
  assign n18 = ~x7 & ~x14 ;
  assign n19 = n18 ^ x13 ;
  assign n20 = n19 ^ x12 ;
  assign n21 = n18 ^ x12 ;
  assign n22 = ~x10 & ~x11 ;
  assign n23 = x9 ^ x8 ;
  assign n24 = n23 ^ x7 ;
  assign n25 = n24 ^ n22 ;
  assign n26 = x14 ^ x8 ;
  assign n27 = ~x7 & n26 ;
  assign n28 = n27 ^ x14 ;
  assign n29 = ~n25 & ~n28 ;
  assign n30 = n29 ^ n27 ;
  assign n31 = n30 ^ x14 ;
  assign n32 = n31 ^ x7 ;
  assign n33 = n22 & n32 ;
  assign n34 = n33 ^ x12 ;
  assign n35 = x12 & n34 ;
  assign n36 = n35 ^ x12 ;
  assign n37 = ~n21 & n36 ;
  assign n38 = n37 ^ n35 ;
  assign n39 = n38 ^ x12 ;
  assign n40 = n39 ^ n33 ;
  assign n41 = ~n20 & n40 ;
  assign n42 = ~x6 & ~n41 ;
  assign n43 = ~x2 & ~x5 ;
  assign n44 = ~n42 & n43 ;
  assign n45 = x1 & ~n44 ;
  assign n46 = n17 & n45 ;
  assign n47 = n46 ^ n17 ;
  assign n48 = n16 & n47 ;
  assign y0 = n48 ;
endmodule
