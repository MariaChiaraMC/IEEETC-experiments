module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n13 = ~x2 & x6 ;
  assign n14 = ~x0 & n13 ;
  assign n15 = ~x3 & ~x4 ;
  assign n16 = n14 & n15 ;
  assign n17 = ~x1 & n16 ;
  assign n18 = x9 ^ x8 ;
  assign n19 = x7 & n18 ;
  assign n20 = n19 ^ x5 ;
  assign n21 = n20 ^ n19 ;
  assign n22 = n21 ^ n17 ;
  assign n23 = ~x10 & ~x11 ;
  assign n24 = n23 ^ x7 ;
  assign n25 = ~n23 & ~n24 ;
  assign n26 = n25 ^ n19 ;
  assign n27 = n26 ^ n23 ;
  assign n28 = n22 & n27 ;
  assign n29 = n28 ^ n25 ;
  assign n30 = n29 ^ n23 ;
  assign n31 = n17 & ~n30 ;
  assign n32 = n31 ^ n17 ;
  assign y0 = n32 ;
endmodule
