// Benchmark "./adr4.pla" written by ABC on Thu Apr 23 10:59:45 2020

module \./adr4.pla  ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z4  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z4;
  assign z4 = 1'b1;
endmodule


