module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 ;
  assign n9 = x5 ^ x4 ;
  assign n10 = x3 ^ x2 ;
  assign n11 = n10 ^ x2 ;
  assign n12 = x6 ^ x2 ;
  assign n13 = ~n11 & ~n12 ;
  assign n14 = n13 ^ x2 ;
  assign n15 = n14 ^ x5 ;
  assign n16 = ~n9 & ~n15 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = n17 ^ x2 ;
  assign n19 = n18 ^ x4 ;
  assign n20 = ~x5 & n19 ;
  assign n21 = n20 ^ x5 ;
  assign n22 = x7 ^ x4 ;
  assign n23 = n22 ^ x2 ;
  assign n24 = n23 ^ x2 ;
  assign n25 = n24 ^ x3 ;
  assign n26 = x2 & n25 ;
  assign n27 = n26 ^ x2 ;
  assign n28 = n27 ^ x3 ;
  assign n29 = n24 ^ x4 ;
  assign n30 = n29 ^ n9 ;
  assign n31 = x6 ^ x4 ;
  assign n32 = n31 ^ n9 ;
  assign n33 = n30 & n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n34 ^ n29 ;
  assign n36 = n29 ^ x3 ;
  assign n37 = ~x3 & n36 ;
  assign n38 = n37 ^ n9 ;
  assign n39 = n38 ^ n31 ;
  assign n40 = n39 ^ x3 ;
  assign n41 = n35 & ~n40 ;
  assign n42 = n41 ^ n9 ;
  assign n43 = n42 ^ n24 ;
  assign n44 = n43 ^ n31 ;
  assign n45 = ~n28 & ~n44 ;
  assign n46 = n45 ^ x3 ;
  assign n47 = n21 & n46 ;
  assign n48 = ~x1 & n47 ;
  assign n49 = ~x0 & ~n48 ;
  assign y0 = n49 ;
endmodule
