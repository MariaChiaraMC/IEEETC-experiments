module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 ;
  assign n11 = ~x2 & x3 ;
  assign n14 = x7 & x8 ;
  assign n15 = x9 & n14 ;
  assign n16 = x5 & ~n15 ;
  assign n12 = ~x2 & x4 ;
  assign n13 = n12 ^ x1 ;
  assign n17 = n16 ^ n13 ;
  assign n18 = ~n11 & n17 ;
  assign n19 = n18 ^ n11 ;
  assign n20 = x2 & ~x3 ;
  assign n21 = x0 & ~n20 ;
  assign n22 = x6 & n21 ;
  assign n23 = n22 ^ n18 ;
  assign n24 = ~n13 & n23 ;
  assign n25 = n24 ^ n13 ;
  assign n26 = n25 ^ n16 ;
  assign n27 = ~n19 & n26 ;
  assign y0 = n27 ;
endmodule
