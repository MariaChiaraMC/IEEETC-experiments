module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ;
  assign n7 = x2 ^ x1 ;
  assign n8 = n7 ^ x3 ;
  assign n9 = n8 ^ x4 ;
  assign n10 = x5 ^ x3 ;
  assign n11 = n10 ^ x2 ;
  assign n12 = ~x2 & ~n11 ;
  assign n13 = n12 ^ x3 ;
  assign n14 = n13 ^ x2 ;
  assign n15 = x4 ^ x3 ;
  assign n16 = n15 ^ n9 ;
  assign n17 = n14 & n16 ;
  assign n18 = n17 ^ n12 ;
  assign n19 = n18 ^ x2 ;
  assign n20 = n9 & ~n19 ;
  assign n21 = n20 ^ x1 ;
  assign n22 = ~x0 & ~n21 ;
  assign n23 = ~x2 & ~x3 ;
  assign n24 = n23 ^ x1 ;
  assign n25 = n23 ^ x0 ;
  assign n26 = n25 ^ n23 ;
  assign n27 = n26 ^ n24 ;
  assign n28 = x4 & x5 ;
  assign n29 = ~x3 & ~n28 ;
  assign n30 = n29 ^ x4 ;
  assign n31 = ~n23 & ~n30 ;
  assign n32 = n31 ^ x4 ;
  assign n33 = n27 & n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n34 ^ x4 ;
  assign n36 = n35 ^ n23 ;
  assign n37 = n24 & ~n36 ;
  assign n38 = n37 ^ x1 ;
  assign n39 = ~n22 & ~n38 ;
  assign y0 = ~n39 ;
endmodule
