module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 ;
  assign n15 = ~x2 & x10 ;
  assign n16 = ~x3 & ~n15 ;
  assign n17 = ~x4 & ~x6 ;
  assign n18 = n17 ^ x6 ;
  assign n19 = ~x1 & n18 ;
  assign n20 = n19 ^ x6 ;
  assign n21 = ~n16 & n20 ;
  assign n22 = x5 & ~n21 ;
  assign n23 = x2 & x6 ;
  assign n24 = x9 & ~x12 ;
  assign n25 = ~x7 & ~x8 ;
  assign n26 = ~x11 & ~x13 ;
  assign n27 = ~x10 & n26 ;
  assign n28 = n25 & n27 ;
  assign n29 = n24 & n28 ;
  assign n30 = x4 & ~n29 ;
  assign n31 = n23 & ~n30 ;
  assign n32 = x3 & ~n31 ;
  assign n33 = ~x2 & n17 ;
  assign n34 = ~x3 & ~n33 ;
  assign n35 = ~x5 & ~n34 ;
  assign n36 = ~x0 & ~n35 ;
  assign n37 = x10 ^ x1 ;
  assign n38 = x2 ^ x1 ;
  assign n39 = n38 ^ x1 ;
  assign n40 = ~n37 & n39 ;
  assign n41 = n40 ^ x1 ;
  assign n42 = x1 & ~x6 ;
  assign n43 = n42 ^ x4 ;
  assign n44 = n41 & ~n43 ;
  assign n45 = n44 ^ n42 ;
  assign n46 = ~x4 & n45 ;
  assign n47 = n46 ^ x4 ;
  assign n48 = n47 ^ x4 ;
  assign n49 = n36 & ~n48 ;
  assign n50 = ~n32 & n49 ;
  assign n51 = ~n22 & n50 ;
  assign y0 = n51 ;
endmodule
