module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 ;
  output y0 ;
  wire n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 ;
  assign n49 = x11 & ~x13 ;
  assign n50 = x8 & ~x14 ;
  assign n51 = n49 & n50 ;
  assign n23 = ~x4 & ~x5 ;
  assign n52 = ~x6 & n23 ;
  assign n53 = x7 & n52 ;
  assign n54 = n51 & n53 ;
  assign n16 = x13 & x14 ;
  assign n17 = x11 & n16 ;
  assign n18 = ~x7 & ~x8 ;
  assign n19 = ~x0 & x14 ;
  assign n20 = ~x11 & ~x14 ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = ~n18 & ~n21 ;
  assign n24 = ~x13 & n23 ;
  assign n25 = x6 & n24 ;
  assign n26 = n22 & n25 ;
  assign n27 = ~x3 & x11 ;
  assign n28 = ~x6 & x14 ;
  assign n29 = n27 & n28 ;
  assign n30 = ~x13 & ~n29 ;
  assign n31 = ~x8 & ~x13 ;
  assign n32 = ~n20 & ~n31 ;
  assign n33 = x7 & ~n32 ;
  assign n34 = ~n30 & ~n33 ;
  assign n35 = x12 & ~n34 ;
  assign n36 = ~n26 & ~n35 ;
  assign n37 = ~n17 & n36 ;
  assign n38 = n37 ^ x11 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = x4 & x14 ;
  assign n41 = ~x13 & n40 ;
  assign n42 = ~x3 & ~n41 ;
  assign n43 = n42 ^ n37 ;
  assign n44 = n43 ^ n37 ;
  assign n45 = ~n39 & ~n44 ;
  assign n46 = n45 ^ n37 ;
  assign n47 = ~x9 & ~n46 ;
  assign n48 = n47 ^ n37 ;
  assign n55 = n54 ^ n48 ;
  assign n56 = n55 ^ n48 ;
  assign n57 = n48 ^ x9 ;
  assign n58 = n57 ^ n48 ;
  assign n59 = n56 & ~n58 ;
  assign n60 = n59 ^ n48 ;
  assign n61 = x10 & ~n60 ;
  assign n62 = n61 ^ n48 ;
  assign n63 = x10 & ~x11 ;
  assign n64 = ~x5 & x7 ;
  assign n65 = x4 & n64 ;
  assign n66 = x3 & n65 ;
  assign n67 = x13 & ~x14 ;
  assign n68 = ~x9 & n67 ;
  assign n69 = ~n66 & n68 ;
  assign n70 = x5 & ~x7 ;
  assign n71 = x4 & ~n70 ;
  assign n72 = x5 & x6 ;
  assign n73 = x0 & ~n72 ;
  assign n74 = n71 & ~n73 ;
  assign n75 = ~x3 & x13 ;
  assign n76 = x14 & n75 ;
  assign n77 = ~x9 & n76 ;
  assign n78 = n77 ^ x14 ;
  assign n79 = n74 & ~n78 ;
  assign n80 = ~n69 & ~n79 ;
  assign n81 = n63 & ~n80 ;
  assign n82 = ~x1 & ~x6 ;
  assign n83 = ~n27 & n82 ;
  assign n84 = n41 & ~n83 ;
  assign n85 = ~x9 & x10 ;
  assign n86 = ~x0 & n85 ;
  assign n87 = x5 & n86 ;
  assign n88 = n84 & n87 ;
  assign n89 = ~n81 & ~n88 ;
  assign n93 = ~x9 & ~x11 ;
  assign n90 = ~x10 & x11 ;
  assign n91 = x5 & ~x13 ;
  assign n92 = n90 & n91 ;
  assign n94 = n93 ^ n92 ;
  assign n95 = n94 ^ x14 ;
  assign n103 = n95 ^ n94 ;
  assign n96 = ~x10 & x13 ;
  assign n97 = n96 ^ n95 ;
  assign n98 = n97 ^ n94 ;
  assign n99 = n95 ^ n92 ;
  assign n100 = n99 ^ n96 ;
  assign n101 = n100 ^ n98 ;
  assign n102 = ~n98 & ~n101 ;
  assign n104 = n103 ^ n102 ;
  assign n105 = n104 ^ n98 ;
  assign n106 = n94 ^ x13 ;
  assign n107 = n102 ^ n98 ;
  assign n108 = ~n106 & ~n107 ;
  assign n109 = n108 ^ n94 ;
  assign n110 = ~n105 & n109 ;
  assign n111 = n110 ^ n94 ;
  assign n112 = n111 ^ n93 ;
  assign n113 = n112 ^ n94 ;
  assign n114 = ~x1 & n113 ;
  assign n115 = ~x0 & x11 ;
  assign n116 = ~x7 & ~x13 ;
  assign n117 = n115 & n116 ;
  assign n118 = ~x3 & x8 ;
  assign n119 = ~x6 & ~n118 ;
  assign n120 = ~x5 & x10 ;
  assign n121 = ~x4 & n120 ;
  assign n122 = ~n119 & n121 ;
  assign n123 = n117 & n122 ;
  assign n124 = ~x10 & ~x13 ;
  assign n125 = x14 & ~n71 ;
  assign n126 = ~n73 & ~n125 ;
  assign n127 = x10 & ~n16 ;
  assign n128 = ~n64 & ~n127 ;
  assign n129 = ~x11 & ~n128 ;
  assign n130 = n126 & n129 ;
  assign n131 = ~n124 & n130 ;
  assign n132 = n116 ^ n18 ;
  assign n133 = n18 ^ x6 ;
  assign n134 = n133 ^ n18 ;
  assign n135 = n134 ^ n121 ;
  assign n136 = ~n132 & n135 ;
  assign n137 = n136 ^ n116 ;
  assign n138 = n121 & n137 ;
  assign n139 = n138 ^ x4 ;
  assign n140 = n131 & n139 ;
  assign n141 = n96 ^ n90 ;
  assign n142 = n141 ^ x0 ;
  assign n150 = n142 ^ n141 ;
  assign n143 = n142 ^ n96 ;
  assign n144 = n143 ^ n142 ;
  assign n145 = n144 ^ n141 ;
  assign n146 = n143 ^ x14 ;
  assign n147 = n146 ^ n143 ;
  assign n148 = n147 ^ n145 ;
  assign n149 = n145 & n148 ;
  assign n151 = n150 ^ n149 ;
  assign n152 = n151 ^ n145 ;
  assign n153 = n141 ^ x1 ;
  assign n154 = n149 ^ n145 ;
  assign n155 = n153 & n154 ;
  assign n156 = n155 ^ n141 ;
  assign n157 = ~n152 & n156 ;
  assign n158 = n157 ^ n141 ;
  assign n159 = n158 ^ n90 ;
  assign n160 = n159 ^ n141 ;
  assign n161 = ~n140 & ~n160 ;
  assign n162 = ~n123 & n161 ;
  assign n163 = n162 ^ x9 ;
  assign n164 = n163 ^ n162 ;
  assign n165 = n164 ^ n114 ;
  assign n166 = x10 ^ x3 ;
  assign n167 = ~x10 & ~n166 ;
  assign n168 = n167 ^ n162 ;
  assign n169 = n168 ^ x10 ;
  assign n170 = n165 & n169 ;
  assign n171 = n170 ^ n167 ;
  assign n172 = n171 ^ x10 ;
  assign n173 = ~n114 & ~n172 ;
  assign n174 = n173 ^ n114 ;
  assign n175 = n89 & ~n174 ;
  assign n176 = n175 ^ x12 ;
  assign n177 = n176 ^ n175 ;
  assign n178 = n31 & n64 ;
  assign n179 = n28 & n178 ;
  assign n180 = ~n49 & ~n179 ;
  assign n181 = ~x4 & ~n180 ;
  assign n182 = ~n82 & n91 ;
  assign n183 = ~x2 & n182 ;
  assign n184 = x1 & n67 ;
  assign n185 = n65 & n184 ;
  assign n186 = ~n183 & ~n185 ;
  assign n187 = n115 & ~n186 ;
  assign n188 = ~n181 & ~n187 ;
  assign n189 = n85 & ~n188 ;
  assign n190 = ~x10 & n93 ;
  assign n191 = n40 & n190 ;
  assign n192 = ~x5 & n124 ;
  assign n193 = x6 & ~x11 ;
  assign n194 = ~x10 & n193 ;
  assign n195 = ~n192 & ~n194 ;
  assign n196 = x9 & ~n195 ;
  assign n197 = n52 & n63 ;
  assign n198 = n76 & n197 ;
  assign n199 = ~n196 & ~n198 ;
  assign n200 = ~x7 & x8 ;
  assign n201 = ~n199 & n200 ;
  assign n202 = ~n191 & ~n201 ;
  assign n203 = ~n189 & n202 ;
  assign n204 = n203 ^ n175 ;
  assign n205 = n177 & n204 ;
  assign n206 = n205 ^ n175 ;
  assign n207 = n62 & n206 ;
  assign y0 = ~n207 ;
endmodule
