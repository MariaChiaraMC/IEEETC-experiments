module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 ;
  assign n17 = x2 & ~x8 ;
  assign n18 = ~x14 & x15 ;
  assign n19 = n17 & n18 ;
  assign n20 = x4 & x9 ;
  assign n21 = n19 & n20 ;
  assign n22 = ~x1 & x10 ;
  assign n23 = x5 & ~x6 ;
  assign n24 = ~x3 & x13 ;
  assign n25 = n23 & n24 ;
  assign n26 = n22 & n25 ;
  assign n27 = n21 & n26 ;
  assign n28 = ~x3 & ~x5 ;
  assign n29 = x6 & n28 ;
  assign n30 = n17 & n29 ;
  assign n31 = ~x10 & ~x14 ;
  assign n32 = ~x4 & x9 ;
  assign n33 = ~x7 & n32 ;
  assign n34 = n31 & n33 ;
  assign n35 = n30 & n34 ;
  assign n36 = x8 ^ x2 ;
  assign n37 = x5 ^ x2 ;
  assign n38 = n36 & n37 ;
  assign n39 = ~x6 & n38 ;
  assign n40 = x7 & n39 ;
  assign n41 = x3 & n40 ;
  assign n42 = ~x14 & ~n41 ;
  assign n43 = n32 & ~n42 ;
  assign n44 = ~x6 & ~x8 ;
  assign n45 = ~x7 & n44 ;
  assign n46 = x6 & x7 ;
  assign n47 = x8 & n46 ;
  assign n48 = ~n45 & ~n47 ;
  assign n49 = x3 & x4 ;
  assign n50 = x2 & ~x9 ;
  assign n51 = n49 & n50 ;
  assign n52 = ~n48 & n51 ;
  assign n53 = x5 & n52 ;
  assign n54 = ~n43 & ~n53 ;
  assign n55 = ~x2 & x8 ;
  assign n56 = ~x7 & x11 ;
  assign n57 = n55 & n56 ;
  assign n58 = n29 & n32 ;
  assign n59 = n57 & n58 ;
  assign n60 = x14 & ~n59 ;
  assign n61 = x10 & ~n60 ;
  assign n62 = ~n54 & n61 ;
  assign n63 = ~n35 & ~n62 ;
  assign n64 = ~x15 & ~n63 ;
  assign n65 = ~x4 & ~x10 ;
  assign n66 = ~x2 & x14 ;
  assign n67 = n65 & n66 ;
  assign n68 = ~x9 & x15 ;
  assign n69 = n28 & n68 ;
  assign n70 = n45 & n69 ;
  assign n71 = n67 & n70 ;
  assign n72 = ~n64 & ~n71 ;
  assign n73 = ~x1 & ~n72 ;
  assign n74 = x6 & ~x7 ;
  assign n75 = x10 & n74 ;
  assign n76 = x5 & x7 ;
  assign n77 = ~x10 & n46 ;
  assign n78 = ~n76 & ~n77 ;
  assign n79 = x1 & x9 ;
  assign n80 = n19 & n79 ;
  assign n81 = n78 & n80 ;
  assign n82 = n49 & n81 ;
  assign n83 = ~n75 & n82 ;
  assign n84 = ~n73 & ~n83 ;
  assign n85 = ~x13 & ~n84 ;
  assign n86 = ~n27 & ~n85 ;
  assign n87 = ~x0 & ~n86 ;
  assign n88 = ~x5 & n18 ;
  assign n89 = x1 & n46 ;
  assign n90 = x0 & ~x13 ;
  assign n91 = n49 & n90 ;
  assign n92 = n89 & n91 ;
  assign n93 = n88 & n92 ;
  assign n94 = ~x2 & n93 ;
  assign n95 = ~n87 & ~n94 ;
  assign n96 = ~x12 & ~n95 ;
  assign y0 = n96 ;
endmodule
