// Benchmark "./wim.pla" written by ABC on Thu Apr 23 11:00:08 2020

module \./wim.pla  ( 
    x0, x1, x2, x3,
    z3  );
  input  x0, x1, x2, x3;
  output z3;
  assign z3 = ~x1 | x2;
endmodule


