module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 ;
  assign n17 = x7 & x12 ;
  assign n18 = x9 & x10 ;
  assign n19 = ~x1 & ~x13 ;
  assign n20 = x0 & ~x2 ;
  assign n21 = ~x3 & ~x4 ;
  assign n22 = n20 & n21 ;
  assign n23 = ~n19 & n22 ;
  assign n24 = ~x13 & ~x14 ;
  assign n25 = ~x0 & ~x3 ;
  assign n26 = ~x4 & x5 ;
  assign n27 = n25 & n26 ;
  assign n28 = x1 & ~x13 ;
  assign n29 = x1 & ~x14 ;
  assign n30 = ~n28 & ~n29 ;
  assign n31 = n27 & n30 ;
  assign n32 = x1 & ~x2 ;
  assign n33 = ~x3 & n32 ;
  assign n34 = ~x0 & ~x5 ;
  assign n35 = n33 & n34 ;
  assign n36 = ~n31 & ~n35 ;
  assign n37 = ~n24 & ~n36 ;
  assign n38 = ~x1 & x3 ;
  assign n39 = ~x5 & x13 ;
  assign n40 = ~x2 & ~x4 ;
  assign n41 = n39 & n40 ;
  assign n42 = x2 & ~x4 ;
  assign n43 = ~x0 & n42 ;
  assign n44 = ~x2 & x14 ;
  assign n45 = ~x0 & ~x13 ;
  assign n46 = ~x5 & n45 ;
  assign n47 = n44 & n46 ;
  assign n48 = ~n43 & ~n47 ;
  assign n49 = ~n41 & n48 ;
  assign n50 = n38 & ~n49 ;
  assign n51 = ~n37 & ~n50 ;
  assign n52 = ~n23 & n51 ;
  assign n53 = n52 ^ x11 ;
  assign n54 = n53 ^ n52 ;
  assign n55 = x1 & ~x3 ;
  assign n56 = ~n38 & ~n55 ;
  assign n57 = ~x1 & x13 ;
  assign n58 = x0 & x2 ;
  assign n59 = ~n57 & n58 ;
  assign n60 = ~x0 & x14 ;
  assign n61 = ~x3 & n60 ;
  assign n62 = ~n59 & ~n61 ;
  assign n63 = n56 & ~n62 ;
  assign n64 = x5 & n63 ;
  assign n65 = x2 & x3 ;
  assign n66 = ~x0 & ~x1 ;
  assign n67 = n65 & n66 ;
  assign n68 = x0 & ~x3 ;
  assign n69 = n32 & n68 ;
  assign n70 = ~n67 & ~n69 ;
  assign n71 = ~n24 & ~n70 ;
  assign n72 = ~x4 & ~n71 ;
  assign n73 = ~n64 & n72 ;
  assign n74 = ~x1 & ~x2 ;
  assign n75 = ~x0 & x5 ;
  assign n76 = ~x13 & x14 ;
  assign n77 = n75 & n76 ;
  assign n78 = n74 & n77 ;
  assign n79 = x1 & ~x5 ;
  assign n80 = ~x3 & n58 ;
  assign n81 = n79 & n80 ;
  assign n82 = x4 & ~n81 ;
  assign n83 = ~n78 & n82 ;
  assign n84 = ~n73 & ~n83 ;
  assign n85 = ~x5 & x14 ;
  assign n86 = ~x0 & n85 ;
  assign n87 = n86 ^ x13 ;
  assign n88 = n87 ^ n86 ;
  assign n89 = x0 & x5 ;
  assign n90 = ~x4 & n89 ;
  assign n91 = n90 ^ n86 ;
  assign n92 = n91 ^ n86 ;
  assign n93 = n88 & n92 ;
  assign n94 = n93 ^ n86 ;
  assign n95 = x2 & n94 ;
  assign n96 = n95 ^ n86 ;
  assign n97 = ~n56 & n96 ;
  assign n98 = ~n84 & ~n97 ;
  assign n99 = n98 ^ n52 ;
  assign n100 = ~n54 & n99 ;
  assign n101 = n100 ^ n52 ;
  assign n102 = x8 & ~n101 ;
  assign n103 = n18 & n102 ;
  assign n104 = ~x9 & x10 ;
  assign n105 = x11 & x13 ;
  assign n106 = ~x4 & x8 ;
  assign n107 = n67 & n106 ;
  assign n108 = n105 & n107 ;
  assign n109 = ~x1 & x11 ;
  assign n110 = x3 & x13 ;
  assign n112 = x2 & ~x8 ;
  assign n111 = ~x2 & x8 ;
  assign n113 = n112 ^ n111 ;
  assign n114 = n113 ^ n112 ;
  assign n115 = n112 ^ x15 ;
  assign n116 = n115 ^ n112 ;
  assign n117 = n114 & n116 ;
  assign n118 = n117 ^ n112 ;
  assign n119 = n110 & n118 ;
  assign n120 = n119 ^ n112 ;
  assign n121 = n109 & n120 ;
  assign n122 = ~x0 & x11 ;
  assign n124 = ~x3 & x8 ;
  assign n123 = x13 & n65 ;
  assign n125 = n124 ^ n123 ;
  assign n126 = x1 & x13 ;
  assign n127 = x15 & n126 ;
  assign n128 = n127 ^ n123 ;
  assign n129 = n123 ^ x1 ;
  assign n130 = ~n123 & ~n129 ;
  assign n131 = n130 ^ n123 ;
  assign n132 = ~n128 & ~n131 ;
  assign n133 = n132 ^ n130 ;
  assign n134 = n133 ^ n123 ;
  assign n135 = n134 ^ x1 ;
  assign n136 = n125 & ~n135 ;
  assign n137 = n136 ^ n124 ;
  assign n138 = n122 & n137 ;
  assign n139 = ~n121 & ~n138 ;
  assign n140 = n26 & ~n139 ;
  assign n145 = x13 & x15 ;
  assign n146 = ~x4 & ~x8 ;
  assign n147 = n145 & n146 ;
  assign n141 = x1 & x2 ;
  assign n142 = ~n74 & ~n141 ;
  assign n143 = x5 & ~n142 ;
  assign n144 = ~n65 & n143 ;
  assign n148 = n147 ^ n144 ;
  assign n149 = n144 ^ n33 ;
  assign n150 = n149 ^ n33 ;
  assign n151 = x8 & ~x13 ;
  assign n152 = x4 & n151 ;
  assign n153 = n152 ^ n33 ;
  assign n154 = n150 & ~n153 ;
  assign n155 = n154 ^ n33 ;
  assign n156 = n148 & ~n155 ;
  assign n157 = n156 ^ n147 ;
  assign n158 = n122 & n157 ;
  assign n159 = ~x1 & x5 ;
  assign n160 = ~n79 & ~n159 ;
  assign n161 = ~x8 & n160 ;
  assign n162 = ~x3 & ~x8 ;
  assign n163 = ~x3 & ~x13 ;
  assign n164 = x1 & x5 ;
  assign n165 = n163 & n164 ;
  assign n166 = ~n162 & ~n165 ;
  assign n167 = ~n161 & ~n166 ;
  assign n168 = x3 & x5 ;
  assign n169 = ~x1 & n168 ;
  assign n170 = ~n167 & ~n169 ;
  assign n171 = n43 & ~n170 ;
  assign n172 = n171 ^ x11 ;
  assign n173 = n172 ^ n171 ;
  assign n174 = n173 ^ n158 ;
  assign n175 = ~x0 & x8 ;
  assign n176 = x2 & ~x13 ;
  assign n177 = x3 & n176 ;
  assign n178 = ~x1 & ~x4 ;
  assign n179 = n177 & n178 ;
  assign n180 = ~x2 & ~x5 ;
  assign n181 = n56 & ~n127 ;
  assign n182 = n180 & ~n181 ;
  assign n183 = ~n179 & ~n182 ;
  assign n184 = n183 ^ n175 ;
  assign n185 = n175 & ~n184 ;
  assign n186 = n185 ^ n171 ;
  assign n187 = n186 ^ n175 ;
  assign n188 = ~n174 & n187 ;
  assign n189 = n188 ^ n185 ;
  assign n190 = n189 ^ n175 ;
  assign n191 = ~n158 & n190 ;
  assign n192 = n191 ^ n158 ;
  assign n193 = ~n140 & ~n192 ;
  assign n194 = x14 & ~n193 ;
  assign n195 = x0 & ~x4 ;
  assign n196 = ~x3 & x5 ;
  assign n197 = x1 & x11 ;
  assign n198 = x2 & x8 ;
  assign n199 = x13 & n198 ;
  assign n200 = ~x8 & n76 ;
  assign n201 = ~n199 & ~n200 ;
  assign n202 = n197 & ~n201 ;
  assign n203 = ~x14 & ~n176 ;
  assign n204 = n109 & ~n112 ;
  assign n205 = x14 & n32 ;
  assign n206 = ~x1 & ~x8 ;
  assign n207 = ~n205 & ~n206 ;
  assign n208 = ~x11 & ~n207 ;
  assign n209 = ~n204 & ~n208 ;
  assign n210 = ~n203 & ~n209 ;
  assign n211 = ~n202 & ~n210 ;
  assign n212 = n196 & ~n211 ;
  assign n213 = x2 & ~x5 ;
  assign n214 = ~x1 & x8 ;
  assign n215 = x11 & n214 ;
  assign n216 = n213 & n215 ;
  assign n217 = ~x3 & x11 ;
  assign n218 = ~n24 & n32 ;
  assign n219 = n217 & n218 ;
  assign n220 = x8 & n219 ;
  assign n221 = ~n216 & ~n220 ;
  assign n222 = ~n212 & n221 ;
  assign n223 = n195 & ~n222 ;
  assign n224 = x0 & x3 ;
  assign n225 = ~x4 & x14 ;
  assign n226 = x2 & ~x11 ;
  assign n227 = x1 & ~x8 ;
  assign n228 = ~x13 & n227 ;
  assign n229 = n226 & n228 ;
  assign n230 = x8 & ~x11 ;
  assign n231 = ~x13 & n230 ;
  assign n232 = ~x2 & x5 ;
  assign n233 = ~x1 & n232 ;
  assign n234 = n231 & n233 ;
  assign n235 = x11 & n232 ;
  assign n236 = n126 & n235 ;
  assign n237 = ~n234 & ~n236 ;
  assign n238 = ~n229 & n237 ;
  assign n239 = n225 & ~n238 ;
  assign n240 = ~x11 & ~x13 ;
  assign n241 = n146 & ~n240 ;
  assign n242 = x4 & ~x11 ;
  assign n243 = ~x5 & n242 ;
  assign n244 = ~n241 & ~n243 ;
  assign n245 = n141 & ~n244 ;
  assign n246 = x5 & x8 ;
  assign n247 = ~x1 & n246 ;
  assign n248 = x11 & ~x13 ;
  assign n249 = x4 & x14 ;
  assign n250 = ~x2 & n249 ;
  assign n251 = n248 & n250 ;
  assign n252 = n247 & n251 ;
  assign n253 = ~n245 & ~n252 ;
  assign n254 = ~n239 & n253 ;
  assign n255 = n224 & ~n254 ;
  assign n256 = ~n223 & ~n255 ;
  assign n257 = ~n194 & n256 ;
  assign n258 = ~n108 & n257 ;
  assign n259 = n104 & ~n258 ;
  assign n260 = ~x11 & x14 ;
  assign n261 = x0 & ~x1 ;
  assign n262 = ~x2 & ~x3 ;
  assign n263 = x8 & x9 ;
  assign n264 = n262 & n263 ;
  assign n265 = ~x8 & ~x9 ;
  assign n266 = n65 & n265 ;
  assign n267 = ~n264 & ~n266 ;
  assign n268 = n261 & ~n267 ;
  assign n269 = ~x8 & n58 ;
  assign n270 = ~x9 & n55 ;
  assign n271 = n269 & n270 ;
  assign n272 = ~n268 & ~n271 ;
  assign n273 = n26 & ~n272 ;
  assign n274 = ~x0 & x15 ;
  assign n275 = ~x3 & n263 ;
  assign n276 = ~x3 & ~x9 ;
  assign n277 = x2 & ~x9 ;
  assign n278 = ~n276 & n277 ;
  assign n279 = ~n275 & ~n278 ;
  assign n280 = n274 & ~n279 ;
  assign n281 = x0 & x15 ;
  assign n282 = ~x8 & x9 ;
  assign n283 = ~x3 & n282 ;
  assign n284 = x3 & ~x9 ;
  assign n285 = ~x2 & n284 ;
  assign n286 = ~n283 & ~n285 ;
  assign n287 = n281 & ~n286 ;
  assign n288 = ~n280 & ~n287 ;
  assign n289 = n26 & ~n288 ;
  assign n290 = x9 & x15 ;
  assign n291 = ~x2 & n224 ;
  assign n292 = ~x5 & ~x8 ;
  assign n293 = n291 & n292 ;
  assign n294 = n290 & n293 ;
  assign n295 = ~n289 & ~n294 ;
  assign n296 = n126 & ~n295 ;
  assign n297 = ~n273 & ~n296 ;
  assign n298 = n260 & ~n297 ;
  assign n299 = ~x8 & n18 ;
  assign n300 = ~x5 & n65 ;
  assign n301 = ~x3 & n44 ;
  assign n302 = ~x4 & x15 ;
  assign n303 = n301 & n302 ;
  assign n304 = ~n300 & ~n303 ;
  assign n305 = n66 & ~n304 ;
  assign n306 = x0 & x1 ;
  assign n307 = x14 & n306 ;
  assign n308 = ~x3 & n26 ;
  assign n309 = n307 & n308 ;
  assign n310 = ~x2 & n306 ;
  assign n311 = x14 & x15 ;
  assign n312 = x3 & ~x4 ;
  assign n313 = n311 & n312 ;
  assign n314 = x3 & ~x14 ;
  assign n315 = ~x5 & ~n314 ;
  assign n316 = ~n313 & ~n315 ;
  assign n317 = n310 & ~n316 ;
  assign n318 = x2 & ~x3 ;
  assign n319 = x5 & x15 ;
  assign n320 = n318 & n319 ;
  assign n321 = n178 & n320 ;
  assign n322 = x14 & n321 ;
  assign n323 = ~n317 & ~n322 ;
  assign n324 = ~n309 & n323 ;
  assign n325 = ~n305 & n324 ;
  assign n326 = n105 & ~n325 ;
  assign n327 = x0 & n74 ;
  assign n328 = ~x3 & x14 ;
  assign n329 = ~x5 & x11 ;
  assign n330 = n328 & n329 ;
  assign n331 = n327 & n330 ;
  assign n332 = ~x1 & x2 ;
  assign n333 = n68 & n332 ;
  assign n334 = ~x13 & n260 ;
  assign n335 = n26 & n334 ;
  assign n336 = n333 & n335 ;
  assign n337 = ~n331 & ~n336 ;
  assign n338 = ~n326 & n337 ;
  assign n339 = n299 & ~n338 ;
  assign n340 = ~n298 & ~n339 ;
  assign n341 = ~n259 & n340 ;
  assign n342 = ~n103 & n341 ;
  assign n343 = n17 & ~n342 ;
  assign n344 = ~x1 & ~x5 ;
  assign n345 = ~x3 & n344 ;
  assign n346 = ~x9 & ~x11 ;
  assign n347 = n345 & n346 ;
  assign n348 = x1 & x3 ;
  assign n349 = x5 & n348 ;
  assign n350 = x2 & n349 ;
  assign n351 = ~n347 & ~n350 ;
  assign n352 = x2 & x4 ;
  assign n353 = n68 & n352 ;
  assign n354 = ~x9 & ~x10 ;
  assign n355 = x8 & ~n354 ;
  assign n356 = ~n353 & n355 ;
  assign n357 = ~n40 & ~n312 ;
  assign n358 = n356 & n357 ;
  assign n359 = ~n351 & n358 ;
  assign n360 = x4 & n318 ;
  assign n361 = ~x0 & ~n360 ;
  assign n362 = n359 & ~n361 ;
  assign n363 = x7 & x14 ;
  assign n364 = x2 & ~x12 ;
  assign n365 = ~x5 & x8 ;
  assign n366 = ~x3 & x4 ;
  assign n367 = ~x0 & n366 ;
  assign n368 = n18 & n248 ;
  assign n369 = n367 & n368 ;
  assign n370 = x1 & x9 ;
  assign n371 = x0 & x10 ;
  assign n372 = n370 & ~n371 ;
  assign n373 = ~x0 & x3 ;
  assign n374 = ~n346 & n373 ;
  assign n375 = x3 & x9 ;
  assign n376 = ~x1 & x4 ;
  assign n377 = ~n375 & n376 ;
  assign n378 = ~n374 & n377 ;
  assign n379 = x10 & n378 ;
  assign n380 = ~n372 & ~n379 ;
  assign n381 = ~x0 & ~x10 ;
  assign n382 = ~n276 & ~n381 ;
  assign n383 = x3 & x11 ;
  assign n384 = ~n66 & ~n383 ;
  assign n385 = n382 & ~n384 ;
  assign n386 = ~n380 & n385 ;
  assign n387 = x13 & n386 ;
  assign n388 = ~n369 & ~n387 ;
  assign n389 = n365 & ~n388 ;
  assign n390 = x4 & x10 ;
  assign n391 = ~x0 & n390 ;
  assign n392 = ~x11 & x13 ;
  assign n393 = ~x9 & n392 ;
  assign n394 = n247 & n393 ;
  assign n395 = ~x1 & x9 ;
  assign n396 = x1 & ~x9 ;
  assign n397 = ~n395 & ~n396 ;
  assign n398 = n163 & ~n263 ;
  assign n399 = ~n230 & n398 ;
  assign n400 = ~n397 & n399 ;
  assign n401 = ~n394 & ~n400 ;
  assign n402 = n391 & ~n401 ;
  assign n403 = ~x5 & n306 ;
  assign n404 = x9 & ~x13 ;
  assign n405 = x3 & x10 ;
  assign n406 = ~x8 & ~x11 ;
  assign n407 = n405 & n406 ;
  assign n408 = n404 & n407 ;
  assign n409 = n403 & n408 ;
  assign n410 = ~n402 & ~n409 ;
  assign n411 = x5 & x10 ;
  assign n412 = n105 & n206 ;
  assign n413 = n281 & n412 ;
  assign n414 = x11 & x15 ;
  assign n415 = ~x8 & n414 ;
  assign n416 = ~n151 & ~n415 ;
  assign n417 = n66 & ~n416 ;
  assign n418 = ~x8 & ~x13 ;
  assign n419 = ~x11 & ~n145 ;
  assign n420 = ~n418 & n419 ;
  assign n421 = ~n248 & n306 ;
  assign n422 = ~n420 & n421 ;
  assign n423 = ~n417 & ~n422 ;
  assign n424 = ~n413 & n423 ;
  assign n425 = n284 & ~n424 ;
  assign n426 = n214 & n375 ;
  assign n427 = ~x11 & x15 ;
  assign n428 = ~n240 & ~n427 ;
  assign n429 = n426 & ~n428 ;
  assign n430 = ~x8 & x13 ;
  assign n431 = n414 & n430 ;
  assign n432 = n55 & n431 ;
  assign n433 = ~n19 & ~n432 ;
  assign n434 = x0 & ~x9 ;
  assign n435 = ~n230 & n434 ;
  assign n436 = ~n433 & n435 ;
  assign n437 = ~n429 & ~n436 ;
  assign n438 = x9 & ~x11 ;
  assign n439 = ~x3 & n438 ;
  assign n440 = n439 ^ x0 ;
  assign n441 = n440 ^ n439 ;
  assign n442 = ~x1 & ~x3 ;
  assign n443 = n442 ^ n439 ;
  assign n444 = ~n441 & n443 ;
  assign n445 = n444 ^ n439 ;
  assign n446 = ~x13 & n445 ;
  assign n447 = x8 & n446 ;
  assign n448 = n437 & ~n447 ;
  assign n449 = ~n425 & n448 ;
  assign n450 = n411 & ~n449 ;
  assign n451 = x10 & n56 ;
  assign n452 = ~x11 & n89 ;
  assign n453 = ~x1 & ~x10 ;
  assign n454 = x9 & ~n453 ;
  assign n455 = n452 & ~n454 ;
  assign n456 = ~x8 & x15 ;
  assign n457 = n456 ^ n151 ;
  assign n458 = n348 & n457 ;
  assign n459 = n458 ^ n151 ;
  assign n460 = n455 & n459 ;
  assign n461 = ~n451 & n460 ;
  assign n462 = x1 & ~x11 ;
  assign n463 = x8 & x10 ;
  assign n464 = ~x13 & n463 ;
  assign n465 = x8 & ~x10 ;
  assign n466 = ~x8 & x10 ;
  assign n467 = ~n465 & ~n466 ;
  assign n468 = n39 & ~n467 ;
  assign n469 = ~n464 & ~n468 ;
  assign n470 = n462 & ~n469 ;
  assign n471 = ~x10 & x11 ;
  assign n472 = n28 & n471 ;
  assign n473 = x10 & x13 ;
  assign n474 = ~x11 & n473 ;
  assign n475 = ~n472 & ~n474 ;
  assign n476 = n365 & ~n475 ;
  assign n477 = ~n470 & ~n476 ;
  assign n478 = n284 & ~n477 ;
  assign n479 = ~x1 & n124 ;
  assign n480 = n368 & n479 ;
  assign n481 = ~n478 & ~n480 ;
  assign n482 = x0 & ~n481 ;
  assign n483 = ~n461 & ~n482 ;
  assign n484 = ~n450 & n483 ;
  assign n485 = ~x4 & ~n484 ;
  assign n486 = n410 & ~n485 ;
  assign n487 = ~n389 & n486 ;
  assign n488 = n364 & ~n487 ;
  assign n489 = ~x0 & x10 ;
  assign n490 = n414 & n489 ;
  assign n491 = ~x1 & n490 ;
  assign n492 = ~x3 & x9 ;
  assign n493 = n246 & n492 ;
  assign n494 = n491 & n493 ;
  assign n495 = n40 & n494 ;
  assign n496 = x4 & ~x9 ;
  assign n497 = x5 & x13 ;
  assign n498 = ~x11 & n497 ;
  assign n499 = n496 & n498 ;
  assign n500 = x5 ^ x4 ;
  assign n501 = n404 ^ x5 ;
  assign n502 = n501 ^ n404 ;
  assign n503 = ~x9 & x13 ;
  assign n504 = n503 ^ n404 ;
  assign n505 = ~n502 & n504 ;
  assign n506 = n505 ^ n404 ;
  assign n507 = n500 & n506 ;
  assign n508 = n462 & n507 ;
  assign n509 = ~n499 & ~n508 ;
  assign n510 = x10 & ~n509 ;
  assign n511 = ~x10 & x15 ;
  assign n512 = n438 & n511 ;
  assign n513 = x1 & ~x4 ;
  assign n514 = x5 & n513 ;
  assign n515 = n512 & n514 ;
  assign n516 = n178 & n411 ;
  assign n517 = x9 & x11 ;
  assign n518 = n145 & n517 ;
  assign n519 = x13 & ~n518 ;
  assign n520 = n516 & ~n519 ;
  assign n521 = ~n515 & ~n520 ;
  assign n522 = ~n510 & n521 ;
  assign n523 = n124 & ~n522 ;
  assign n537 = n196 & n513 ;
  assign n524 = x10 & x11 ;
  assign n525 = ~x13 & n524 ;
  assign n526 = x5 & x9 ;
  assign n527 = ~n276 & ~n526 ;
  assign n528 = n525 & n527 ;
  assign n529 = ~x3 & x10 ;
  assign n530 = x9 & x13 ;
  assign n531 = ~x5 & n530 ;
  assign n532 = n529 & n531 ;
  assign n533 = ~n528 & ~n532 ;
  assign n534 = n376 & ~n533 ;
  assign n538 = n537 ^ n534 ;
  assign n539 = n538 ^ n534 ;
  assign n535 = n534 ^ n414 ;
  assign n536 = n535 ^ n534 ;
  assign n540 = n539 ^ n536 ;
  assign n541 = n534 ^ n104 ;
  assign n542 = n541 ^ n534 ;
  assign n543 = n542 ^ n539 ;
  assign n544 = n539 & n543 ;
  assign n545 = n544 ^ n539 ;
  assign n546 = n540 & n545 ;
  assign n547 = n546 ^ n544 ;
  assign n548 = n547 ^ n534 ;
  assign n549 = n548 ^ n539 ;
  assign n550 = ~x8 & n549 ;
  assign n551 = n550 ^ n534 ;
  assign n552 = ~n523 & ~n551 ;
  assign n553 = n20 & ~n552 ;
  assign n554 = ~x9 & x11 ;
  assign n555 = ~n438 & ~n554 ;
  assign n556 = x4 & ~x8 ;
  assign n557 = ~x10 & ~x13 ;
  assign n558 = ~x3 & n261 ;
  assign n559 = n557 & n558 ;
  assign n560 = n556 & n559 ;
  assign n561 = x3 & ~x5 ;
  assign n562 = x1 & x8 ;
  assign n563 = n489 & n562 ;
  assign n564 = n145 & n563 ;
  assign n565 = n561 & n564 ;
  assign n566 = ~n560 & ~n565 ;
  assign n567 = x2 & ~n566 ;
  assign n568 = x1 & x10 ;
  assign n569 = x8 & n568 ;
  assign n570 = n195 & n196 ;
  assign n571 = x0 & ~x5 ;
  assign n572 = ~x2 & n571 ;
  assign n573 = x3 & n572 ;
  assign n574 = ~n570 & ~n573 ;
  assign n575 = n145 & ~n574 ;
  assign n576 = n569 & n575 ;
  assign n577 = ~n567 & ~n576 ;
  assign n578 = ~n555 & ~n577 ;
  assign n579 = x13 & n263 ;
  assign n580 = n570 & n579 ;
  assign n581 = x1 & n524 ;
  assign n582 = n580 & n581 ;
  assign n583 = ~n578 & ~n582 ;
  assign n584 = ~n553 & n583 ;
  assign n585 = ~n495 & n584 ;
  assign n586 = ~x12 & ~n585 ;
  assign n587 = ~x13 & n197 ;
  assign n588 = n124 & n277 ;
  assign n589 = n90 & n588 ;
  assign n590 = n295 & ~n589 ;
  assign n591 = n587 & ~n590 ;
  assign n592 = n112 & n224 ;
  assign n593 = n329 & n404 ;
  assign n594 = n592 & n593 ;
  assign n595 = n75 & n346 ;
  assign n596 = x8 & x13 ;
  assign n597 = n262 & n596 ;
  assign n598 = n595 & n597 ;
  assign n599 = ~n594 & ~n598 ;
  assign n600 = n376 & ~n599 ;
  assign n601 = ~n591 & ~n600 ;
  assign n602 = n601 ^ x10 ;
  assign n603 = n602 ^ n601 ;
  assign n604 = n603 ^ n586 ;
  assign n605 = x15 & n248 ;
  assign n606 = n90 & ~n279 ;
  assign n607 = x9 & n175 ;
  assign n608 = n300 & n607 ;
  assign n609 = ~n606 & ~n608 ;
  assign n610 = n605 & ~n609 ;
  assign n611 = n610 ^ x1 ;
  assign n612 = x1 & n611 ;
  assign n613 = n612 ^ n601 ;
  assign n614 = n613 ^ x1 ;
  assign n615 = n604 & ~n614 ;
  assign n616 = n615 ^ n612 ;
  assign n617 = n616 ^ x1 ;
  assign n618 = ~n586 & n617 ;
  assign n619 = n618 ^ n586 ;
  assign n620 = ~n488 & ~n619 ;
  assign n621 = n363 & ~n620 ;
  assign n622 = x7 & ~x10 ;
  assign n623 = x11 & x14 ;
  assign n624 = ~x5 & ~x13 ;
  assign n625 = n623 & n624 ;
  assign n626 = n26 & n392 ;
  assign n627 = ~n625 & ~n626 ;
  assign n628 = n434 & ~n627 ;
  assign n629 = ~n24 & n571 ;
  assign n630 = n438 & n629 ;
  assign n631 = ~n628 & ~n630 ;
  assign n632 = n227 & ~n631 ;
  assign n633 = ~x9 & x14 ;
  assign n634 = n105 & n633 ;
  assign n635 = n89 & n513 ;
  assign n636 = n634 & n635 ;
  assign n637 = ~n632 & ~n636 ;
  assign n638 = n65 & ~n637 ;
  assign n639 = ~x9 & n226 ;
  assign n640 = n366 & n639 ;
  assign n641 = ~x11 & n530 ;
  assign n642 = ~n105 & ~n240 ;
  assign n643 = x9 & ~n642 ;
  assign n644 = x11 & ~n145 ;
  assign n645 = ~x9 & ~n644 ;
  assign n646 = ~n643 & ~n645 ;
  assign n647 = x14 & ~n646 ;
  assign n648 = ~n641 & ~n647 ;
  assign n649 = n308 & ~n648 ;
  assign n650 = ~x3 & x13 ;
  assign n651 = n517 & n650 ;
  assign n652 = x3 & x14 ;
  assign n653 = n645 & n652 ;
  assign n654 = ~n651 & ~n653 ;
  assign n655 = n180 & ~n654 ;
  assign n656 = ~x9 & ~x14 ;
  assign n657 = ~x13 & n656 ;
  assign n658 = ~x2 & ~n531 ;
  assign n659 = x3 & ~x11 ;
  assign n660 = ~x4 & n659 ;
  assign n661 = ~n658 & n660 ;
  assign n662 = ~n657 & n661 ;
  assign n663 = ~n655 & ~n662 ;
  assign n664 = ~n649 & n663 ;
  assign n665 = ~n640 & n664 ;
  assign n666 = n306 & ~n665 ;
  assign n667 = n623 ^ n26 ;
  assign n668 = ~x2 & x9 ;
  assign n669 = ~x5 & n668 ;
  assign n670 = n669 ^ n667 ;
  assign n671 = n670 ^ n623 ;
  assign n672 = n671 ^ n670 ;
  assign n673 = x13 & ~x14 ;
  assign n674 = n639 & ~n673 ;
  assign n675 = n674 ^ n670 ;
  assign n676 = n675 ^ n667 ;
  assign n677 = n672 & ~n676 ;
  assign n678 = n677 ^ n674 ;
  assign n679 = ~x2 & x15 ;
  assign n680 = n530 & n679 ;
  assign n681 = ~n674 & ~n680 ;
  assign n682 = n681 ^ n667 ;
  assign n683 = ~n678 & ~n682 ;
  assign n684 = n683 ^ n681 ;
  assign n685 = ~n667 & n684 ;
  assign n686 = n685 ^ n677 ;
  assign n687 = n686 ^ n26 ;
  assign n688 = n687 ^ n674 ;
  assign n689 = n558 & ~n688 ;
  assign n690 = ~x1 & x14 ;
  assign n691 = ~x0 & n690 ;
  assign n692 = ~n639 & ~n680 ;
  assign n693 = n308 & ~n692 ;
  assign n694 = n691 & n693 ;
  assign n695 = ~n689 & ~n694 ;
  assign n696 = n260 & n526 ;
  assign n697 = n179 & n696 ;
  assign n698 = x13 & n517 ;
  assign n699 = ~n645 & ~n698 ;
  assign n700 = x1 & x14 ;
  assign n701 = n300 & n700 ;
  assign n702 = ~x1 & n65 ;
  assign n703 = n517 & n702 ;
  assign n704 = n39 & n703 ;
  assign n705 = ~n701 & ~n704 ;
  assign n706 = ~n699 & ~n705 ;
  assign n707 = ~x0 & n706 ;
  assign n708 = ~n697 & ~n707 ;
  assign n709 = n695 & n708 ;
  assign n710 = ~n666 & n709 ;
  assign n711 = x8 & ~n710 ;
  assign n712 = x2 & x5 ;
  assign n713 = ~x9 & n712 ;
  assign n714 = n328 & n713 ;
  assign n715 = ~x4 & n714 ;
  assign n716 = n306 & n431 ;
  assign n717 = n715 & n716 ;
  assign n718 = x13 & x14 ;
  assign n719 = x15 & n718 ;
  assign n720 = x5 & ~x8 ;
  assign n721 = ~x9 & n720 ;
  assign n722 = ~x4 & n721 ;
  assign n723 = n719 & n722 ;
  assign n724 = n69 & n723 ;
  assign n725 = ~n717 & ~n724 ;
  assign n726 = n178 & n311 ;
  assign n727 = ~x0 & x13 ;
  assign n728 = x5 & n727 ;
  assign n729 = n726 & n728 ;
  assign n730 = n105 & n311 ;
  assign n731 = n159 & n195 ;
  assign n732 = n730 & n731 ;
  assign n733 = ~n729 & ~n732 ;
  assign n734 = n266 & ~n733 ;
  assign n735 = n725 & ~n734 ;
  assign n736 = ~n711 & n735 ;
  assign n737 = ~n638 & n736 ;
  assign n738 = n622 & ~n737 ;
  assign n739 = ~x4 & ~x5 ;
  assign n740 = ~x0 & x2 ;
  assign n741 = ~n20 & ~n740 ;
  assign n742 = n348 & ~n741 ;
  assign n743 = x10 & ~n24 ;
  assign n744 = n554 & n743 ;
  assign n745 = n742 & n744 ;
  assign n746 = ~x11 & n442 ;
  assign n747 = n718 & n746 ;
  assign n748 = ~x1 & ~x11 ;
  assign n749 = ~n197 & ~n748 ;
  assign n750 = ~n110 & ~n652 ;
  assign n751 = n749 & ~n750 ;
  assign n752 = ~n57 & n751 ;
  assign n753 = ~n747 & ~n752 ;
  assign n754 = n371 & n668 ;
  assign n755 = ~n753 & n754 ;
  assign n756 = ~n745 & ~n755 ;
  assign n757 = x2 & x9 ;
  assign n758 = ~x10 & n306 ;
  assign n759 = ~x13 & n623 ;
  assign n760 = ~n383 & ~n759 ;
  assign n761 = n758 & ~n760 ;
  assign n762 = x0 & x11 ;
  assign n763 = ~x1 & n762 ;
  assign n764 = n60 & ~n126 ;
  assign n765 = n642 & n764 ;
  assign n766 = ~n763 & ~n765 ;
  assign n767 = n529 & ~n766 ;
  assign n768 = ~x14 & n240 ;
  assign n769 = n348 & n489 ;
  assign n770 = ~n768 & n769 ;
  assign n771 = ~n767 & ~n770 ;
  assign n772 = ~n761 & n771 ;
  assign n773 = n757 & ~n772 ;
  assign n774 = n756 & ~n773 ;
  assign n775 = x8 & ~n774 ;
  assign n776 = x0 & ~n467 ;
  assign n777 = x2 & n776 ;
  assign n778 = ~x2 & ~x8 ;
  assign n779 = x10 & x14 ;
  assign n780 = n274 & n779 ;
  assign n781 = n778 & n780 ;
  assign n782 = ~n777 & ~n781 ;
  assign n783 = n698 & ~n782 ;
  assign n784 = ~x2 & x10 ;
  assign n785 = ~x9 & n784 ;
  assign n786 = x8 & x14 ;
  assign n787 = ~x0 & ~x11 ;
  assign n788 = ~x13 & n787 ;
  assign n789 = n786 & n788 ;
  assign n790 = n785 & n789 ;
  assign n791 = ~n783 & ~n790 ;
  assign n792 = ~n56 & ~n791 ;
  assign n793 = ~n775 & ~n792 ;
  assign n794 = n739 & ~n793 ;
  assign n795 = x4 & x5 ;
  assign n796 = x11 & ~n467 ;
  assign n797 = n66 & n796 ;
  assign n798 = x0 & ~x8 ;
  assign n799 = ~x10 & n798 ;
  assign n800 = n462 & n799 ;
  assign n801 = ~n797 & ~n800 ;
  assign n802 = x3 & n757 ;
  assign n803 = ~n801 & n802 ;
  assign n804 = ~x0 & n562 ;
  assign n805 = n744 & n804 ;
  assign n806 = x11 & n776 ;
  assign n807 = ~n19 & n806 ;
  assign n808 = ~n563 & ~n807 ;
  assign n809 = x9 & ~n768 ;
  assign n810 = ~n808 & n809 ;
  assign n811 = ~n805 & ~n810 ;
  assign n812 = n262 & ~n811 ;
  assign n813 = ~n803 & ~n812 ;
  assign n814 = n795 & ~n813 ;
  assign n815 = ~x4 & n463 ;
  assign n816 = n301 & n815 ;
  assign n817 = x0 & x9 ;
  assign n818 = x11 & n817 ;
  assign n819 = ~n595 & ~n818 ;
  assign n820 = n816 & ~n819 ;
  assign n821 = n19 & n820 ;
  assign n822 = ~n814 & ~n821 ;
  assign n823 = ~n794 & n822 ;
  assign n824 = ~n738 & n823 ;
  assign n825 = x12 & ~n824 ;
  assign n826 = x2 & n348 ;
  assign n827 = x7 & x10 ;
  assign n828 = ~x12 & ~x13 ;
  assign n829 = n517 & n828 ;
  assign n830 = x0 & ~n346 ;
  assign n831 = ~n829 & ~n830 ;
  assign n832 = n365 & ~n831 ;
  assign n833 = n554 & n828 ;
  assign n834 = n90 & n833 ;
  assign n835 = ~n832 & ~n834 ;
  assign n836 = n827 & ~n835 ;
  assign n837 = n826 & n836 ;
  assign n838 = ~n825 & ~n837 ;
  assign n839 = ~n621 & n838 ;
  assign n840 = ~n362 & n839 ;
  assign n841 = ~n343 & n840 ;
  assign n842 = ~x6 & ~n841 ;
  assign n843 = ~x5 & x6 ;
  assign n844 = ~x4 & n843 ;
  assign n845 = ~x10 & ~x11 ;
  assign n846 = ~x3 & x12 ;
  assign n847 = n845 & n846 ;
  assign n848 = x8 & n757 ;
  assign n849 = n66 & n848 ;
  assign n850 = ~n111 & ~n112 ;
  assign n851 = ~x9 & n141 ;
  assign n852 = ~x1 & n668 ;
  assign n853 = ~n851 & ~n852 ;
  assign n854 = x0 & ~n853 ;
  assign n855 = ~n850 & n854 ;
  assign n856 = ~n849 & ~n855 ;
  assign n857 = n847 & ~n856 ;
  assign n858 = x7 & ~x9 ;
  assign n859 = n240 & n858 ;
  assign n860 = n332 & n859 ;
  assign n861 = n776 & n860 ;
  assign n1002 = ~x0 & x7 ;
  assign n1003 = ~x2 & n463 ;
  assign n1004 = n240 & n1003 ;
  assign n1005 = n370 & n1004 ;
  assign n1006 = ~n415 & ~n503 ;
  assign n1007 = ~x1 & n784 ;
  assign n1008 = ~n265 & n1007 ;
  assign n1009 = ~n1006 & n1008 ;
  assign n1010 = x10 & ~x11 ;
  assign n863 = ~x13 & ~x15 ;
  assign n864 = n396 & ~n863 ;
  assign n865 = ~x8 & n864 ;
  assign n1011 = n214 & ~n530 ;
  assign n1012 = ~n865 & ~n1011 ;
  assign n1013 = n1010 & ~n1012 ;
  assign n1014 = n265 & n524 ;
  assign n1015 = n28 & n1014 ;
  assign n1016 = ~x9 & ~n19 ;
  assign n1017 = n456 & n1016 ;
  assign n1018 = n471 & n1017 ;
  assign n1019 = ~n1015 & ~n1018 ;
  assign n1020 = ~n1013 & n1019 ;
  assign n1021 = x2 & ~n1020 ;
  assign n1022 = ~n1009 & ~n1021 ;
  assign n1023 = ~n1005 & n1022 ;
  assign n1024 = n1002 & ~n1023 ;
  assign n1025 = ~x7 & x9 ;
  assign n1026 = ~x1 & n1025 ;
  assign n1027 = ~n393 & ~n1026 ;
  assign n1028 = ~n748 & ~n1027 ;
  assign n1029 = n463 & n1028 ;
  assign n1030 = x9 & ~x10 ;
  assign n1031 = ~n104 & ~n1030 ;
  assign n1032 = ~x15 & ~n473 ;
  assign n1033 = ~n1031 & ~n1032 ;
  assign n1034 = x1 & x7 ;
  assign n1035 = n406 & n1034 ;
  assign n1036 = n1033 & n1035 ;
  assign n1037 = ~n105 & ~n418 ;
  assign n900 = ~x1 & x10 ;
  assign n1038 = ~n404 & ~n503 ;
  assign n1039 = n900 & ~n1038 ;
  assign n1040 = ~n1037 & n1039 ;
  assign n1041 = ~n1036 & ~n1040 ;
  assign n869 = ~n248 & ~n392 ;
  assign n870 = ~x9 & ~x13 ;
  assign n871 = ~n473 & ~n870 ;
  assign n872 = ~n869 & ~n871 ;
  assign n1042 = ~x1 & x7 ;
  assign n1043 = n872 & n1042 ;
  assign n1044 = x8 & n1043 ;
  assign n1045 = n1041 & ~n1044 ;
  assign n1046 = ~n1029 & n1045 ;
  assign n1047 = n20 & ~n1046 ;
  assign n995 = x10 & n58 ;
  assign n996 = n392 & n995 ;
  assign n1048 = ~x7 & n282 ;
  assign n1049 = n996 & n1048 ;
  assign n1050 = x7 & ~x11 ;
  assign n1051 = n430 & n1050 ;
  assign n1052 = n18 & n1051 ;
  assign n1053 = n332 & n1052 ;
  assign n1054 = ~n1049 & ~n1053 ;
  assign n1055 = ~n1047 & n1054 ;
  assign n1056 = ~n1024 & n1055 ;
  assign n862 = x2 & x7 ;
  assign n866 = x0 & ~x10 ;
  assign n867 = n865 & n866 ;
  assign n868 = ~n419 & n867 ;
  assign n873 = n804 & n872 ;
  assign n874 = x0 & x13 ;
  assign n875 = ~x10 & n874 ;
  assign n876 = n215 & n875 ;
  assign n877 = n66 & n104 ;
  assign n878 = ~n151 & ~n431 ;
  assign n879 = n877 & ~n878 ;
  assign n880 = ~n876 & ~n879 ;
  assign n881 = ~n873 & n880 ;
  assign n882 = ~n868 & n881 ;
  assign n883 = n862 & ~n882 ;
  assign n884 = x0 & x7 ;
  assign n885 = ~x2 & ~x9 ;
  assign n886 = n463 ^ n19 ;
  assign n887 = n886 ^ n463 ;
  assign n888 = ~x10 & x13 ;
  assign n889 = x10 & ~x13 ;
  assign n890 = ~n888 & ~n889 ;
  assign n891 = x1 & n890 ;
  assign n892 = n415 & ~n453 ;
  assign n893 = ~n891 & n892 ;
  assign n894 = n893 ^ n463 ;
  assign n895 = ~n887 & n894 ;
  assign n896 = n895 ^ n463 ;
  assign n897 = n885 & n896 ;
  assign n898 = n884 & n897 ;
  assign n899 = n568 & n727 ;
  assign n901 = n900 ^ n758 ;
  assign n902 = n900 ^ x13 ;
  assign n903 = n902 ^ n901 ;
  assign n904 = n798 ^ x8 ;
  assign n905 = ~x13 & n904 ;
  assign n906 = n905 ^ x8 ;
  assign n907 = n903 & ~n906 ;
  assign n908 = n907 ^ n905 ;
  assign n909 = n908 ^ x8 ;
  assign n910 = n909 ^ x13 ;
  assign n911 = n901 & n910 ;
  assign n912 = n911 ^ n758 ;
  assign n913 = ~n899 & ~n912 ;
  assign n914 = n554 & ~n913 ;
  assign n915 = x2 & n914 ;
  assign n916 = ~n898 & ~n915 ;
  assign n917 = ~n883 & n916 ;
  assign n918 = x10 ^ x8 ;
  assign n919 = ~x2 & x7 ;
  assign n920 = ~x0 & n919 ;
  assign n921 = x15 ^ x10 ;
  assign n922 = n918 & n921 ;
  assign n923 = n922 ^ x10 ;
  assign n924 = n920 & n923 ;
  assign n925 = n924 ^ n918 ;
  assign n926 = n58 ^ x8 ;
  assign n927 = n926 ^ n58 ;
  assign n928 = ~x0 & ~x2 ;
  assign n929 = ~n58 & ~n928 ;
  assign n930 = n929 ^ n58 ;
  assign n931 = n927 & n930 ;
  assign n932 = n931 ^ n58 ;
  assign n933 = n932 ^ n918 ;
  assign n934 = ~n925 & n933 ;
  assign n935 = n934 ^ n931 ;
  assign n936 = n935 ^ n58 ;
  assign n937 = n936 ^ n924 ;
  assign n938 = n918 & ~n937 ;
  assign n939 = n938 ^ n918 ;
  assign n940 = n939 ^ n924 ;
  assign n941 = n105 & n940 ;
  assign n942 = ~x11 & n465 ;
  assign n943 = n145 & n919 ;
  assign n944 = ~n176 & ~n943 ;
  assign n945 = n942 & ~n944 ;
  assign n946 = x2 & ~x10 ;
  assign n947 = ~n784 & ~n946 ;
  assign n948 = ~x7 & x8 ;
  assign n949 = n248 & ~n466 ;
  assign n950 = ~n948 & n949 ;
  assign n951 = ~n947 & n950 ;
  assign n952 = ~n945 & ~n951 ;
  assign n953 = x0 & ~n952 ;
  assign n954 = x10 & ~n928 ;
  assign n955 = x7 & x13 ;
  assign n956 = ~x8 & n955 ;
  assign n957 = ~n231 & ~n956 ;
  assign n958 = n954 & ~n957 ;
  assign n959 = ~n58 & n958 ;
  assign n960 = ~n953 & ~n959 ;
  assign n961 = ~n941 & n960 ;
  assign n962 = n395 & ~n961 ;
  assign n963 = n917 & ~n962 ;
  assign n964 = ~x2 & ~x13 ;
  assign n965 = x10 & n230 ;
  assign n966 = n964 & n965 ;
  assign n967 = n431 & n946 ;
  assign n968 = ~n966 & ~n967 ;
  assign n969 = n884 & ~n968 ;
  assign n970 = n112 ^ x11 ;
  assign n971 = n970 ^ n112 ;
  assign n972 = n114 & ~n971 ;
  assign n973 = n972 ^ n112 ;
  assign n974 = x13 & n973 ;
  assign n975 = n974 ^ n112 ;
  assign n976 = n489 & n975 ;
  assign n977 = x11 & n175 ;
  assign n978 = x0 & ~x11 ;
  assign n979 = n430 & n978 ;
  assign n980 = ~n977 & ~n979 ;
  assign n981 = ~x7 & x10 ;
  assign n982 = x2 & n981 ;
  assign n983 = n511 & n919 ;
  assign n984 = ~n982 & ~n983 ;
  assign n985 = ~n980 & ~n984 ;
  assign n986 = x13 & ~x15 ;
  assign n987 = x7 & n471 ;
  assign n988 = ~x0 & n198 ;
  assign n989 = n987 & n988 ;
  assign n990 = ~n986 & n989 ;
  assign n991 = ~n985 & ~n990 ;
  assign n992 = ~n976 & n991 ;
  assign n993 = ~n969 & n992 ;
  assign n994 = n370 & ~n993 ;
  assign n997 = x7 & ~x8 ;
  assign n998 = n996 & n997 ;
  assign n999 = x9 & n998 ;
  assign n1000 = ~n994 & ~n999 ;
  assign n1001 = n963 & n1000 ;
  assign n1057 = n1056 ^ n1001 ;
  assign n1058 = n1057 ^ n1001 ;
  assign n1059 = x2 & n434 ;
  assign n1060 = x1 & ~x10 ;
  assign n1061 = ~n900 & ~n1060 ;
  assign n1062 = ~x10 & n248 ;
  assign n1063 = n948 & n1062 ;
  assign n1064 = ~n1051 & ~n1063 ;
  assign n1065 = ~n1061 & ~n1064 ;
  assign n1066 = ~n419 & ~n863 ;
  assign n1067 = n1066 ^ n105 ;
  assign n1068 = n1067 ^ n105 ;
  assign n1069 = n105 ^ x7 ;
  assign n1070 = n1069 ^ n105 ;
  assign n1071 = n1068 & n1070 ;
  assign n1072 = n1071 ^ n105 ;
  assign n1073 = ~x8 & n1072 ;
  assign n1074 = n1073 ^ n105 ;
  assign n1075 = n453 & n1074 ;
  assign n1076 = ~n1065 & ~n1075 ;
  assign n1077 = n1059 & ~n1076 ;
  assign n1078 = ~x0 & n463 ;
  assign n1079 = n392 & ~n853 ;
  assign n1080 = n1078 & n1079 ;
  assign n1081 = ~n1077 & ~n1080 ;
  assign n1082 = n1081 ^ n1001 ;
  assign n1083 = n1082 ^ n1001 ;
  assign n1084 = n1058 & n1083 ;
  assign n1085 = n1084 ^ n1001 ;
  assign n1086 = x3 & n1085 ;
  assign n1087 = n1086 ^ n1001 ;
  assign n1088 = ~n861 & n1087 ;
  assign n1089 = ~x12 & ~n1088 ;
  assign n1090 = n25 & n141 ;
  assign n1091 = n74 & n224 ;
  assign n1092 = ~n1090 & ~n1091 ;
  assign n1093 = n393 & ~n1092 ;
  assign n1094 = ~n467 & n1093 ;
  assign n1095 = ~x2 & x12 ;
  assign n1096 = x15 ^ x11 ;
  assign n1097 = x11 ^ x0 ;
  assign n1098 = n1096 & n1097 ;
  assign n1099 = n1098 ^ x11 ;
  assign n1100 = n1060 & n1099 ;
  assign n1101 = ~n491 & ~n1100 ;
  assign n1102 = x13 & n162 ;
  assign n1103 = ~n1101 & n1102 ;
  assign n1104 = ~x11 & n866 ;
  assign n1105 = n66 & n473 ;
  assign n1106 = ~n1104 & ~n1105 ;
  assign n1107 = n124 & ~n1106 ;
  assign n1108 = ~x8 & n371 ;
  assign n1109 = n442 & n1108 ;
  assign n1110 = ~n1107 & ~n1109 ;
  assign n1111 = ~n1103 & n1110 ;
  assign n1112 = ~x9 & ~n1111 ;
  assign n1113 = x0 & ~x13 ;
  assign n1114 = ~x11 & n1113 ;
  assign n1115 = n568 & n1114 ;
  assign n1116 = ~n395 & ~n1115 ;
  assign n1117 = x3 & ~x8 ;
  assign n1118 = n145 & n381 ;
  assign n1119 = ~n525 & ~n978 ;
  assign n1120 = ~n1118 & n1119 ;
  assign n1121 = n1117 & ~n1120 ;
  assign n1122 = ~n1116 & n1121 ;
  assign n1123 = ~x13 & n263 ;
  assign n1124 = ~x1 & n471 ;
  assign n1125 = ~x1 & ~n511 ;
  assign n1126 = n787 & ~n1125 ;
  assign n1127 = ~n1124 & ~n1126 ;
  assign n1128 = n1123 & ~n1127 ;
  assign n1129 = x3 & n1128 ;
  assign n1130 = ~n1122 & ~n1129 ;
  assign n1131 = n438 & n888 ;
  assign n1132 = n175 & n1131 ;
  assign n1133 = n55 & n1132 ;
  assign n1134 = x10 & ~n418 ;
  assign n1135 = n763 & ~n1134 ;
  assign n1136 = ~n489 & ~n866 ;
  assign n1137 = x1 & ~n978 ;
  assign n1138 = ~n1136 & n1137 ;
  assign n1139 = ~n105 & n1138 ;
  assign n1140 = ~n1135 & ~n1139 ;
  assign n1141 = n284 & ~n1140 ;
  assign n1142 = ~n1133 & ~n1141 ;
  assign n1143 = n1130 & n1142 ;
  assign n1144 = ~n1112 & n1143 ;
  assign n1145 = n1095 & ~n1144 ;
  assign n1146 = x2 & x12 ;
  assign n1147 = n214 & n346 ;
  assign n1148 = n396 & ~n406 ;
  assign n1149 = x11 ^ x3 ;
  assign n1150 = n1149 ^ x13 ;
  assign n1151 = x13 ^ x11 ;
  assign n1152 = n1151 ^ n1148 ;
  assign n1153 = n1150 & n1152 ;
  assign n1154 = n1153 ^ x11 ;
  assign n1155 = x11 & n263 ;
  assign n1156 = n1155 ^ n1148 ;
  assign n1157 = n1154 & ~n1156 ;
  assign n1158 = n1157 ^ n1155 ;
  assign n1159 = ~n1148 & n1158 ;
  assign n1160 = n1159 ^ n1153 ;
  assign n1161 = n1160 ^ x11 ;
  assign n1162 = ~n1147 & ~n1161 ;
  assign n1163 = n381 & ~n1162 ;
  assign n1164 = n405 & n787 ;
  assign n1165 = ~x10 & n762 ;
  assign n1166 = ~x3 & n1165 ;
  assign n1167 = ~n1164 & ~n1166 ;
  assign n1168 = n28 & ~n1167 ;
  assign n1169 = ~x1 & ~x9 ;
  assign n1170 = ~x0 & n529 ;
  assign n1171 = n1169 & n1170 ;
  assign n1172 = x0 & ~n38 ;
  assign n1173 = ~n524 & ~n762 ;
  assign n1174 = ~x13 & ~n405 ;
  assign n1175 = ~n1173 & n1174 ;
  assign n1176 = ~n1172 & n1175 ;
  assign n1177 = ~n1171 & ~n1176 ;
  assign n1178 = n462 & n492 ;
  assign n1179 = ~x0 & n1178 ;
  assign n1180 = n748 & ~n1136 ;
  assign n1181 = n1180 ^ x9 ;
  assign n1182 = n1181 ^ n1180 ;
  assign n1183 = n1182 ^ n1179 ;
  assign n1184 = n1124 ^ x3 ;
  assign n1185 = ~x3 & ~n1184 ;
  assign n1186 = n1185 ^ n1180 ;
  assign n1187 = n1186 ^ x3 ;
  assign n1188 = ~n1183 & ~n1187 ;
  assign n1189 = n1188 ^ n1185 ;
  assign n1190 = n1189 ^ x3 ;
  assign n1191 = ~n1179 & ~n1190 ;
  assign n1192 = n1191 ^ n1179 ;
  assign n1193 = n1177 & ~n1192 ;
  assign n1194 = ~n1168 & n1193 ;
  assign n1195 = ~x8 & ~n1194 ;
  assign n1196 = ~n1163 & ~n1195 ;
  assign n1197 = n1146 & ~n1196 ;
  assign n1198 = ~x11 & n1030 ;
  assign n1199 = n333 & n430 ;
  assign n1200 = n1198 & n1199 ;
  assign n1201 = ~x9 & n105 ;
  assign n1202 = ~x3 & ~x10 ;
  assign n1203 = n740 & n1202 ;
  assign n1204 = n1201 & n1203 ;
  assign n1205 = n214 & n1204 ;
  assign n1206 = ~n1200 & ~n1205 ;
  assign n1207 = ~n1197 & n1206 ;
  assign n1208 = ~n1145 & n1207 ;
  assign n1209 = ~n1094 & n1208 ;
  assign n1210 = x7 & ~n1209 ;
  assign n1211 = ~n1089 & ~n1210 ;
  assign n1212 = ~n857 & n1211 ;
  assign n1213 = x14 & ~n1212 ;
  assign n1214 = x12 & x13 ;
  assign n1215 = n517 & n1214 ;
  assign n1216 = n988 & n1215 ;
  assign n1217 = x0 & x8 ;
  assign n1218 = x12 ^ x2 ;
  assign n1219 = x12 ^ x9 ;
  assign n1220 = n1219 ^ x9 ;
  assign n1221 = n698 ^ x9 ;
  assign n1222 = ~n1220 & ~n1221 ;
  assign n1223 = n1222 ^ x9 ;
  assign n1224 = ~n1218 & ~n1223 ;
  assign n1225 = n1217 & n1224 ;
  assign n1226 = ~x11 & x12 ;
  assign n1227 = ~x14 & n145 ;
  assign n1228 = x9 ^ x2 ;
  assign n1229 = n1227 & n1228 ;
  assign n1230 = n1226 & n1229 ;
  assign n1231 = n175 & n1230 ;
  assign n1232 = ~n1225 & ~n1231 ;
  assign n1233 = ~x8 & x12 ;
  assign n1234 = n105 & n1233 ;
  assign n1235 = n58 & n1234 ;
  assign n1236 = n1232 & ~n1235 ;
  assign n1237 = x1 & ~n1236 ;
  assign n1238 = ~n1216 & ~n1237 ;
  assign n1239 = n1202 & ~n1238 ;
  assign n1250 = x8 & x12 ;
  assign n1264 = ~x8 & x11 ;
  assign n1265 = x13 & n1264 ;
  assign n1281 = ~n1250 & ~n1265 ;
  assign n1282 = ~x12 & x14 ;
  assign n1283 = ~x12 & ~x15 ;
  assign n1284 = ~n1282 & ~n1283 ;
  assign n1285 = n1169 & n1284 ;
  assign n1286 = ~n1281 & n1285 ;
  assign n1287 = ~x1 & n263 ;
  assign n1270 = ~x14 & x15 ;
  assign n1271 = n828 & n1270 ;
  assign n1288 = ~x11 & ~n1271 ;
  assign n1289 = n1287 & ~n1288 ;
  assign n1290 = n346 & n1270 ;
  assign n1291 = n240 & ~n1290 ;
  assign n1292 = n1291 ^ x12 ;
  assign n1293 = n1292 ^ n1291 ;
  assign n1294 = n1293 ^ n227 ;
  assign n1295 = ~n76 & ~n863 ;
  assign n1296 = n554 ^ n227 ;
  assign n1297 = n1295 & ~n1296 ;
  assign n1298 = n1297 ^ n1291 ;
  assign n1299 = ~n1294 & ~n1298 ;
  assign n1300 = n1299 ^ n1297 ;
  assign n1301 = ~n227 & n1300 ;
  assign n1302 = n1301 ^ n1297 ;
  assign n1303 = n1302 ^ n1299 ;
  assign n1304 = ~n1289 & ~n1303 ;
  assign n1305 = ~n1286 & n1304 ;
  assign n1240 = ~x12 & n105 ;
  assign n1241 = x12 & x15 ;
  assign n1242 = n768 & n1241 ;
  assign n1243 = ~n1240 & ~n1242 ;
  assign n1244 = n55 & ~n1243 ;
  assign n1245 = n263 & n1244 ;
  assign n1246 = x11 & x12 ;
  assign n1247 = x13 & n1246 ;
  assign n1248 = n265 & n348 ;
  assign n1249 = n1247 & n1248 ;
  assign n1251 = n284 & n1250 ;
  assign n1252 = ~n462 & n1251 ;
  assign n1253 = n869 & n1252 ;
  assign n1254 = ~n1249 & ~n1253 ;
  assign n1255 = x12 & n263 ;
  assign n1256 = x3 & ~n240 ;
  assign n1257 = ~n105 & ~n1227 ;
  assign n1258 = n442 & ~n1257 ;
  assign n1259 = ~n1256 & ~n1258 ;
  assign n1260 = n1255 & ~n1259 ;
  assign n1261 = n1254 & ~n1260 ;
  assign n1262 = ~n1245 & n1261 ;
  assign n1306 = n1305 ^ n1262 ;
  assign n1263 = x9 & x12 ;
  assign n1266 = n418 & n748 ;
  assign n1267 = ~n1265 & ~n1266 ;
  assign n1268 = n1263 & ~n1267 ;
  assign n1269 = n396 & n1250 ;
  assign n1272 = x8 & n197 ;
  assign n1273 = n1271 & n1272 ;
  assign n1274 = ~n1269 & ~n1273 ;
  assign n1275 = n265 & n1214 ;
  assign n1276 = ~n263 & ~n1275 ;
  assign n1277 = n197 & ~n1276 ;
  assign n1278 = n1274 & ~n1277 ;
  assign n1279 = ~n1268 & n1278 ;
  assign n1280 = n1279 ^ n1262 ;
  assign n1307 = n1306 ^ n1280 ;
  assign n1308 = n1280 ^ x3 ;
  assign n1309 = n1308 ^ n1280 ;
  assign n1310 = n1307 & n1309 ;
  assign n1311 = n1310 ^ n1280 ;
  assign n1312 = x2 & n1311 ;
  assign n1313 = n1312 ^ n1262 ;
  assign n1314 = n489 & ~n1313 ;
  assign n1315 = ~x12 & n1270 ;
  assign n1316 = ~x3 & ~n1315 ;
  assign n1317 = ~n364 & ~n1095 ;
  assign n1318 = n265 & ~n1317 ;
  assign n1319 = ~n1316 & n1318 ;
  assign n1320 = n105 & n1319 ;
  assign n1321 = n198 & ~n492 ;
  assign n1322 = ~n1251 & ~n1321 ;
  assign n1323 = n264 & n1240 ;
  assign n1324 = n1322 & ~n1323 ;
  assign n1325 = ~n1320 & n1324 ;
  assign n1326 = n261 & ~n1325 ;
  assign n1327 = ~x12 & x13 ;
  assign n1328 = ~x11 & n1327 ;
  assign n1329 = n275 & n1328 ;
  assign n1330 = ~n1201 & ~n1256 ;
  assign n1331 = n1233 & ~n1330 ;
  assign n1332 = ~n1329 & ~n1331 ;
  assign n1333 = n310 & ~n1332 ;
  assign n1334 = n778 & n1215 ;
  assign n1335 = n38 & n1334 ;
  assign n1336 = ~x12 & n240 ;
  assign n1337 = n266 & ~n1336 ;
  assign n1338 = n306 & n1337 ;
  assign n1339 = ~n1335 & ~n1338 ;
  assign n1340 = ~n1333 & n1339 ;
  assign n1341 = ~n1326 & n1340 ;
  assign n1342 = n1341 ^ x10 ;
  assign n1343 = n1342 ^ n1341 ;
  assign n1344 = n1343 ^ n1314 ;
  assign n1345 = n277 & n1315 ;
  assign n1346 = x9 & n1095 ;
  assign n1347 = ~n1345 & ~n1346 ;
  assign n1348 = n227 & ~n1347 ;
  assign n1349 = ~x1 & ~x12 ;
  assign n1350 = n848 & n1349 ;
  assign n1351 = ~n1348 & ~n1350 ;
  assign n1352 = n392 & ~n1351 ;
  assign n1353 = ~x13 & n1270 ;
  assign n1354 = n852 & n1353 ;
  assign n1355 = ~n277 & ~n1354 ;
  assign n1356 = x12 & n230 ;
  assign n1357 = ~n1355 & n1356 ;
  assign n1358 = x9 & n562 ;
  assign n1359 = x1 & n1201 ;
  assign n1360 = ~n1358 & ~n1359 ;
  assign n1361 = n1095 & ~n1360 ;
  assign n1362 = ~n1357 & ~n1361 ;
  assign n1363 = x2 & x11 ;
  assign n1364 = x9 & ~x12 ;
  assign n1365 = n227 & ~n1364 ;
  assign n1366 = ~n1233 & ~n1365 ;
  assign n1367 = ~n828 & ~n1366 ;
  assign n1368 = ~n19 & n1367 ;
  assign n1369 = ~n1287 & ~n1368 ;
  assign n1370 = n1363 & ~n1369 ;
  assign n1371 = n1362 & ~n1370 ;
  assign n1372 = ~n1352 & n1371 ;
  assign n1373 = x0 & ~n1372 ;
  assign n1374 = n263 & n740 ;
  assign n1375 = n749 & n1327 ;
  assign n1376 = n1374 & n1375 ;
  assign n1377 = ~x0 & n141 ;
  assign n1378 = n503 & n1246 ;
  assign n1379 = n1377 & n1378 ;
  assign n1380 = ~x1 & n1095 ;
  assign n1381 = n105 & n1380 ;
  assign n1382 = x1 & x12 ;
  assign n1383 = n740 & n1382 ;
  assign n1384 = ~n1381 & ~n1383 ;
  assign n1385 = n263 & ~n1384 ;
  assign n1386 = ~n1379 & ~n1385 ;
  assign n1387 = ~n1376 & n1386 ;
  assign n1388 = ~n1373 & n1387 ;
  assign n1389 = n1388 ^ x3 ;
  assign n1390 = ~n1388 & ~n1389 ;
  assign n1391 = n1390 ^ n1341 ;
  assign n1392 = n1391 ^ n1388 ;
  assign n1393 = n1344 & n1392 ;
  assign n1394 = n1393 ^ n1390 ;
  assign n1395 = n1394 ^ n1388 ;
  assign n1396 = ~n1314 & ~n1395 ;
  assign n1397 = n1396 ^ n1314 ;
  assign n1398 = ~n1239 & ~n1397 ;
  assign n1399 = x7 & ~n1398 ;
  assign n1400 = x12 & n20 ;
  assign n1401 = n263 & n748 ;
  assign n1402 = n405 & n1401 ;
  assign n1403 = n1400 & n1402 ;
  assign n1404 = n1124 & n1255 ;
  assign n1405 = n462 & n1263 ;
  assign n1406 = ~n562 & ~n1405 ;
  assign n1407 = ~x8 & ~x12 ;
  assign n1408 = n395 & ~n1407 ;
  assign n1409 = ~n406 & n1408 ;
  assign n1410 = n1406 & ~n1409 ;
  assign n1411 = x10 & ~n1410 ;
  assign n1412 = ~n1404 & ~n1411 ;
  assign n1413 = n80 & ~n1412 ;
  assign n1414 = ~x11 & n1263 ;
  assign n1415 = n1090 & n1414 ;
  assign n1416 = n463 & n1415 ;
  assign n1417 = ~n1413 & ~n1416 ;
  assign n1418 = ~n1403 & n1417 ;
  assign n1419 = ~n1399 & n1418 ;
  assign n1420 = ~n1213 & n1419 ;
  assign n1421 = n844 & ~n1420 ;
  assign n1422 = ~x6 & ~x7 ;
  assign n1423 = x10 & x12 ;
  assign n1424 = x11 & n366 ;
  assign n1425 = n1424 ^ x14 ;
  assign n1426 = n1425 ^ n1424 ;
  assign n1427 = ~x5 & n312 ;
  assign n1428 = n1427 ^ n1424 ;
  assign n1429 = n1428 ^ n1424 ;
  assign n1430 = n1426 & n1429 ;
  assign n1431 = n1430 ^ n1424 ;
  assign n1432 = ~x9 & n1431 ;
  assign n1433 = n1432 ^ n1424 ;
  assign n1434 = n206 & n1433 ;
  assign n1435 = x5 & x11 ;
  assign n1436 = n312 & n1435 ;
  assign n1437 = x4 & n439 ;
  assign n1438 = ~n1436 & ~n1437 ;
  assign n1439 = n227 & ~n1438 ;
  assign n1440 = x3 & x8 ;
  assign n1441 = n1440 ^ n438 ;
  assign n1442 = n1440 ^ x1 ;
  assign n1443 = n1442 ^ n1440 ;
  assign n1444 = n1443 ^ n1441 ;
  assign n1445 = ~n1149 & ~n1440 ;
  assign n1446 = n1445 ^ x11 ;
  assign n1447 = ~n1444 & n1446 ;
  assign n1448 = n1447 ^ n1445 ;
  assign n1449 = n1448 ^ x11 ;
  assign n1450 = n1449 ^ n1440 ;
  assign n1451 = n1441 & ~n1450 ;
  assign n1452 = n1451 ^ n438 ;
  assign n1453 = n739 & n1452 ;
  assign n1454 = ~n1439 & ~n1453 ;
  assign n1455 = ~n1434 & n1454 ;
  assign n1456 = n58 & ~n1455 ;
  assign n1457 = n561 & n1147 ;
  assign n1458 = x1 & n530 ;
  assign n1459 = n196 & n1458 ;
  assign n1460 = n1264 & n1459 ;
  assign n1461 = ~n1457 & ~n1460 ;
  assign n1462 = n195 & ~n1461 ;
  assign n1463 = n328 & n498 ;
  assign n1464 = ~x3 & ~x5 ;
  assign n1465 = n334 & n1464 ;
  assign n1466 = ~n1463 & ~n1465 ;
  assign n1467 = n740 & ~n1466 ;
  assign n1468 = n151 & n652 ;
  assign n1469 = n235 & n1468 ;
  assign n1470 = ~n105 & ~n260 ;
  assign n1471 = n175 & n300 ;
  assign n1472 = ~n1470 & n1471 ;
  assign n1473 = ~n1469 & ~n1472 ;
  assign n1474 = ~n1467 & n1473 ;
  assign n1475 = n178 & ~n1474 ;
  assign n1476 = ~x0 & x4 ;
  assign n1477 = n235 & n1440 ;
  assign n1478 = x2 & x13 ;
  assign n1479 = n1478 ^ n700 ;
  assign n1480 = n1479 ^ n700 ;
  assign n1481 = n700 ^ n168 ;
  assign n1482 = n1481 ^ n700 ;
  assign n1483 = n1480 & ~n1482 ;
  assign n1484 = n1483 ^ n700 ;
  assign n1485 = ~n1464 & n1484 ;
  assign n1486 = n1485 ^ n700 ;
  assign n1487 = n1264 & n1486 ;
  assign n1488 = ~n168 & n230 ;
  assign n1489 = n141 & n1488 ;
  assign n1490 = ~n1487 & ~n1489 ;
  assign n1491 = ~n1477 & n1490 ;
  assign n1492 = n1476 & ~n1491 ;
  assign n1493 = ~n85 & ~n497 ;
  assign n1494 = x3 & x4 ;
  assign n1495 = ~x2 & n1494 ;
  assign n1496 = n1264 & n1495 ;
  assign n1497 = ~n1493 & n1496 ;
  assign n1498 = ~x1 & n1497 ;
  assign n1499 = ~x0 & ~x4 ;
  assign n1500 = n65 & n1435 ;
  assign n1501 = n1499 & n1500 ;
  assign n1502 = x8 & n1501 ;
  assign n1503 = ~n1498 & ~n1502 ;
  assign n1504 = ~n1492 & n1503 ;
  assign n1505 = ~n1475 & n1504 ;
  assign n1506 = x9 & ~n1505 ;
  assign n1507 = ~n1462 & ~n1506 ;
  assign n1508 = ~n1456 & n1507 ;
  assign n1509 = n513 & n571 ;
  assign n1510 = n75 & n376 ;
  assign n1511 = ~n1509 & ~n1510 ;
  assign n1512 = ~n267 & ~n1470 ;
  assign n1513 = n112 & n492 ;
  assign n1514 = ~x2 & x3 ;
  assign n1515 = x8 & ~x9 ;
  assign n1516 = n1514 & n1515 ;
  assign n1517 = ~n1513 & ~n1516 ;
  assign n1518 = n240 & ~n1517 ;
  assign n1519 = ~n1512 & ~n1518 ;
  assign n1520 = ~n1511 & ~n1519 ;
  assign n1521 = n247 & n352 ;
  assign n1522 = ~x4 & n365 ;
  assign n1523 = n332 & n1522 ;
  assign n1524 = ~x2 & ~x11 ;
  assign n1525 = n164 ^ x8 ;
  assign n1526 = n1525 ^ n164 ;
  assign n1527 = n164 ^ n160 ;
  assign n1528 = n1527 ^ n164 ;
  assign n1529 = n1526 & ~n1528 ;
  assign n1530 = n1529 ^ n164 ;
  assign n1531 = ~x4 & n1530 ;
  assign n1532 = n1531 ^ n164 ;
  assign n1533 = n1524 & n1532 ;
  assign n1534 = ~n1523 & ~n1533 ;
  assign n1535 = x14 & ~n1534 ;
  assign n1536 = x8 & n42 ;
  assign n1537 = n497 & n1536 ;
  assign n1538 = x4 & ~x5 ;
  assign n1539 = n205 & n1538 ;
  assign n1540 = ~n1537 & ~n1539 ;
  assign n1541 = x11 & ~n1540 ;
  assign n1542 = ~n1535 & ~n1541 ;
  assign n1543 = ~n1521 & n1542 ;
  assign n1544 = n284 & ~n1543 ;
  assign n1545 = x4 & n65 ;
  assign n1546 = n164 & n1264 ;
  assign n1547 = n1545 & n1546 ;
  assign n1548 = n346 & n712 ;
  assign n1549 = n479 & n1548 ;
  assign n1550 = ~n1547 & ~n1549 ;
  assign n1551 = ~n1544 & n1550 ;
  assign n1552 = n1551 ^ x0 ;
  assign n1553 = n1552 ^ n1551 ;
  assign n1554 = n1553 ^ n1520 ;
  assign n1555 = ~x11 & ~x14 ;
  assign n1556 = n530 & ~n1264 ;
  assign n1557 = ~n1555 & n1556 ;
  assign n1558 = n308 & n1557 ;
  assign n1559 = ~x9 & n328 ;
  assign n1560 = ~n230 & ~n1559 ;
  assign n1561 = n795 & ~n1515 ;
  assign n1562 = ~n1560 & n1561 ;
  assign n1563 = x8 & x11 ;
  assign n1564 = ~x9 & n1563 ;
  assign n1565 = x9 & x14 ;
  assign n1566 = ~x3 & n1565 ;
  assign n1567 = ~n1564 & ~n1566 ;
  assign n1568 = ~x13 & n739 ;
  assign n1569 = ~n217 & n1568 ;
  assign n1570 = ~n1567 & n1569 ;
  assign n1571 = ~n1562 & ~n1570 ;
  assign n1572 = ~n1558 & n1571 ;
  assign n1573 = ~x1 & ~n1572 ;
  assign n1574 = n246 & n1178 ;
  assign n1575 = n365 & n438 ;
  assign n1576 = ~n1546 & ~n1575 ;
  assign n1577 = x3 & ~n1576 ;
  assign n1578 = ~n1574 & ~n1577 ;
  assign n1579 = x4 & ~n1578 ;
  assign n1580 = n514 & n1155 ;
  assign n1581 = x1 & x4 ;
  assign n1582 = n292 & n698 ;
  assign n1583 = n196 & n265 ;
  assign n1584 = ~n1470 & n1583 ;
  assign n1585 = ~n1582 & ~n1584 ;
  assign n1586 = n1581 & ~n1585 ;
  assign n1587 = ~n1580 & ~n1586 ;
  assign n1588 = ~n1579 & n1587 ;
  assign n1589 = ~n1573 & n1588 ;
  assign n1590 = n1589 ^ x2 ;
  assign n1591 = ~x2 & n1590 ;
  assign n1592 = n1591 ^ n1551 ;
  assign n1593 = n1592 ^ x2 ;
  assign n1594 = ~n1554 & n1593 ;
  assign n1595 = n1594 ^ n1591 ;
  assign n1596 = n1595 ^ x2 ;
  assign n1597 = ~n1520 & ~n1596 ;
  assign n1598 = n1597 ^ n1520 ;
  assign n1599 = n1508 & ~n1598 ;
  assign n1600 = n1423 & ~n1599 ;
  assign n1601 = ~x10 & n1214 ;
  assign n1602 = n282 & n1514 ;
  assign n1603 = ~n1511 & n1602 ;
  assign n1604 = n1601 & n1603 ;
  assign n1605 = ~x12 & n263 ;
  assign n1606 = ~x5 & n195 ;
  assign n1607 = ~n1061 & n1606 ;
  assign n1608 = ~x10 & n1510 ;
  assign n1609 = ~n1607 & ~n1608 ;
  assign n1610 = n262 & ~n1609 ;
  assign n1611 = ~x0 & n561 ;
  assign n1612 = x4 ^ x1 ;
  assign n1613 = n946 & ~n1612 ;
  assign n1614 = n1611 & n1613 ;
  assign n1615 = ~n1610 & ~n1614 ;
  assign n1616 = x13 & ~n1615 ;
  assign n1617 = n164 & n740 ;
  assign n1618 = x4 & ~x10 ;
  assign n1619 = n650 & n1618 ;
  assign n1620 = n1617 & n1619 ;
  assign n1621 = ~n1616 & ~n1620 ;
  assign n1622 = n1605 & ~n1621 ;
  assign n1623 = ~x3 & n795 ;
  assign n1624 = ~x5 & n42 ;
  assign n1625 = ~n1623 & ~n1624 ;
  assign n1626 = ~n318 & ~n1625 ;
  assign n1627 = x1 & ~x12 ;
  assign n1628 = n381 & n1627 ;
  assign n1629 = n1626 & n1628 ;
  assign n1630 = ~x5 & x12 ;
  assign n1631 = ~x4 & n1630 ;
  assign n1632 = n126 & n1202 ;
  assign n1633 = n19 & n405 ;
  assign n1634 = ~n1632 & ~n1633 ;
  assign n1635 = n1631 & ~n1634 ;
  assign n1636 = n928 & n1635 ;
  assign n1637 = ~n1629 & ~n1636 ;
  assign n1638 = n263 & ~n1637 ;
  assign n1639 = ~n1622 & ~n1638 ;
  assign n1640 = n1639 ^ x8 ;
  assign n1641 = x5 & ~x12 ;
  assign n1642 = ~x9 & n163 ;
  assign n1643 = ~n947 & n1642 ;
  assign n1644 = n306 & n1643 ;
  assign n1645 = ~x1 & n58 ;
  assign n1646 = n284 & n557 ;
  assign n1647 = n1645 & n1646 ;
  assign n1648 = n18 & n74 ;
  assign n1649 = ~x10 & n141 ;
  assign n1650 = ~x9 & n1649 ;
  assign n1651 = ~n1648 & ~n1650 ;
  assign n1652 = n373 & ~n1651 ;
  assign n1653 = ~n1647 & ~n1652 ;
  assign n1654 = ~n1644 & n1653 ;
  assign n1655 = n1641 & ~n1654 ;
  assign n1656 = ~x10 & x12 ;
  assign n1657 = x10 & ~x12 ;
  assign n1658 = ~n1656 & ~n1657 ;
  assign n1659 = ~n160 & n291 ;
  assign n1660 = ~x3 & n164 ;
  assign n1661 = n740 & n1660 ;
  assign n1662 = ~n1659 & ~n1661 ;
  assign n1663 = ~n1658 & ~n1662 ;
  assign n1664 = ~x0 & n784 ;
  assign n1665 = ~x3 & ~x12 ;
  assign n1666 = n159 & n1665 ;
  assign n1667 = x3 & x12 ;
  assign n1668 = n79 & n1667 ;
  assign n1669 = ~n1666 & ~n1668 ;
  assign n1670 = n1664 & ~n1669 ;
  assign n1671 = ~x10 & ~x12 ;
  assign n1672 = x1 & n58 ;
  assign n1673 = n196 & n1672 ;
  assign n1674 = n1671 & n1673 ;
  assign n1675 = ~n1670 & ~n1674 ;
  assign n1676 = ~n1663 & n1675 ;
  assign n1677 = n530 & ~n1676 ;
  assign n1678 = ~x0 & ~x12 ;
  assign n1679 = x3 & ~x10 ;
  assign n1680 = n332 & n1679 ;
  assign n1681 = n1678 & n1680 ;
  assign n1682 = ~x0 & x12 ;
  assign n1683 = x0 & ~x12 ;
  assign n1684 = ~n1682 & ~n1683 ;
  assign n1685 = ~x2 & ~n1684 ;
  assign n1686 = ~x0 & n364 ;
  assign n1687 = ~x1 & n1686 ;
  assign n1688 = ~n1685 & ~n1687 ;
  assign n1689 = ~x3 & ~n1061 ;
  assign n1690 = ~n1688 & n1689 ;
  assign n1691 = ~n1681 & ~n1690 ;
  assign n1692 = x5 & ~x9 ;
  assign n1693 = x13 & n1692 ;
  assign n1694 = ~n1691 & n1693 ;
  assign n1695 = ~n1677 & ~n1694 ;
  assign n1696 = ~n1655 & n1695 ;
  assign n1697 = n1696 ^ x4 ;
  assign n1698 = n1697 ^ n1696 ;
  assign n1699 = n375 & n1683 ;
  assign n1700 = n180 & n568 ;
  assign n1701 = n1699 & n1700 ;
  assign n1702 = x12 & n75 ;
  assign n1703 = ~x9 & ~x12 ;
  assign n1704 = ~n1263 & ~n1703 ;
  assign n1705 = n571 & n1704 ;
  assign n1706 = ~n1702 & ~n1705 ;
  assign n1707 = n262 & ~n1706 ;
  assign n1708 = ~x2 & n1667 ;
  assign n1709 = n34 & n1708 ;
  assign n1710 = ~n1707 & ~n1709 ;
  assign n1711 = n568 & ~n1710 ;
  assign n1712 = ~n56 & n995 ;
  assign n1713 = n1703 & n1712 ;
  assign n1714 = ~x5 & n1713 ;
  assign n1715 = ~x9 & ~n1684 ;
  assign n1716 = ~x5 & n348 ;
  assign n1717 = n946 & n1716 ;
  assign n1718 = n1715 & n1717 ;
  assign n1719 = n1648 & n1702 ;
  assign n1720 = ~n1718 & ~n1719 ;
  assign n1721 = ~n1714 & n1720 ;
  assign n1722 = ~n1711 & n1721 ;
  assign n1723 = x13 & ~n1722 ;
  assign n1724 = ~n1701 & ~n1723 ;
  assign n1725 = n1724 ^ n1696 ;
  assign n1726 = ~n1698 & n1725 ;
  assign n1727 = n1726 ^ n1696 ;
  assign n1728 = n1727 ^ n1639 ;
  assign n1729 = ~n1640 & ~n1728 ;
  assign n1730 = n1729 ^ n1726 ;
  assign n1731 = n1730 ^ n1696 ;
  assign n1732 = n1731 ^ x8 ;
  assign n1733 = n1639 & n1732 ;
  assign n1734 = n1733 ^ n1639 ;
  assign n1735 = n1734 ^ n1639 ;
  assign n1736 = n1735 ^ x11 ;
  assign n1737 = n1736 ^ n1735 ;
  assign n1738 = n106 & n561 ;
  assign n1739 = x13 & n364 ;
  assign n1740 = n261 & n1739 ;
  assign n1741 = n28 & n1400 ;
  assign n1742 = ~x1 & x12 ;
  assign n1743 = ~x0 & n1742 ;
  assign n1744 = n1478 & n1743 ;
  assign n1745 = ~n1741 & ~n1744 ;
  assign n1746 = ~n1740 & n1745 ;
  assign n1747 = n1030 & ~n1746 ;
  assign n1748 = n1738 & n1747 ;
  assign n1749 = ~x2 & n1704 ;
  assign n1750 = ~n227 & ~n1287 ;
  assign n1751 = n1749 & ~n1750 ;
  assign n1752 = n851 & n1407 ;
  assign n1753 = ~n1751 & ~n1752 ;
  assign n1754 = n875 & ~n1753 ;
  assign n1755 = ~x3 & ~n1754 ;
  assign n1756 = ~x12 & n265 ;
  assign n1757 = n332 & n875 ;
  assign n1758 = ~x13 & n568 ;
  assign n1759 = n929 & n1758 ;
  assign n1760 = ~n1757 & ~n1759 ;
  assign n1761 = n1756 & ~n1760 ;
  assign n1762 = ~x10 & n20 ;
  assign n1763 = n1627 & n1762 ;
  assign n1764 = n282 & n1763 ;
  assign n1765 = n151 & n1682 ;
  assign n1766 = n74 & n1030 ;
  assign n1767 = n1765 & n1766 ;
  assign n1768 = x3 & ~n1767 ;
  assign n1769 = ~n1764 & n1768 ;
  assign n1770 = ~n1761 & n1769 ;
  assign n1771 = n795 & ~n1770 ;
  assign n1772 = ~n1755 & n1771 ;
  assign n1773 = ~n1748 & ~n1772 ;
  assign n1774 = n1773 ^ n1735 ;
  assign n1775 = ~n1737 & n1774 ;
  assign n1776 = n1775 ^ n1735 ;
  assign n1777 = ~n1604 & n1776 ;
  assign n1778 = n311 & ~n1777 ;
  assign n1779 = ~n1600 & ~n1778 ;
  assign n1780 = n556 & n779 ;
  assign n1781 = x13 & n20 ;
  assign n1782 = ~x5 & n55 ;
  assign n1783 = ~x12 & n517 ;
  assign n1784 = n1782 & n1783 ;
  assign n1785 = ~x11 & n1692 ;
  assign n1786 = n38 & n1785 ;
  assign n1787 = ~n1784 & ~n1786 ;
  assign n1788 = n1781 & ~n1787 ;
  assign n1789 = n1780 & n1788 ;
  assign n1790 = x8 ^ x0 ;
  assign n1791 = ~n55 & ~n159 ;
  assign n1792 = n1791 ^ x8 ;
  assign n1793 = n1792 ^ n1791 ;
  assign n1794 = n1793 ^ n1790 ;
  assign n1795 = ~n55 & ~n126 ;
  assign n1796 = n1795 ^ x5 ;
  assign n1797 = x5 & n1796 ;
  assign n1798 = n1797 ^ n1791 ;
  assign n1799 = n1798 ^ x5 ;
  assign n1800 = n1794 & ~n1799 ;
  assign n1801 = n1800 ^ n1797 ;
  assign n1802 = n1801 ^ x5 ;
  assign n1803 = n1790 & n1802 ;
  assign n1804 = n346 & n1803 ;
  assign n1805 = n607 & n746 ;
  assign n1806 = ~x1 & n196 ;
  assign n1807 = ~x8 & n517 ;
  assign n1808 = n1806 & n1807 ;
  assign n1809 = ~n1805 & ~n1808 ;
  assign n1810 = ~n1804 & n1809 ;
  assign n1811 = n249 & ~n1810 ;
  assign n1814 = n1424 ^ n739 ;
  assign n1815 = n1814 ^ n1424 ;
  assign n1812 = n1424 ^ n392 ;
  assign n1813 = n1812 ^ n1424 ;
  assign n1816 = n1815 ^ n1813 ;
  assign n1817 = n1424 ^ x3 ;
  assign n1818 = n1817 ^ n1424 ;
  assign n1819 = n1818 ^ n1815 ;
  assign n1820 = n1815 & n1819 ;
  assign n1821 = n1820 ^ n1815 ;
  assign n1822 = n1816 & n1821 ;
  assign n1823 = n1822 ^ n1820 ;
  assign n1824 = n1823 ^ n1424 ;
  assign n1825 = n1824 ^ n1815 ;
  assign n1826 = x1 & n1825 ;
  assign n1827 = n1826 ^ n1424 ;
  assign n1828 = n263 & n1827 ;
  assign n1829 = x0 & n1828 ;
  assign n1830 = n375 & n513 ;
  assign n1831 = ~x9 & n746 ;
  assign n1832 = ~n1830 & ~n1831 ;
  assign n1833 = n1217 & ~n1832 ;
  assign n1841 = x4 & x8 ;
  assign n1837 = ~n55 & ~n346 ;
  assign n1838 = x0 & ~n517 ;
  assign n1839 = ~n1837 & n1838 ;
  assign n1834 = ~x4 & ~n503 ;
  assign n1835 = n306 & n383 ;
  assign n1836 = ~n1834 & n1835 ;
  assign n1840 = n1839 ^ n1836 ;
  assign n1842 = n1841 ^ n1840 ;
  assign n1852 = n1842 ^ n1840 ;
  assign n1843 = ~n217 & ~n659 ;
  assign n1844 = x13 & ~n1843 ;
  assign n1845 = ~n348 & ~n1844 ;
  assign n1846 = n1845 ^ n1842 ;
  assign n1847 = n1846 ^ n1840 ;
  assign n1848 = n1842 ^ n1836 ;
  assign n1849 = n1848 ^ n1845 ;
  assign n1850 = n1849 ^ n1847 ;
  assign n1851 = n1847 & n1850 ;
  assign n1853 = n1852 ^ n1851 ;
  assign n1854 = n1853 ^ n1847 ;
  assign n1855 = ~x0 & x9 ;
  assign n1856 = n1855 ^ n1840 ;
  assign n1857 = n1851 ^ n1847 ;
  assign n1858 = n1856 & n1857 ;
  assign n1859 = n1858 ^ n1840 ;
  assign n1860 = ~n1854 & n1859 ;
  assign n1861 = n1860 ^ n1840 ;
  assign n1862 = n1861 ^ n1839 ;
  assign n1863 = n1862 ^ n1840 ;
  assign n1864 = ~n1833 & ~n1863 ;
  assign n1865 = n1864 ^ x5 ;
  assign n1866 = n1865 ^ n1864 ;
  assign n1867 = n1866 ^ n1829 ;
  assign n1868 = n346 & n1440 ;
  assign n1869 = ~x1 & n492 ;
  assign n1870 = ~n1037 & n1869 ;
  assign n1871 = ~n1401 & ~n1870 ;
  assign n1872 = ~n1868 & n1871 ;
  assign n1873 = n195 & ~n1872 ;
  assign n1874 = ~x0 & n348 ;
  assign n1875 = n106 & n641 ;
  assign n1876 = x4 & x11 ;
  assign n1877 = ~x9 & n1876 ;
  assign n1878 = ~n1875 & ~n1877 ;
  assign n1879 = n1874 & ~n1878 ;
  assign n1880 = ~x4 & ~x11 ;
  assign n1881 = n68 & n1880 ;
  assign n1882 = n562 & n1881 ;
  assign n1883 = ~n1879 & ~n1882 ;
  assign n1884 = ~n1873 & n1883 ;
  assign n1885 = n1884 ^ x14 ;
  assign n1886 = ~n1884 & ~n1885 ;
  assign n1887 = n1886 ^ n1864 ;
  assign n1888 = n1887 ^ n1884 ;
  assign n1889 = n1867 & n1888 ;
  assign n1890 = n1889 ^ n1886 ;
  assign n1891 = n1890 ^ n1884 ;
  assign n1892 = ~n1829 & ~n1891 ;
  assign n1893 = n1892 ^ n1829 ;
  assign n1894 = ~n1811 & ~n1893 ;
  assign n1895 = n946 & ~n1894 ;
  assign n1896 = ~x8 & n438 ;
  assign n1897 = n1581 & n1896 ;
  assign n1898 = ~x4 & n214 ;
  assign n1899 = n1201 & n1898 ;
  assign n1900 = ~n1897 & ~n1899 ;
  assign n1901 = n572 & ~n1900 ;
  assign n1902 = n652 & n1901 ;
  assign n1903 = ~x5 & n517 ;
  assign n1904 = n1581 & n1903 ;
  assign n1905 = ~x10 & x14 ;
  assign n1906 = ~x0 & n124 ;
  assign n1907 = n1905 & n1906 ;
  assign n1908 = n1904 & n1907 ;
  assign n1909 = ~x8 & x14 ;
  assign n1910 = n517 & n1909 ;
  assign n1911 = n1464 & n1910 ;
  assign n1912 = ~x5 & n623 ;
  assign n1913 = ~n263 & n497 ;
  assign n1914 = ~n1912 & ~n1913 ;
  assign n1915 = n1514 & ~n1914 ;
  assign n1916 = ~n555 & n1915 ;
  assign n1917 = ~n1911 & ~n1916 ;
  assign n1918 = n1581 & ~n1917 ;
  assign n1919 = n795 & n1358 ;
  assign n1920 = ~x5 & ~x9 ;
  assign n1921 = n1920 ^ x11 ;
  assign n1922 = n1921 ^ n1920 ;
  assign n1923 = n1920 ^ n526 ;
  assign n1924 = n1923 ^ n1920 ;
  assign n1925 = ~n1922 & n1924 ;
  assign n1926 = n1925 ^ n1920 ;
  assign n1927 = x4 & n1926 ;
  assign n1928 = n1927 ^ n1920 ;
  assign n1929 = n786 & n1928 ;
  assign n1930 = n19 & n1929 ;
  assign n1931 = ~n1919 & ~n1930 ;
  assign n1932 = n1514 & ~n1931 ;
  assign n1933 = n105 & n227 ;
  assign n1934 = ~n230 & ~n1933 ;
  assign n1935 = ~n1401 & ~n1692 ;
  assign n1936 = n44 & n366 ;
  assign n1937 = ~n1935 & n1936 ;
  assign n1938 = ~n1934 & n1937 ;
  assign n1939 = ~n1932 & ~n1938 ;
  assign n1940 = ~n1918 & n1939 ;
  assign n1941 = n866 & ~n1940 ;
  assign n1942 = ~n1908 & ~n1941 ;
  assign n1943 = ~n1902 & n1942 ;
  assign n1944 = ~n1895 & n1943 ;
  assign n1945 = x12 & ~n1944 ;
  assign n1946 = ~x0 & n38 ;
  assign n1947 = n499 & n1946 ;
  assign n1948 = x4 & ~x12 ;
  assign n1949 = ~x13 & n438 ;
  assign n1950 = ~x1 & n392 ;
  assign n1951 = ~n1949 & ~n1950 ;
  assign n1952 = ~x0 & n870 ;
  assign n1953 = n1951 & ~n1952 ;
  assign n1954 = ~x0 & x1 ;
  assign n1955 = ~n261 & ~n1954 ;
  assign n1956 = n168 & ~n1955 ;
  assign n1957 = ~n1953 & n1956 ;
  assign n1958 = n306 & n561 ;
  assign n1959 = n392 & n1958 ;
  assign n1960 = n163 & n261 ;
  assign n1961 = ~n438 & ~n1692 ;
  assign n1962 = n1960 & ~n1961 ;
  assign n1963 = ~n1959 & ~n1962 ;
  assign n1964 = ~n1957 & n1963 ;
  assign n1965 = n1948 & ~n1964 ;
  assign n1966 = n224 & n346 ;
  assign n1967 = ~n126 & ~n1349 ;
  assign n1968 = n739 & ~n1967 ;
  assign n1969 = n1966 & n1968 ;
  assign n1970 = ~n1965 & ~n1969 ;
  assign n1971 = ~n1947 & n1970 ;
  assign n1972 = n779 & ~n1971 ;
  assign n1973 = x11 & n18 ;
  assign n1974 = n1623 & n1973 ;
  assign n1975 = n1327 & ~n1955 ;
  assign n1976 = n1974 & n1975 ;
  assign n1977 = ~x12 & n718 ;
  assign n1978 = ~x12 & n497 ;
  assign n1979 = ~n1977 & ~n1978 ;
  assign n1980 = ~x10 & n517 ;
  assign n1981 = n68 & n1581 ;
  assign n1982 = n1980 & n1981 ;
  assign n1983 = ~n1979 & n1982 ;
  assign n1984 = ~n1976 & ~n1983 ;
  assign n1985 = ~n1972 & n1984 ;
  assign n1986 = n111 & ~n1985 ;
  assign n1987 = ~n1945 & ~n1986 ;
  assign n1988 = ~n1789 & n1987 ;
  assign n1989 = n277 & n524 ;
  assign n2007 = n106 & n1464 ;
  assign n1990 = ~x0 & n55 ;
  assign n1991 = x5 & ~x13 ;
  assign n1992 = n1841 & n1991 ;
  assign n1993 = n1990 & n1992 ;
  assign n1994 = x5 & n1494 ;
  assign n1995 = n66 & n1994 ;
  assign n1996 = ~x1 & n795 ;
  assign n1997 = ~n1427 & ~n1996 ;
  assign n1998 = n1172 & ~n1997 ;
  assign n1999 = ~n1995 & ~n1998 ;
  assign n2000 = n430 & ~n1999 ;
  assign n2001 = n45 & n227 ;
  assign n2002 = n1994 & n2001 ;
  assign n2003 = ~n2000 & ~n2002 ;
  assign n2004 = ~n1993 & n2003 ;
  assign n2008 = n2007 ^ n2004 ;
  assign n2009 = n2008 ^ n2004 ;
  assign n2005 = n2004 ^ n126 ;
  assign n2006 = n2005 ^ n2004 ;
  assign n2010 = n2009 ^ n2006 ;
  assign n2011 = n2004 ^ x0 ;
  assign n2012 = n2011 ^ n2004 ;
  assign n2013 = n2012 ^ n2009 ;
  assign n2014 = n2009 & ~n2013 ;
  assign n2015 = n2014 ^ n2009 ;
  assign n2016 = n2010 & n2015 ;
  assign n2017 = n2016 ^ n2014 ;
  assign n2018 = n2017 ^ n2004 ;
  assign n2019 = n2018 ^ n2009 ;
  assign n2020 = x12 & ~n2019 ;
  assign n2021 = n2020 ^ n2004 ;
  assign n2022 = n1989 & ~n2021 ;
  assign n2023 = ~x13 & n1657 ;
  assign n2024 = n434 & n2023 ;
  assign n2025 = n1427 & n2024 ;
  assign n2026 = n214 & n2025 ;
  assign n2027 = n739 & n1214 ;
  assign n2028 = n795 & n828 ;
  assign n2029 = ~n2027 & ~n2028 ;
  assign n2030 = x10 & ~n2029 ;
  assign n2031 = n66 & n263 ;
  assign n2032 = n2030 & n2031 ;
  assign n2033 = n265 & n795 ;
  assign n2034 = n263 & n739 ;
  assign n2035 = ~n2033 & ~n2034 ;
  assign n2036 = x12 & ~x13 ;
  assign n2037 = n489 & n2036 ;
  assign n2038 = ~n2035 & n2037 ;
  assign n2039 = ~x13 & n18 ;
  assign n2040 = n1522 & n2039 ;
  assign n2041 = n496 & n720 ;
  assign n2042 = n888 & n2041 ;
  assign n2043 = ~n2040 & ~n2042 ;
  assign n2044 = n1683 & ~n2043 ;
  assign n2045 = ~n2038 & ~n2044 ;
  assign n2048 = n2045 ^ n1601 ;
  assign n2049 = n2048 ^ n2045 ;
  assign n2046 = n2045 ^ n1606 ;
  assign n2047 = n2046 ^ n2045 ;
  assign n2050 = n2049 ^ n2047 ;
  assign n2051 = n2045 ^ n263 ;
  assign n2052 = n2051 ^ n2045 ;
  assign n2053 = n2052 ^ n2049 ;
  assign n2054 = n2049 & n2053 ;
  assign n2055 = n2054 ^ n2049 ;
  assign n2056 = n2050 & n2055 ;
  assign n2057 = n2056 ^ n2054 ;
  assign n2058 = n2057 ^ n2045 ;
  assign n2059 = n2058 ^ n2049 ;
  assign n2060 = ~x1 & ~n2059 ;
  assign n2061 = n2060 ^ n2045 ;
  assign n2062 = ~n2032 & n2061 ;
  assign n2063 = n65 & ~n2062 ;
  assign n2064 = ~x0 & n795 ;
  assign n2065 = n579 & n2064 ;
  assign n2066 = n739 & ~n1920 ;
  assign n2067 = ~n721 & ~n2066 ;
  assign n2068 = n1113 & ~n2067 ;
  assign n2069 = ~n2065 & ~n2068 ;
  assign n2070 = n262 & n900 ;
  assign n2071 = ~n2069 & n2070 ;
  assign n2072 = n1618 & n1991 ;
  assign n2073 = n1091 & n2072 ;
  assign n2074 = n263 & n2073 ;
  assign n2075 = n75 & n1581 ;
  assign n2076 = n888 & n2075 ;
  assign n2077 = n1476 & n1991 ;
  assign n2078 = n568 & n2077 ;
  assign n2079 = ~n2076 & ~n2078 ;
  assign n2080 = n264 & ~n2079 ;
  assign n2081 = ~n2074 & ~n2080 ;
  assign n2082 = ~n776 & ~n1078 ;
  assign n2083 = ~x1 & n284 ;
  assign n2084 = n1568 & n2083 ;
  assign n2085 = ~n2082 & n2084 ;
  assign n2086 = n2081 & ~n2085 ;
  assign n2087 = ~n2071 & n2086 ;
  assign n2088 = x12 & ~n2087 ;
  assign n2089 = n1606 ^ x0 ;
  assign n2090 = n2089 ^ n1606 ;
  assign n2091 = n1606 ^ n246 ;
  assign n2092 = n2091 ^ n1606 ;
  assign n2093 = ~n2090 & n2092 ;
  assign n2094 = n2093 ^ n1606 ;
  assign n2095 = ~x9 & n2094 ;
  assign n2096 = n2095 ^ n1606 ;
  assign n2097 = ~n1658 & n2096 ;
  assign n2098 = x9 & n489 ;
  assign n2099 = n1631 & n2098 ;
  assign n2100 = n434 & n465 ;
  assign n2101 = n1641 & n2100 ;
  assign n2102 = ~n2099 & ~n2101 ;
  assign n2103 = ~n2097 & n2102 ;
  assign n2104 = n19 & ~n2103 ;
  assign n2105 = n1601 & n2075 ;
  assign n2106 = n1515 & n2105 ;
  assign n2107 = ~n2104 & ~n2106 ;
  assign n2108 = n318 & ~n2107 ;
  assign n2109 = ~n2088 & ~n2108 ;
  assign n2110 = ~n2063 & n2109 ;
  assign n2111 = ~n2026 & n2110 ;
  assign n2112 = ~x11 & ~n2111 ;
  assign n2113 = ~n2022 & ~n2112 ;
  assign n2114 = n1270 & ~n2113 ;
  assign n2115 = ~x10 & n1246 ;
  assign n2116 = x11 & ~x12 ;
  assign n2117 = ~x13 & n2116 ;
  assign n2118 = ~x10 & n392 ;
  assign n2119 = ~n2117 & ~n2118 ;
  assign n2120 = x8 & ~n2119 ;
  assign n2121 = ~n2115 & ~n2120 ;
  assign n2122 = n2121 ^ n105 ;
  assign n2123 = n2122 ^ n2121 ;
  assign n2124 = n2121 ^ n1657 ;
  assign n2125 = n2124 ^ n2121 ;
  assign n2126 = n2123 & n2125 ;
  assign n2127 = n2126 ^ n2121 ;
  assign n2128 = ~x5 & ~n2127 ;
  assign n2129 = n2128 ^ n2121 ;
  assign n2130 = n633 & ~n2129 ;
  assign n2131 = n696 & n1233 ;
  assign n2132 = ~n240 & ~n1423 ;
  assign n2133 = n1692 & ~n2132 ;
  assign n2134 = x12 ^ x10 ;
  assign n2135 = n2134 ^ x12 ;
  assign n2136 = n1247 ^ x12 ;
  assign n2137 = n2135 & ~n2136 ;
  assign n2138 = n2137 ^ x12 ;
  assign n2139 = n918 & ~n2138 ;
  assign n2140 = n2139 ^ x8 ;
  assign n2141 = n2133 & n2140 ;
  assign n2142 = ~n246 & n1657 ;
  assign n2143 = ~n430 & n2142 ;
  assign n2144 = ~n231 & n2143 ;
  assign n2145 = n1565 & n2144 ;
  assign n2146 = ~n2141 & ~n2145 ;
  assign n2147 = ~n2131 & n2146 ;
  assign n2148 = ~n2130 & n2147 ;
  assign n2151 = n2148 ^ x5 ;
  assign n2152 = n2151 ^ n2148 ;
  assign n2149 = n2148 ^ x10 ;
  assign n2150 = n2149 ^ n2148 ;
  assign n2153 = n2152 ^ n2150 ;
  assign n2154 = ~x9 & x12 ;
  assign n2155 = n1563 & ~n2154 ;
  assign n2156 = n2155 ^ x14 ;
  assign n2157 = n2155 ^ x12 ;
  assign n2158 = n2157 ^ x12 ;
  assign n2159 = n1414 ^ x12 ;
  assign n2160 = ~n2158 & ~n2159 ;
  assign n2161 = n2160 ^ x12 ;
  assign n2162 = n2156 & n2161 ;
  assign n2163 = n2162 ^ x14 ;
  assign n2164 = x13 & n2163 ;
  assign n2165 = n76 & n1226 ;
  assign n2166 = ~x8 & n2165 ;
  assign n2167 = ~n2164 & ~n2166 ;
  assign n2168 = n2167 ^ n2148 ;
  assign n2169 = n2168 ^ n2148 ;
  assign n2170 = n2169 ^ n2152 ;
  assign n2171 = ~n2152 & n2170 ;
  assign n2172 = n2171 ^ n2152 ;
  assign n2173 = ~n2153 & ~n2172 ;
  assign n2174 = n2173 ^ n2171 ;
  assign n2175 = n2174 ^ n2148 ;
  assign n2176 = n2175 ^ n2152 ;
  assign n2177 = ~x4 & n2176 ;
  assign n2178 = n2177 ^ n2148 ;
  assign n2179 = ~n1092 & ~n2178 ;
  assign n2180 = ~x0 & n1246 ;
  assign n2181 = n21 & n2180 ;
  assign n2182 = ~x4 & x12 ;
  assign n2183 = ~n1948 & ~n2182 ;
  assign n2184 = n978 & ~n1494 ;
  assign n2185 = ~n2183 & n2184 ;
  assign n2186 = ~n2181 & ~n2185 ;
  assign n2187 = n411 & ~n2186 ;
  assign n2188 = n571 & n2115 ;
  assign n2189 = x4 & n2188 ;
  assign n2190 = n367 & n524 ;
  assign n2191 = n1630 & n2190 ;
  assign n2192 = ~n2189 & ~n2191 ;
  assign n2193 = ~n2187 & n2192 ;
  assign n2194 = n668 & ~n2193 ;
  assign n2195 = x10 ^ x9 ;
  assign n2196 = n2195 ^ n1246 ;
  assign n2197 = n570 ^ x9 ;
  assign n2198 = n2197 ^ n570 ;
  assign n2199 = n20 & n26 ;
  assign n2200 = n2199 ^ n570 ;
  assign n2201 = ~n2198 & n2200 ;
  assign n2202 = n2201 ^ n570 ;
  assign n2203 = n2202 ^ n2195 ;
  assign n2204 = n2196 & n2203 ;
  assign n2205 = n2204 ^ n2201 ;
  assign n2206 = n2205 ^ n570 ;
  assign n2207 = n2206 ^ n1246 ;
  assign n2208 = n2195 & n2207 ;
  assign n2209 = n2208 ^ n2195 ;
  assign n2210 = ~n2194 & ~n2209 ;
  assign n2211 = n562 & ~n2210 ;
  assign n2212 = n106 & n1414 ;
  assign n2213 = ~x11 & n263 ;
  assign n2214 = n1349 & n2213 ;
  assign n2215 = x12 ^ x11 ;
  assign n2216 = n1365 & n2215 ;
  assign n2217 = ~n2214 & ~n2216 ;
  assign n2218 = x4 & ~n2217 ;
  assign n2219 = ~n2212 & ~n2218 ;
  assign n2220 = n489 & ~n2219 ;
  assign n2221 = n471 & n1287 ;
  assign n2222 = ~x4 & n2221 ;
  assign n2223 = x12 & n2222 ;
  assign n2224 = ~x8 & ~x10 ;
  assign n2225 = n1246 & n2224 ;
  assign n2226 = x4 & n261 ;
  assign n2227 = n2225 & n2226 ;
  assign n2228 = x12 & n1954 ;
  assign n2229 = n354 & n1876 ;
  assign n2230 = n2228 & n2229 ;
  assign n2231 = ~n2227 & ~n2230 ;
  assign n2232 = ~n263 & n513 ;
  assign n2233 = n776 & n2232 ;
  assign n2234 = n1226 & n2233 ;
  assign n2235 = n2231 & ~n2234 ;
  assign n2236 = ~n2223 & n2235 ;
  assign n2237 = ~n2220 & n2236 ;
  assign n2238 = n712 & ~n2237 ;
  assign n2239 = x0 & x4 ;
  assign n2240 = ~n197 & n1657 ;
  assign n2241 = ~x4 & ~n2240 ;
  assign n2242 = n263 & ~n2241 ;
  assign n2243 = ~n2239 & ~n2242 ;
  assign n2244 = ~n227 & n2239 ;
  assign n2245 = n213 & ~n748 ;
  assign n2246 = x4 & ~n1656 ;
  assign n2247 = n2245 & ~n2246 ;
  assign n2248 = ~n2244 & n2247 ;
  assign n2249 = ~x0 & ~n1876 ;
  assign n2250 = ~n346 & ~n2249 ;
  assign n2251 = n2248 & n2250 ;
  assign n2252 = ~n2243 & n2251 ;
  assign n2253 = n175 & ~n555 ;
  assign n2254 = n1097 ^ x11 ;
  assign n2255 = n554 ^ x11 ;
  assign n2256 = ~n2254 & ~n2255 ;
  assign n2257 = n2256 ^ x11 ;
  assign n2258 = n227 & ~n2257 ;
  assign n2259 = ~n2253 & ~n2258 ;
  assign n2260 = x10 & ~n2259 ;
  assign n2261 = ~n2221 & ~n2260 ;
  assign n2262 = n795 & ~n2261 ;
  assign n2263 = n122 & n568 ;
  assign n2264 = n2034 & n2263 ;
  assign n2265 = ~n2262 & ~n2264 ;
  assign n2266 = n1095 & ~n2265 ;
  assign n2267 = ~n2252 & ~n2266 ;
  assign n2268 = ~n2238 & n2267 ;
  assign n2269 = x3 & ~n2268 ;
  assign n2270 = n366 & n720 ;
  assign n2271 = x0 & x12 ;
  assign n2272 = n141 & n2271 ;
  assign n2273 = n471 & n2272 ;
  assign n2274 = n2270 & n2273 ;
  assign n2275 = ~n2269 & ~n2274 ;
  assign n2276 = ~n2211 & n2275 ;
  assign n2277 = ~n24 & ~n2276 ;
  assign n2278 = ~n2179 & ~n2277 ;
  assign n2279 = ~x4 & x10 ;
  assign n2280 = x5 & ~x11 ;
  assign n2281 = ~n870 & ~n2280 ;
  assign n2282 = x0 & x14 ;
  assign n2283 = ~n1991 & n2282 ;
  assign n2284 = n1349 & n2283 ;
  assign n2285 = ~n2281 & n2284 ;
  assign n2286 = ~x9 & n260 ;
  assign n2287 = ~n1783 & ~n2286 ;
  assign n2288 = n34 & n126 ;
  assign n2289 = ~n2287 & n2288 ;
  assign n2290 = ~x11 & ~x12 ;
  assign n2291 = n76 & n2290 ;
  assign n2292 = ~x9 & n2291 ;
  assign n2293 = ~n329 & ~n2292 ;
  assign n2294 = n306 & ~n1920 ;
  assign n2295 = ~n2293 & n2294 ;
  assign n2296 = ~n2289 & ~n2295 ;
  assign n2297 = ~n2285 & n2296 ;
  assign n2298 = n2297 ^ n261 ;
  assign n2299 = n2298 ^ x3 ;
  assign n2309 = n2299 ^ n2298 ;
  assign n2300 = ~x5 & ~x11 ;
  assign n2301 = n828 & n1565 ;
  assign n2302 = n2300 & n2301 ;
  assign n2303 = n2302 ^ n2299 ;
  assign n2304 = n2303 ^ n2298 ;
  assign n2305 = n2299 ^ n2297 ;
  assign n2306 = n2305 ^ n2302 ;
  assign n2307 = n2306 ^ n2304 ;
  assign n2308 = ~n2304 & ~n2307 ;
  assign n2310 = n2309 ^ n2308 ;
  assign n2311 = n2310 ^ n2304 ;
  assign n2312 = n248 & n1282 ;
  assign n2313 = n2312 ^ x11 ;
  assign n2314 = ~n1692 & ~n2313 ;
  assign n2315 = n2314 ^ x11 ;
  assign n2316 = n2315 ^ n2298 ;
  assign n2317 = n2308 ^ n2304 ;
  assign n2318 = ~n2316 & ~n2317 ;
  assign n2319 = n2318 ^ n2298 ;
  assign n2320 = ~n2311 & ~n2319 ;
  assign n2321 = n2320 ^ n2298 ;
  assign n2322 = n2321 ^ n261 ;
  assign n2323 = n2322 ^ n2298 ;
  assign n2324 = n2279 & ~n2323 ;
  assign n2325 = ~n659 & ~n759 ;
  assign n2326 = x3 & ~x13 ;
  assign n2327 = ~n1955 & ~n2326 ;
  assign n2328 = ~n2325 & n2327 ;
  assign n2329 = x13 & n109 ;
  assign n2330 = ~n328 & ~n373 ;
  assign n2331 = n2329 & ~n2330 ;
  assign n2332 = ~n2328 & ~n2331 ;
  assign n2333 = n1364 & ~n2332 ;
  assign n2334 = n375 & n763 ;
  assign n2335 = ~n2333 & ~n2334 ;
  assign n2336 = n795 & ~n2335 ;
  assign n2337 = n978 & n1692 ;
  assign n2338 = x14 & ~n348 ;
  assign n2339 = n2337 & n2338 ;
  assign n2340 = ~n57 & n2339 ;
  assign n2341 = ~n19 & ~n329 ;
  assign n2342 = n68 & ~n2341 ;
  assign n2343 = ~x1 & n561 ;
  assign n2344 = x11 & n2343 ;
  assign n2345 = ~n2342 & ~n2344 ;
  assign n2346 = ~n248 & n1565 ;
  assign n2347 = ~n2345 & n2346 ;
  assign n2348 = ~n2340 & ~n2347 ;
  assign n2349 = n1948 & ~n2348 ;
  assign n2350 = n762 & n1327 ;
  assign n2351 = ~x5 & n2350 ;
  assign n2352 = n1830 & n2351 ;
  assign n2353 = ~x10 & ~n2352 ;
  assign n2354 = ~n2349 & n2353 ;
  assign n2355 = ~n2336 & n2354 ;
  assign n2356 = ~x12 & n76 ;
  assign n2357 = n439 & n2356 ;
  assign n2358 = x3 & ~x12 ;
  assign n2359 = n2286 & n2358 ;
  assign n2360 = n383 ^ x9 ;
  assign n2361 = n2360 ^ n383 ;
  assign n2362 = n76 & n1665 ;
  assign n2363 = n2362 ^ n383 ;
  assign n2364 = ~n2361 & n2363 ;
  assign n2365 = n2364 ^ n383 ;
  assign n2366 = ~n2359 & ~n2365 ;
  assign n2367 = x5 & ~n2366 ;
  assign n2368 = ~n2357 & ~n2367 ;
  assign n2369 = n66 & ~n2368 ;
  assign n2370 = ~n196 & ~n561 ;
  assign n2371 = n517 & ~n2370 ;
  assign n2372 = n39 & n2358 ;
  assign n2373 = n260 & n2372 ;
  assign n2374 = n718 & n1703 ;
  assign n2375 = n2280 & n2374 ;
  assign n2376 = ~n2373 & ~n2375 ;
  assign n2377 = ~n2371 & n2376 ;
  assign n2378 = n1954 & ~n2377 ;
  assign n2379 = n390 & ~n492 ;
  assign n2380 = n1791 & n2379 ;
  assign n2381 = ~n391 & ~n2380 ;
  assign n2382 = ~n2378 & ~n2381 ;
  assign n2383 = ~n2369 & n2382 ;
  assign n2384 = x8 & ~n2383 ;
  assign n2385 = ~n2355 & n2384 ;
  assign n2386 = ~n2324 & n2385 ;
  assign n2387 = n168 & n396 ;
  assign n2388 = n787 & n2387 ;
  assign n2389 = ~x1 & n517 ;
  assign n2390 = ~n2370 & n2389 ;
  assign n2391 = ~n2388 & ~n2390 ;
  assign n2392 = n1327 & ~n2391 ;
  assign n2393 = n1780 & n2392 ;
  assign n2394 = ~x8 & n795 ;
  assign n2395 = ~x10 & n328 ;
  assign n2396 = n57 & ~n555 ;
  assign n2397 = n2395 & n2396 ;
  assign n2398 = x10 & n197 ;
  assign n2399 = n284 & n2398 ;
  assign n2400 = ~n2397 & ~n2399 ;
  assign n2401 = n2394 & ~n2400 ;
  assign n2402 = n109 & n492 ;
  assign n2403 = n739 & n2402 ;
  assign n2404 = n348 & n1880 ;
  assign n2405 = ~n1424 & ~n2404 ;
  assign n2406 = x9 & n292 ;
  assign n2407 = ~n2405 & n2406 ;
  assign n2408 = n556 & n2083 ;
  assign n2409 = n2280 & n2408 ;
  assign n2410 = ~n2407 & ~n2409 ;
  assign n2411 = ~n2403 & n2410 ;
  assign n2412 = n779 & ~n2411 ;
  assign n2413 = ~n471 & ~n1010 ;
  assign n2414 = n2413 ^ n524 ;
  assign n2415 = x1 & ~n2414 ;
  assign n2416 = n2415 ^ n524 ;
  assign n2417 = n1994 & n2416 ;
  assign n2418 = n265 & n2417 ;
  assign n2419 = n1692 & n2224 ;
  assign n2420 = n2419 ^ n249 ;
  assign n2421 = n383 ^ x1 ;
  assign n2422 = n2421 ^ n383 ;
  assign n2423 = n1843 ^ n383 ;
  assign n2424 = n2422 & ~n2423 ;
  assign n2425 = n2424 ^ n383 ;
  assign n2426 = n2425 ^ n2419 ;
  assign n2427 = n2420 & n2426 ;
  assign n2428 = n2427 ^ n2424 ;
  assign n2429 = n2428 ^ n383 ;
  assign n2430 = n2429 ^ n249 ;
  assign n2431 = n2419 & n2430 ;
  assign n2432 = n2431 ^ n2419 ;
  assign n2433 = ~n2418 & ~n2432 ;
  assign n2434 = ~n2412 & n2433 ;
  assign n2435 = n1327 & ~n2434 ;
  assign n2436 = n418 & n690 ;
  assign n2437 = ~n1031 & n1948 ;
  assign n2438 = ~n217 & ~n1785 ;
  assign n2439 = n2437 & ~n2438 ;
  assign n2440 = n2436 & n2439 ;
  assign n2441 = ~n2435 & ~n2440 ;
  assign n2442 = ~n2401 & n2441 ;
  assign n2443 = x0 & ~n2442 ;
  assign n2444 = ~n2393 & ~n2443 ;
  assign n2445 = ~n2386 & n2444 ;
  assign n2446 = x2 & ~n2445 ;
  assign n2447 = n2278 & ~n2446 ;
  assign n2448 = ~n2114 & n2447 ;
  assign n2449 = n1988 & n2448 ;
  assign n2450 = n1779 & n2449 ;
  assign n2451 = n1422 & ~n2450 ;
  assign n2452 = ~n1421 & ~n2451 ;
  assign n2453 = ~n842 & n2452 ;
  assign n2454 = n1422 & n1515 ;
  assign n2455 = ~x11 & n779 ;
  assign n2456 = n1499 & n2455 ;
  assign n2457 = n2454 & n2456 ;
  assign n2458 = ~x0 & ~x7 ;
  assign n2459 = n260 & n354 ;
  assign n2460 = n556 & n2459 ;
  assign n2461 = ~x10 & n1563 ;
  assign n2462 = n249 & n2461 ;
  assign n2463 = n1703 & n2462 ;
  assign n2464 = ~n2460 & ~n2463 ;
  assign n2465 = n2458 & ~n2464 ;
  assign n2466 = ~x12 & ~x14 ;
  assign n2467 = ~x7 & x11 ;
  assign n2468 = ~n438 & ~n2467 ;
  assign n2469 = n489 & ~n2468 ;
  assign n2470 = ~x7 & n471 ;
  assign n2471 = ~x11 & n18 ;
  assign n2472 = ~n2470 & ~n2471 ;
  assign n2473 = x0 & ~n2472 ;
  assign n2474 = ~n1025 & n2473 ;
  assign n2475 = ~n2469 & ~n2474 ;
  assign n2476 = n1841 & ~n2475 ;
  assign n2480 = ~x7 & ~x9 ;
  assign n2481 = n463 & ~n2480 ;
  assign n2482 = n1838 & n2481 ;
  assign n2477 = ~n524 & ~n845 ;
  assign n2478 = ~x9 & n798 ;
  assign n2479 = ~n2477 & n2478 ;
  assign n2483 = n2482 ^ n2479 ;
  assign n2484 = n2483 ^ x4 ;
  assign n2491 = n2484 ^ n2483 ;
  assign n2485 = n2484 ^ n390 ;
  assign n2486 = n2485 ^ n2483 ;
  assign n2487 = n2479 ^ n390 ;
  assign n2488 = n2487 ^ n390 ;
  assign n2489 = n2488 ^ n2486 ;
  assign n2490 = n2486 & n2489 ;
  assign n2492 = n2491 ^ n2490 ;
  assign n2493 = n2492 ^ n2486 ;
  assign n2494 = n2483 ^ x7 ;
  assign n2495 = n2490 ^ n2486 ;
  assign n2496 = n2494 & n2495 ;
  assign n2497 = n2496 ^ n2483 ;
  assign n2498 = ~n2493 & n2497 ;
  assign n2499 = n2498 ^ n2483 ;
  assign n2500 = n2499 ^ n2479 ;
  assign n2501 = n2500 ^ n2483 ;
  assign n2502 = ~n2476 & ~n2501 ;
  assign n2503 = n2466 & ~n2502 ;
  assign n2504 = ~n2465 & ~n2503 ;
  assign n2505 = x6 & ~n2504 ;
  assign n2506 = ~n2457 & ~n2505 ;
  assign n2507 = n39 & ~n2506 ;
  assign n2508 = x9 & ~x14 ;
  assign n2509 = x6 & x11 ;
  assign n2510 = ~x10 & n17 ;
  assign n2511 = n1841 & n2510 ;
  assign n2512 = ~x7 & x12 ;
  assign n2513 = n1108 & ~n2512 ;
  assign n2514 = ~n2183 & n2513 ;
  assign n2515 = ~n2511 & ~n2514 ;
  assign n2516 = n2509 & ~n2515 ;
  assign n2517 = n1880 & n2271 ;
  assign n2518 = n1422 & n2517 ;
  assign n2519 = n466 & n2518 ;
  assign n2520 = ~n2516 & ~n2519 ;
  assign n2521 = n2508 & ~n2520 ;
  assign n2522 = x4 & x12 ;
  assign n2523 = n2522 ^ n2183 ;
  assign n2524 = ~x0 & ~n2523 ;
  assign n2525 = n2524 ^ n2183 ;
  assign n2526 = n2224 & ~n2525 ;
  assign n2527 = x8 & ~x12 ;
  assign n2528 = ~x0 & n2279 ;
  assign n2529 = n2527 & n2528 ;
  assign n2530 = ~n2526 & ~n2529 ;
  assign n2531 = n2286 & ~n2530 ;
  assign n2532 = n2531 ^ x7 ;
  assign n2533 = n2532 ^ n2531 ;
  assign n2534 = n2533 ^ n2521 ;
  assign n2535 = ~x4 & ~x6 ;
  assign n2536 = n2271 & n2535 ;
  assign n2537 = x6 & ~x12 ;
  assign n2538 = n1476 & n2537 ;
  assign n2539 = ~n2536 & ~n2538 ;
  assign n2540 = ~x8 & n554 ;
  assign n2541 = ~n1198 & ~n2540 ;
  assign n2542 = ~n2539 & ~n2541 ;
  assign n2543 = ~n1564 & ~n2471 ;
  assign n2544 = n2535 & ~n2543 ;
  assign n2545 = ~n1684 & n2544 ;
  assign n2546 = ~n2542 & ~n2545 ;
  assign n2547 = n2546 ^ x14 ;
  assign n2548 = ~n2546 & ~n2547 ;
  assign n2549 = n2548 ^ n2531 ;
  assign n2550 = n2549 ^ n2546 ;
  assign n2551 = n2534 & ~n2550 ;
  assign n2552 = n2551 ^ n2548 ;
  assign n2553 = n2552 ^ n2546 ;
  assign n2554 = ~n2521 & ~n2553 ;
  assign n2555 = n2554 ^ n2521 ;
  assign n2556 = n624 & n2555 ;
  assign n2557 = ~x7 & x13 ;
  assign n2558 = x7 & ~x13 ;
  assign n2559 = ~n2557 & ~n2558 ;
  assign n2560 = x10 & ~x14 ;
  assign n2561 = ~n2559 & n2560 ;
  assign n2562 = x0 & ~x6 ;
  assign n2563 = n1841 & n2562 ;
  assign n2564 = ~x12 & n438 ;
  assign n2565 = n2563 & n2564 ;
  assign n2566 = n2561 & n2565 ;
  assign n2567 = ~n2556 & ~n2566 ;
  assign n2568 = x0 & ~x14 ;
  assign n2569 = x4 & ~x7 ;
  assign n2570 = ~n299 & ~n2461 ;
  assign n2571 = n2569 & ~n2570 ;
  assign n2572 = n438 & n815 ;
  assign n2573 = ~n2571 & ~n2572 ;
  assign n2574 = n2537 & ~n2573 ;
  assign n2575 = x4 & ~x6 ;
  assign n2576 = n18 & n2575 ;
  assign n2577 = n1264 & n2512 ;
  assign n2578 = n2576 & n2577 ;
  assign n2579 = ~n2574 & ~n2578 ;
  assign n2580 = n2568 & ~n2579 ;
  assign n2581 = ~x7 & ~x8 ;
  assign n2582 = n1905 & n2581 ;
  assign n2583 = x7 & ~x14 ;
  assign n2584 = ~n1002 & ~n2583 ;
  assign n2585 = n815 & ~n2584 ;
  assign n2586 = ~n2582 & ~n2585 ;
  assign n2587 = x6 & x10 ;
  assign n2588 = n1226 & ~n2587 ;
  assign n2589 = x6 ^ x0 ;
  assign n2590 = n2589 ^ x6 ;
  assign n2591 = x6 & x14 ;
  assign n2592 = ~n779 & ~n2591 ;
  assign n2593 = n2592 ^ x6 ;
  assign n2594 = ~n2590 & n2593 ;
  assign n2595 = n2594 ^ x6 ;
  assign n2596 = n2588 & ~n2595 ;
  assign n2597 = ~n2586 & n2596 ;
  assign n2598 = ~n799 & ~n1078 ;
  assign n2599 = ~x0 & x6 ;
  assign n2600 = ~n2562 & ~n2599 ;
  assign n2601 = ~x7 & ~x11 ;
  assign n2602 = n1282 & n2601 ;
  assign n2603 = n2600 & n2602 ;
  assign n2604 = ~n2598 & n2603 ;
  assign n2605 = x12 & n762 ;
  assign n2606 = x7 & n2605 ;
  assign n2607 = ~x10 & ~x14 ;
  assign n2608 = x4 & x6 ;
  assign n2609 = n2607 & n2608 ;
  assign n2610 = n2609 ^ x14 ;
  assign n2611 = n2610 ^ n2609 ;
  assign n2612 = ~x6 & x10 ;
  assign n2613 = ~x4 & n2612 ;
  assign n2614 = n2613 ^ n2609 ;
  assign n2615 = n2614 ^ n2609 ;
  assign n2616 = n2611 & n2615 ;
  assign n2617 = n2616 ^ n2609 ;
  assign n2618 = x8 & n2617 ;
  assign n2619 = n2618 ^ n2609 ;
  assign n2620 = n2606 & n2619 ;
  assign n2621 = ~n2604 & ~n2620 ;
  assign n2622 = ~n2597 & n2621 ;
  assign n2623 = ~x9 & ~n2622 ;
  assign n2624 = ~x8 & n2608 ;
  assign n2625 = n18 & n1226 ;
  assign n2626 = n2624 & n2625 ;
  assign n2627 = n2583 & n2626 ;
  assign n2628 = ~n2623 & ~n2627 ;
  assign n2629 = ~n2580 & n2628 ;
  assign n2630 = n1991 & ~n2629 ;
  assign n2631 = x10 & n1683 ;
  assign n2632 = n2454 & n2631 ;
  assign n2633 = x0 & ~x7 ;
  assign n2634 = ~x8 & n104 ;
  assign n2635 = ~n942 & ~n2634 ;
  assign n2636 = n2633 & ~n2635 ;
  assign n2637 = x7 & x9 ;
  assign n2638 = ~x8 & n2637 ;
  assign n2639 = n524 & n2638 ;
  assign n2640 = ~n2636 & ~n2639 ;
  assign n2641 = n2537 & ~n2640 ;
  assign n2642 = n2509 & n2638 ;
  assign n2643 = n1656 & n2642 ;
  assign n2644 = ~n2641 & ~n2643 ;
  assign n2645 = ~n2632 & n2644 ;
  assign n2646 = x4 & n673 ;
  assign n2647 = ~n2645 & n2646 ;
  assign n2648 = x5 & n2647 ;
  assign n2649 = ~n2630 & ~n2648 ;
  assign n2650 = n2567 & n2649 ;
  assign n2651 = ~n2507 & n2650 ;
  assign n2652 = n1514 & ~n2651 ;
  assign n2653 = x5 & x7 ;
  assign n2654 = ~x9 & n2653 ;
  assign n2655 = ~n104 & ~n2654 ;
  assign n2656 = ~x0 & n2655 ;
  assign n2657 = ~n105 & ~n2608 ;
  assign n2658 = n739 & n1422 ;
  assign n2659 = ~n381 & ~n2658 ;
  assign n2660 = n2657 & ~n2659 ;
  assign n2661 = ~n2656 & n2660 ;
  assign n2662 = ~x9 & ~n240 ;
  assign n2663 = ~x12 & ~n371 ;
  assign n2664 = ~n1949 & n2663 ;
  assign n2665 = ~n2662 & n2664 ;
  assign n2666 = n2661 & n2665 ;
  assign n2667 = n328 & n2666 ;
  assign n2668 = ~x6 & x12 ;
  assign n2669 = ~x4 & n2668 ;
  assign n2670 = ~n110 & n1104 ;
  assign n2671 = ~n163 & ~n1679 ;
  assign n2672 = x11 & ~n557 ;
  assign n2673 = ~n2671 & n2672 ;
  assign n2674 = ~n2670 & ~n2673 ;
  assign n2675 = x9 & n2653 ;
  assign n2676 = ~x14 & n2675 ;
  assign n2677 = ~n2674 & n2676 ;
  assign n2678 = ~x7 & ~x13 ;
  assign n2679 = ~x5 & n25 ;
  assign n2680 = n2459 & n2679 ;
  assign n2681 = n2678 & n2680 ;
  assign n2682 = ~n2677 & ~n2681 ;
  assign n2683 = n2669 & ~n2682 ;
  assign n2684 = ~x6 & x7 ;
  assign n2685 = n525 & n2684 ;
  assign n2686 = x6 & x9 ;
  assign n2687 = n2118 & n2686 ;
  assign n2688 = ~n2685 & ~n2687 ;
  assign n2689 = n196 & ~n2688 ;
  assign n2690 = ~x6 & n411 ;
  assign n2691 = n240 & n2690 ;
  assign n2692 = n2637 & n2691 ;
  assign n2693 = ~x6 & ~x10 ;
  assign n2694 = n650 & n2693 ;
  assign n2695 = n329 & n2694 ;
  assign n2696 = n2480 & n2695 ;
  assign n2697 = ~n2692 & ~n2696 ;
  assign n2698 = ~n2689 & n2697 ;
  assign n2699 = n195 & ~n2698 ;
  assign n2700 = x13 & n489 ;
  assign n2701 = ~x4 & x6 ;
  assign n2702 = ~n2575 & ~n2701 ;
  assign n2703 = ~n843 & ~n2569 ;
  assign n2704 = ~n2702 & n2703 ;
  assign n2705 = n439 & n2704 ;
  assign n2706 = n2700 & n2705 ;
  assign n2707 = x5 & ~x6 ;
  assign n2708 = x7 & n2707 ;
  assign n2709 = n312 & n2708 ;
  assign n2710 = n18 & n2709 ;
  assign n2711 = ~n168 & ~n1464 ;
  assign n2712 = x6 & n2458 ;
  assign n2713 = n1618 & n2712 ;
  assign n2714 = n2711 & n2713 ;
  assign n2715 = ~n2710 & ~n2714 ;
  assign n2716 = n105 & ~n2715 ;
  assign n2717 = ~n2706 & ~n2716 ;
  assign n2718 = n870 & n2279 ;
  assign n2719 = n2708 & n2718 ;
  assign n2720 = n105 & n1030 ;
  assign n2721 = n843 & n2569 ;
  assign n2722 = n2720 & n2721 ;
  assign n2723 = ~n2719 & ~n2722 ;
  assign n2724 = x3 & ~n2723 ;
  assign n2725 = n1619 & n2684 ;
  assign n2726 = n438 & n2725 ;
  assign n2727 = ~n2724 & ~n2726 ;
  assign n2728 = x0 & ~n2727 ;
  assign n2729 = n2717 & ~n2728 ;
  assign n2730 = ~n2699 & n2729 ;
  assign n2731 = n2466 & ~n2730 ;
  assign n2732 = ~n2683 & ~n2731 ;
  assign n2733 = ~n2667 & n2732 ;
  assign n2734 = n198 & ~n2733 ;
  assign n2735 = ~x10 & ~n869 ;
  assign n2736 = ~x12 & n607 ;
  assign n2737 = n2735 & n2736 ;
  assign n2738 = ~x13 & n346 ;
  assign n2739 = ~n698 & ~n2738 ;
  assign n2740 = n866 & ~n2739 ;
  assign n2741 = x11 & n404 ;
  assign n2742 = n104 & n869 ;
  assign n2743 = ~n2741 & ~n2742 ;
  assign n2744 = ~x0 & ~n2743 ;
  assign n2745 = ~n2740 & ~n2744 ;
  assign n2746 = n1407 & ~n2745 ;
  assign n2747 = ~x0 & ~x9 ;
  assign n2748 = n418 & n1656 ;
  assign n2749 = n2747 & n2748 ;
  assign n2750 = ~x11 & n2749 ;
  assign n2751 = ~n2746 & ~n2750 ;
  assign n2752 = ~n2737 & n2751 ;
  assign n2753 = n843 & ~n2752 ;
  assign n2754 = ~x8 & n2036 ;
  assign n2755 = ~x6 & x9 ;
  assign n2756 = n489 & n2755 ;
  assign n2757 = n2754 & n2756 ;
  assign n2758 = n2280 & n2757 ;
  assign n2759 = ~n2753 & ~n2758 ;
  assign n2760 = ~x7 & ~n2759 ;
  assign n2761 = n240 & n265 ;
  assign n2762 = n2761 ^ n2708 ;
  assign n2763 = n1658 ^ x0 ;
  assign n2764 = n2763 ^ n1658 ;
  assign n2765 = n1658 ^ n1423 ;
  assign n2766 = ~n2764 & ~n2765 ;
  assign n2767 = n2766 ^ n1658 ;
  assign n2768 = n2767 ^ n2761 ;
  assign n2769 = n2762 & ~n2768 ;
  assign n2770 = n2769 ^ n2766 ;
  assign n2771 = n2770 ^ n1658 ;
  assign n2772 = n2771 ^ n2708 ;
  assign n2773 = n2761 & ~n2772 ;
  assign n2774 = n2773 ^ n2761 ;
  assign n2775 = ~n2760 & ~n2774 ;
  assign n2776 = n1936 & ~n2775 ;
  assign n2777 = ~n354 & n2512 ;
  assign n2778 = ~x6 & n571 ;
  assign n2779 = n555 & n2778 ;
  assign n2780 = n2777 & n2779 ;
  assign n2781 = n34 & n2686 ;
  assign n2782 = n1423 & n2781 ;
  assign n2783 = ~x9 & n1656 ;
  assign n2784 = n89 & n2783 ;
  assign n2785 = ~x6 & n1263 ;
  assign n2786 = x0 & n2785 ;
  assign n2787 = ~n1715 & ~n2786 ;
  assign n2788 = n411 & ~n2787 ;
  assign n2789 = ~n2784 & ~n2788 ;
  assign n2790 = ~n2782 & n2789 ;
  assign n2791 = n1050 & ~n2790 ;
  assign n2792 = ~n2780 & ~n2791 ;
  assign n2793 = n225 & n418 ;
  assign n2794 = ~n2792 & n2793 ;
  assign n2795 = n262 & n2794 ;
  assign n2838 = x4 & n492 ;
  assign n2839 = x6 & ~x10 ;
  assign n2822 = ~x7 & n34 ;
  assign n2840 = n1328 & n2822 ;
  assign n2841 = ~x13 & n2653 ;
  assign n2842 = n1246 & n2841 ;
  assign n2810 = ~x12 & n762 ;
  assign n2843 = ~n497 & n2810 ;
  assign n2844 = ~n2559 & n2843 ;
  assign n2845 = ~n2842 & ~n2844 ;
  assign n2846 = ~n2840 & n2845 ;
  assign n2847 = n2839 & ~n2846 ;
  assign n2848 = x5 & ~x7 ;
  assign n2849 = ~x0 & n2848 ;
  assign n2850 = x6 & x13 ;
  assign n2851 = n1657 & n2850 ;
  assign n2852 = n2849 & n2851 ;
  assign n2853 = ~x6 & n89 ;
  assign n2854 = n471 & n2512 ;
  assign n2855 = n2853 & n2854 ;
  assign n2856 = ~n2852 & ~n2855 ;
  assign n2857 = ~n2847 & n2856 ;
  assign n2858 = n2838 & ~n2857 ;
  assign n2859 = n1201 & n2631 ;
  assign n2860 = n2704 & n2859 ;
  assign n2861 = n471 & n843 ;
  assign n2862 = ~n2691 & ~n2861 ;
  assign n2863 = x9 & n884 ;
  assign n2864 = n2182 & n2863 ;
  assign n2865 = ~n2862 & n2864 ;
  assign n2866 = ~n2860 & ~n2865 ;
  assign n2867 = ~x3 & ~n2866 ;
  assign n2868 = ~x0 & n405 ;
  assign n2869 = n1327 & n2868 ;
  assign n2870 = ~x5 & n2608 ;
  assign n2871 = n1025 & n2870 ;
  assign n2872 = n2869 & n2871 ;
  assign n2873 = ~x5 & ~x12 ;
  assign n2874 = n888 & n2608 ;
  assign n2875 = n2873 & n2874 ;
  assign n2876 = n827 & n2036 ;
  assign n2877 = ~x4 & n2707 ;
  assign n2878 = n2876 & n2877 ;
  assign n2879 = ~n2875 & ~n2878 ;
  assign n2880 = n284 & ~n2879 ;
  assign n2881 = x6 & ~x7 ;
  assign n2882 = n795 & n2881 ;
  assign n2883 = n404 & n2882 ;
  assign n2884 = n1671 & n2883 ;
  assign n2885 = ~n2880 & ~n2884 ;
  assign n2886 = n762 & ~n2885 ;
  assign n2887 = ~n2872 & ~n2886 ;
  assign n2888 = ~n2867 & n2887 ;
  assign n2889 = ~n2858 & n2888 ;
  assign n2796 = ~x12 & n874 ;
  assign n2797 = n1618 & n2480 ;
  assign n2798 = n2796 & n2797 ;
  assign n2799 = ~x4 & n1423 ;
  assign n2800 = n1002 & n2799 ;
  assign n2801 = n404 & n2800 ;
  assign n2802 = ~n2798 & ~n2801 ;
  assign n2803 = ~x3 & ~x11 ;
  assign n2804 = n2707 & n2803 ;
  assign n2805 = ~n2802 & n2804 ;
  assign n2806 = x6 & x7 ;
  assign n2807 = ~x9 & n2806 ;
  assign n2808 = n2118 & n2807 ;
  assign n2809 = n1683 & n2808 ;
  assign n2811 = ~x6 & ~x13 ;
  assign n2812 = n1025 & n2811 ;
  assign n2813 = n2810 & n2812 ;
  assign n2814 = n517 & n2036 ;
  assign n2815 = ~x0 & ~x6 ;
  assign n2816 = ~x7 & n2815 ;
  assign n2817 = n2814 & n2816 ;
  assign n2818 = ~n2813 & ~n2817 ;
  assign n2819 = ~n2809 & n2818 ;
  assign n2820 = ~x3 & n739 ;
  assign n2821 = ~n2819 & n2820 ;
  assign n2823 = ~x10 & n2608 ;
  assign n2824 = ~x9 & n1327 ;
  assign n2825 = n2823 & n2824 ;
  assign n2826 = ~x4 & n2755 ;
  assign n2827 = ~x13 & n1423 ;
  assign n2828 = n2826 & n2827 ;
  assign n2829 = ~n2825 & ~n2828 ;
  assign n2830 = n659 & ~n2829 ;
  assign n2831 = x6 & n366 ;
  assign n2832 = n2720 & n2831 ;
  assign n2833 = ~x12 & n2832 ;
  assign n2834 = ~n2830 & ~n2833 ;
  assign n2835 = n2822 & ~n2834 ;
  assign n2836 = ~n2821 & ~n2835 ;
  assign n2837 = ~n2805 & n2836 ;
  assign n2890 = n2889 ^ n2837 ;
  assign n2891 = n2889 ^ x14 ;
  assign n2892 = n2891 ^ n2889 ;
  assign n2893 = n2892 ^ n112 ;
  assign n2894 = n2893 ^ x8 ;
  assign n2895 = n2890 & ~n2894 ;
  assign n2896 = n2895 ^ n2889 ;
  assign n2897 = n112 & n2896 ;
  assign n2898 = n2897 ^ n112 ;
  assign n2899 = ~n2795 & ~n2898 ;
  assign n2900 = ~n2776 & n2899 ;
  assign n2901 = ~x5 & x7 ;
  assign n2902 = ~n2848 & ~n2901 ;
  assign n2903 = n106 & n2562 ;
  assign n2904 = n1010 & n1514 ;
  assign n2905 = ~x10 & n1363 ;
  assign n2906 = ~n110 & n2905 ;
  assign n2907 = ~n2904 & ~n2906 ;
  assign n2908 = n2903 & ~n2907 ;
  assign n2909 = ~n525 & ~n1104 ;
  assign n2910 = x6 & ~x8 ;
  assign n2911 = n1495 & n2910 ;
  assign n2912 = ~n2909 & n2911 ;
  assign n2913 = x11 & n58 ;
  assign n2914 = ~n2613 & ~n2874 ;
  assign n2915 = n2913 & ~n2914 ;
  assign n2916 = n471 & n2608 ;
  assign n2917 = ~x6 & n1880 ;
  assign n2918 = n889 & n2917 ;
  assign n2919 = ~n2916 & ~n2918 ;
  assign n2920 = ~n741 & ~n2919 ;
  assign n2921 = ~n2915 & ~n2920 ;
  assign n2922 = n162 & ~n2921 ;
  assign n2923 = ~n2912 & ~n2922 ;
  assign n2924 = ~n2908 & n2923 ;
  assign n2927 = n2924 ^ x13 ;
  assign n2928 = n2927 ^ n2924 ;
  assign n2925 = n2924 ^ n2917 ;
  assign n2926 = n2925 ^ n2924 ;
  assign n2929 = n2928 ^ n2926 ;
  assign n2930 = n262 & ~n1136 ;
  assign n2931 = n1108 & n1514 ;
  assign n2932 = ~n1203 & ~n2931 ;
  assign n2933 = ~n2930 & n2932 ;
  assign n2934 = n2933 ^ n2924 ;
  assign n2935 = n2934 ^ n2924 ;
  assign n2936 = n2935 ^ n2928 ;
  assign n2937 = ~n2928 & n2936 ;
  assign n2938 = n2937 ^ n2928 ;
  assign n2939 = ~n2929 & ~n2938 ;
  assign n2940 = n2939 ^ n2937 ;
  assign n2941 = n2940 ^ n2924 ;
  assign n2942 = n2941 ^ n2928 ;
  assign n2943 = x14 & n2942 ;
  assign n2944 = n2943 ^ n2924 ;
  assign n2945 = n1263 & ~n2944 ;
  assign n2952 = n248 & n1678 ;
  assign n2953 = n727 & n845 ;
  assign n2954 = ~n2952 & ~n2953 ;
  assign n2955 = ~x6 & n106 ;
  assign n2956 = ~n2954 & n2955 ;
  assign n2957 = n471 & n1327 ;
  assign n2958 = n2903 & n2957 ;
  assign n2959 = n1407 & n2608 ;
  assign n2960 = n381 & ~n869 ;
  assign n2961 = n2959 & n2960 ;
  assign n2962 = ~n2958 & ~n2961 ;
  assign n2963 = ~n2956 & n2962 ;
  assign n2946 = n642 & n1671 ;
  assign n2947 = n2608 & n2946 ;
  assign n2948 = ~x13 & n1246 ;
  assign n2949 = ~n474 & ~n2948 ;
  assign n2950 = n2535 & ~n2949 ;
  assign n2951 = ~n2947 & ~n2950 ;
  assign n2964 = n2963 ^ n2951 ;
  assign n2965 = n2964 ^ n2963 ;
  assign n2966 = n2963 ^ n798 ;
  assign n2967 = n2966 ^ n2963 ;
  assign n2968 = ~n2965 & n2967 ;
  assign n2969 = n2968 ^ n2963 ;
  assign n2970 = ~x2 & ~n2969 ;
  assign n2971 = n2970 ^ n2963 ;
  assign n2972 = n1559 & ~n2971 ;
  assign n2973 = ~x6 & n195 ;
  assign n2974 = n946 & n2973 ;
  assign n2975 = n2224 & n2608 ;
  assign n2976 = ~n2613 & ~n2975 ;
  assign n2977 = ~n741 & ~n2976 ;
  assign n2978 = ~n2974 & ~n2977 ;
  assign n2979 = n2978 ^ x13 ;
  assign n2980 = n2979 ^ n2978 ;
  assign n2981 = n2980 ^ n1151 ;
  assign n2982 = n2975 ^ n58 ;
  assign n2983 = n2975 & n2982 ;
  assign n2984 = n2983 ^ n2978 ;
  assign n2985 = n2984 ^ n2975 ;
  assign n2986 = ~n2981 & ~n2985 ;
  assign n2987 = n2986 ^ n2983 ;
  assign n2988 = n2987 ^ n2975 ;
  assign n2989 = ~n1151 & n2988 ;
  assign n2990 = n328 & n2989 ;
  assign n2991 = ~x3 & ~x14 ;
  assign n2992 = n1876 & n2991 ;
  assign n2993 = n2850 & n2992 ;
  assign n2994 = n777 & n2993 ;
  assign n2995 = n58 & n2535 ;
  assign n2996 = ~x14 & n473 ;
  assign n2997 = n230 & n2996 ;
  assign n2998 = n2995 & n2997 ;
  assign n2999 = ~n2994 & ~n2998 ;
  assign n3000 = ~n2990 & n2999 ;
  assign n3001 = n1364 & ~n3000 ;
  assign n3002 = ~x3 & n2535 ;
  assign n3003 = ~x12 & n673 ;
  assign n3004 = n2913 & n3003 ;
  assign n3005 = n3002 & n3004 ;
  assign n3006 = n463 & n3005 ;
  assign n3007 = ~n3001 & ~n3006 ;
  assign n3008 = ~n2972 & n3007 ;
  assign n3009 = ~x12 & n596 ;
  assign n3010 = x2 & ~x14 ;
  assign n3011 = n471 & n3010 ;
  assign n3012 = ~n1905 & ~n2560 ;
  assign n3013 = ~n20 & ~n784 ;
  assign n3014 = ~n978 & ~n3013 ;
  assign n3015 = ~n3012 & n3014 ;
  assign n3016 = ~n3011 & ~n3015 ;
  assign n3017 = n3009 & ~n3016 ;
  assign n3018 = n2608 & n3017 ;
  assign n3019 = x2 & x14 ;
  assign n3020 = ~n1658 & n3019 ;
  assign n3021 = x12 & ~x14 ;
  assign n3022 = n784 & n3021 ;
  assign n3023 = ~n3020 & ~n3022 ;
  assign n3024 = n240 & ~n3023 ;
  assign n3025 = n2535 & n3024 ;
  assign n3026 = ~x2 & n3021 ;
  assign n3027 = n2916 & n3026 ;
  assign n3028 = ~n3025 & ~n3027 ;
  assign n3029 = n798 & ~n3028 ;
  assign n3030 = x12 & x14 ;
  assign n3031 = n2535 & n3030 ;
  assign n3032 = n740 & n1010 ;
  assign n3033 = n418 & n3032 ;
  assign n3034 = n3031 & n3033 ;
  assign n3035 = ~n3029 & ~n3034 ;
  assign n3036 = ~n3018 & n3035 ;
  assign n3037 = n2290 & n2560 ;
  assign n3038 = n964 & n3037 ;
  assign n3039 = n76 & n845 ;
  assign n3040 = ~n2996 & ~n3039 ;
  assign n3041 = n364 & ~n3040 ;
  assign n3042 = n890 ^ x10 ;
  assign n3043 = n890 ^ x11 ;
  assign n3044 = n3043 ^ n890 ;
  assign n3045 = n3042 & n3044 ;
  assign n3046 = n3045 ^ n890 ;
  assign n3047 = n3026 & n3046 ;
  assign n3048 = ~n3041 & ~n3047 ;
  assign n3049 = ~n3038 & n3048 ;
  assign n3050 = n3049 ^ n3024 ;
  assign n3051 = n3024 ^ x0 ;
  assign n3052 = n3051 ^ n3024 ;
  assign n3053 = n3052 ^ n2955 ;
  assign n3054 = n3053 ^ n106 ;
  assign n3055 = ~n3050 & n3054 ;
  assign n3056 = n3055 ^ n3024 ;
  assign n3057 = n2955 & ~n3056 ;
  assign n3058 = n3057 ^ n2955 ;
  assign n3059 = n3036 & ~n3058 ;
  assign n3060 = n284 & ~n3059 ;
  assign n3061 = n3008 & ~n3060 ;
  assign n3062 = ~n2945 & n3061 ;
  assign n3063 = ~n2902 & ~n3062 ;
  assign n3064 = n2900 & ~n3063 ;
  assign n3065 = ~n2734 & n3064 ;
  assign n3123 = n26 & n2562 ;
  assign n3124 = n859 & n3123 ;
  assign n3125 = ~x5 & n105 ;
  assign n3126 = n2686 & n3125 ;
  assign n3127 = n1476 & n3126 ;
  assign n3128 = x6 ^ x4 ;
  assign n3129 = n3128 ^ n818 ;
  assign n3130 = ~n39 & ~n1991 ;
  assign n3131 = n3130 ^ n2559 ;
  assign n3132 = n2559 ^ x4 ;
  assign n3133 = n3132 ^ n2559 ;
  assign n3134 = n3131 & ~n3133 ;
  assign n3135 = n3134 ^ n2559 ;
  assign n3136 = n3135 ^ n3128 ;
  assign n3137 = n3129 & ~n3136 ;
  assign n3138 = n3137 ^ n3134 ;
  assign n3139 = n3138 ^ n2559 ;
  assign n3140 = n3139 ^ n818 ;
  assign n3141 = n3128 & ~n3140 ;
  assign n3142 = n3141 ^ n3128 ;
  assign n3143 = ~n3127 & ~n3142 ;
  assign n3144 = ~n3124 & n3143 ;
  assign n3145 = n1665 & ~n3144 ;
  assign n3146 = ~x9 & n1226 ;
  assign n3147 = n26 & n2684 ;
  assign n3148 = n224 & n3147 ;
  assign n3149 = n3146 & n3148 ;
  assign n3150 = n17 & n346 ;
  assign n3151 = n650 & n3150 ;
  assign n3152 = n3123 & n3151 ;
  assign n3153 = ~n3149 & ~n3152 ;
  assign n3154 = ~n3145 & n3153 ;
  assign n3066 = n818 & n3003 ;
  assign n3067 = n1464 & n2608 ;
  assign n3068 = n3066 & n3067 ;
  assign n3069 = n3068 ^ x3 ;
  assign n3070 = n243 & n2356 ;
  assign n3071 = n858 & n3070 ;
  assign n3072 = ~x14 & n2608 ;
  assign n3073 = n1025 & n1246 ;
  assign n3074 = n3072 & n3073 ;
  assign n3075 = ~x4 & ~x9 ;
  assign n3076 = n334 & n3075 ;
  assign n3077 = n17 & n3076 ;
  assign n3078 = ~n3074 & ~n3077 ;
  assign n3079 = ~x5 & ~n3078 ;
  assign n3080 = ~n2537 & ~n2668 ;
  assign n3081 = n76 & n346 ;
  assign n3082 = n2848 & n3081 ;
  assign n3083 = ~n3080 & n3082 ;
  assign n3084 = ~n3079 & ~n3083 ;
  assign n3085 = ~n3071 & n3084 ;
  assign n3086 = n3085 ^ x0 ;
  assign n3087 = n3086 ^ n3085 ;
  assign n3088 = n76 & n1422 ;
  assign n3089 = n346 & n3088 ;
  assign n3090 = n1641 & n3089 ;
  assign n3091 = ~x7 & x14 ;
  assign n3092 = ~x5 & n3091 ;
  assign n3093 = n2535 & n3092 ;
  assign n3094 = ~x12 & n2608 ;
  assign n3095 = n2583 & n3094 ;
  assign n3096 = ~n3093 & ~n3095 ;
  assign n3097 = n346 & ~n3096 ;
  assign n3098 = x6 & ~x14 ;
  assign n3099 = n517 & n2512 ;
  assign n3100 = n1538 & n3099 ;
  assign n3101 = n3098 & n3100 ;
  assign n3102 = ~n3097 & ~n3101 ;
  assign n3103 = x13 & ~n3102 ;
  assign n3104 = ~x4 & x7 ;
  assign n3105 = ~n1630 & ~n1641 ;
  assign n3106 = x5 & x6 ;
  assign n3107 = n3081 & ~n3106 ;
  assign n3108 = n3105 & n3107 ;
  assign n3109 = n3104 & n3108 ;
  assign n3110 = ~n3103 & ~n3109 ;
  assign n3111 = ~n3090 & n3110 ;
  assign n3112 = n3111 ^ n3085 ;
  assign n3113 = n3087 & n3112 ;
  assign n3114 = n3113 ^ n3085 ;
  assign n3115 = n3114 ^ n3068 ;
  assign n3116 = ~n3069 & n3115 ;
  assign n3117 = n3116 ^ n3113 ;
  assign n3118 = n3117 ^ n3085 ;
  assign n3119 = n3118 ^ x3 ;
  assign n3120 = ~n3068 & ~n3119 ;
  assign n3121 = n3120 ^ n3068 ;
  assign n3122 = n3121 ^ n3068 ;
  assign n3155 = n3154 ^ n3122 ;
  assign n3156 = n3155 ^ n3122 ;
  assign n3157 = n3122 ^ x14 ;
  assign n3158 = n3157 ^ n3122 ;
  assign n3159 = ~n3156 & ~n3158 ;
  assign n3160 = n3159 ^ n3122 ;
  assign n3161 = x2 & ~n3160 ;
  assign n3162 = n3161 ^ n3122 ;
  assign n3163 = ~n467 & ~n3162 ;
  assign n3164 = n20 & n2991 ;
  assign n3165 = x7 & x8 ;
  assign n3166 = n1328 & n3165 ;
  assign n3167 = n2576 & n3166 ;
  assign n3168 = ~n105 & n263 ;
  assign n3169 = ~n2761 & ~n3168 ;
  assign n3170 = n17 & n2613 ;
  assign n3171 = ~n3169 & n3170 ;
  assign n3172 = n392 & n1657 ;
  assign n3173 = n263 & n3172 ;
  assign n3174 = n2701 & n3173 ;
  assign n3175 = ~x7 & n1327 ;
  assign n3176 = ~n2570 & n3175 ;
  assign n3177 = n471 & n2036 ;
  assign n3178 = n2638 & n3177 ;
  assign n3179 = ~n3176 & ~n3178 ;
  assign n3180 = n2608 & ~n3179 ;
  assign n3181 = ~n3174 & ~n3180 ;
  assign n3182 = ~n3171 & n3181 ;
  assign n3183 = x5 & ~n3182 ;
  assign n3184 = ~n3167 & ~n3183 ;
  assign n3185 = n3164 & ~n3184 ;
  assign n3225 = ~x14 & n828 ;
  assign n3226 = n224 & n3225 ;
  assign n3227 = ~x0 & ~n328 ;
  assign n3228 = ~x14 & n1665 ;
  assign n3229 = ~n1282 & ~n3021 ;
  assign n3230 = x3 & ~n3229 ;
  assign n3231 = x0 & ~n3230 ;
  assign n3232 = ~n3228 & n3231 ;
  assign n3233 = x13 & ~n3232 ;
  assign n3234 = ~n3227 & n3233 ;
  assign n3235 = ~n3226 & ~n3234 ;
  assign n3186 = ~x6 & x8 ;
  assign n3187 = ~x4 & n3186 ;
  assign n3188 = n1423 & n3187 ;
  assign n3189 = n673 & n2653 ;
  assign n3190 = n3188 & n3189 ;
  assign n3191 = n673 & n2806 ;
  assign n3192 = n76 & n2848 ;
  assign n3193 = ~x6 & n3192 ;
  assign n3194 = ~n3191 & ~n3193 ;
  assign n3195 = n1948 & ~n3194 ;
  assign n3196 = ~x5 & ~x7 ;
  assign n3197 = n718 & n3196 ;
  assign n3198 = n2535 & n3197 ;
  assign n3199 = n363 & n828 ;
  assign n3200 = n844 & n3199 ;
  assign n3201 = ~n3198 & ~n3200 ;
  assign n3202 = ~n3195 & n3201 ;
  assign n3203 = n2224 & ~n3202 ;
  assign n3204 = ~n3190 & ~n3203 ;
  assign n3205 = n68 & ~n3204 ;
  assign n3206 = ~x5 & ~x10 ;
  assign n3207 = n2608 & n3206 ;
  assign n3208 = n76 & n1407 ;
  assign n3209 = x3 & n2458 ;
  assign n3210 = n3208 & n3209 ;
  assign n3211 = n3207 & n3210 ;
  assign n3212 = ~x14 & n1423 ;
  assign n3213 = n151 & n2709 ;
  assign n3214 = n2653 & n3002 ;
  assign n3215 = n175 & n3214 ;
  assign n3216 = ~n3213 & ~n3215 ;
  assign n3217 = n3212 & ~n3216 ;
  assign n3218 = n799 & n3003 ;
  assign n3219 = n2882 & n3218 ;
  assign n3220 = ~n3217 & ~n3219 ;
  assign n3221 = ~n3211 & n3220 ;
  assign n3222 = ~n3205 & n3221 ;
  assign n3236 = n3235 ^ n3222 ;
  assign n3237 = n3236 ^ n3222 ;
  assign n3223 = n3222 ^ n2721 ;
  assign n3224 = n3223 ^ n3222 ;
  assign n3238 = n3237 ^ n3224 ;
  assign n3239 = n3222 ^ n2224 ;
  assign n3240 = n3239 ^ n3222 ;
  assign n3241 = n3240 ^ n3237 ;
  assign n3242 = ~n3237 & ~n3241 ;
  assign n3243 = n3242 ^ n3237 ;
  assign n3244 = ~n3238 & ~n3243 ;
  assign n3245 = n3244 ^ n3242 ;
  assign n3246 = n3245 ^ n3222 ;
  assign n3247 = n3246 ^ n3237 ;
  assign n3248 = ~x2 & n3247 ;
  assign n3249 = n3248 ^ n3222 ;
  assign n3250 = ~n555 & ~n3249 ;
  assign n3251 = ~n3185 & ~n3250 ;
  assign n3252 = ~n3163 & n3251 ;
  assign n3253 = n3065 & n3252 ;
  assign n3254 = ~n2652 & n3253 ;
  assign n3255 = ~x1 & ~n3254 ;
  assign n3256 = x8 & ~x14 ;
  assign n3257 = ~x0 & n757 ;
  assign n3258 = ~x7 & n2608 ;
  assign n3259 = n3125 & n3258 ;
  assign n3260 = n3257 & n3259 ;
  assign n3261 = ~x0 & n213 ;
  assign n3262 = n859 & n3261 ;
  assign n3263 = x2 & ~x7 ;
  assign n3264 = ~x0 & n3263 ;
  assign n3265 = n2738 & n3264 ;
  assign n3266 = ~n1524 & n2863 ;
  assign n3267 = n869 & n3266 ;
  assign n3268 = ~n3265 & ~n3267 ;
  assign n3269 = x5 & ~n3268 ;
  assign n3270 = ~n3262 & ~n3269 ;
  assign n3271 = n2535 & ~n3270 ;
  assign n3272 = ~n3260 & ~n3271 ;
  assign n3273 = n3256 & ~n3272 ;
  assign n3274 = n1807 & n3191 ;
  assign n3275 = n2064 & n3274 ;
  assign n3276 = ~n3273 & ~n3275 ;
  assign n3277 = ~n1658 & ~n3276 ;
  assign n3278 = n784 & n3125 ;
  assign n3279 = x5 & n946 ;
  assign n3280 = ~n869 & n3279 ;
  assign n3281 = ~n572 & ~n3280 ;
  assign n3282 = ~n3278 & n3281 ;
  assign n3283 = ~x10 & n105 ;
  assign n3284 = n180 & n3283 ;
  assign n3285 = x0 & ~n3284 ;
  assign n3286 = ~x7 & ~x12 ;
  assign n3287 = x6 & x8 ;
  assign n3288 = x4 & ~x14 ;
  assign n3289 = n3287 & n3288 ;
  assign n3290 = n3286 & n3289 ;
  assign n3291 = ~n3285 & n3290 ;
  assign n3292 = ~n3282 & n3291 ;
  assign n3293 = ~x0 & ~n1658 ;
  assign n3294 = ~x5 & n1025 ;
  assign n3295 = ~x6 & n42 ;
  assign n3296 = n3294 & n3295 ;
  assign n3297 = ~n1538 & ~n2881 ;
  assign n3298 = ~n720 & ~n997 ;
  assign n3299 = ~n3297 & ~n3298 ;
  assign n3300 = n885 & n3299 ;
  assign n3301 = ~n3296 & ~n3300 ;
  assign n3302 = n334 & ~n3301 ;
  assign n3303 = n3293 & n3302 ;
  assign n3304 = ~n3292 & ~n3303 ;
  assign n3305 = ~n175 & ~n798 ;
  assign n3306 = x13 & n2653 ;
  assign n3307 = x11 & ~x14 ;
  assign n3308 = n3306 & n3307 ;
  assign n3309 = ~n3305 & n3308 ;
  assign n3310 = x11 ^ x5 ;
  assign n3311 = n44 ^ x11 ;
  assign n3312 = n3311 ^ n44 ;
  assign n3313 = n3010 ^ n44 ;
  assign n3314 = n3312 & n3313 ;
  assign n3315 = n3314 ^ n44 ;
  assign n3316 = ~n3310 & n3315 ;
  assign n3317 = n798 & n3316 ;
  assign n3318 = ~x14 & n740 ;
  assign n3319 = ~x5 & n406 ;
  assign n3320 = n3318 & n3319 ;
  assign n3321 = n86 & n1524 ;
  assign n3322 = ~n3320 & ~n3321 ;
  assign n3323 = ~n3317 & n3322 ;
  assign n3324 = n2678 & ~n3323 ;
  assign n3325 = ~n3309 & ~n3324 ;
  assign n3326 = ~n2587 & ~n2693 ;
  assign n3327 = ~n2669 & ~n3094 ;
  assign n3328 = n3326 & ~n3327 ;
  assign n3329 = ~n3325 & n3328 ;
  assign n3330 = x2 & n866 ;
  assign n3331 = x8 ^ x5 ;
  assign n3332 = n3331 ^ x13 ;
  assign n3342 = n3332 ^ x5 ;
  assign n3339 = n2467 ^ n1151 ;
  assign n3343 = n3339 ^ n2653 ;
  assign n3344 = n3343 ^ x5 ;
  assign n3345 = ~n3342 & n3344 ;
  assign n3333 = x13 ^ x5 ;
  assign n3334 = n3333 ^ n3332 ;
  assign n3335 = n3334 ^ n1151 ;
  assign n3336 = n3335 ^ n1151 ;
  assign n3337 = n3336 ^ n3332 ;
  assign n3338 = n3337 ^ x5 ;
  assign n3340 = n3339 ^ n1151 ;
  assign n3341 = n3338 & n3340 ;
  assign n3346 = n3345 ^ n3341 ;
  assign n3347 = n3346 ^ n3339 ;
  assign n3348 = n3347 ^ n2653 ;
  assign n3349 = n3348 ^ n3338 ;
  assign n3350 = n3341 ^ n1151 ;
  assign n3351 = n3345 ^ n3339 ;
  assign n3352 = n3351 ^ n2653 ;
  assign n3353 = n3352 ^ n1151 ;
  assign n3354 = n3353 ^ n3342 ;
  assign n3355 = n3350 & n3354 ;
  assign n3356 = n3355 ^ n3341 ;
  assign n3357 = ~n3349 & n3356 ;
  assign n3358 = n3094 & n3357 ;
  assign n3359 = n3330 & n3358 ;
  assign n3360 = ~x6 & ~n2559 ;
  assign n3361 = ~x5 & n2806 ;
  assign n3362 = x13 & n3361 ;
  assign n3363 = ~n3360 & ~n3362 ;
  assign n3364 = n1948 & ~n3363 ;
  assign n3365 = ~x13 & n2537 ;
  assign n3366 = ~x7 & n2668 ;
  assign n3367 = ~n3365 & ~n3366 ;
  assign n3368 = n26 & ~n3367 ;
  assign n3369 = ~n17 & ~n1327 ;
  assign n3370 = n739 & ~n3080 ;
  assign n3371 = ~n3369 & n3370 ;
  assign n3372 = ~n3368 & ~n3371 ;
  assign n3373 = ~n3364 & n3372 ;
  assign n3374 = n463 & ~n3373 ;
  assign n3375 = ~n39 & n2902 ;
  assign n3376 = n2975 & ~n3375 ;
  assign n3377 = x12 & n3376 ;
  assign n3378 = x8 & n2875 ;
  assign n3379 = ~n3377 & ~n3378 ;
  assign n3380 = ~n3374 & n3379 ;
  assign n3381 = n226 & ~n3380 ;
  assign n3382 = ~n40 & n843 ;
  assign n3383 = n2512 ^ x13 ;
  assign n3384 = n3383 ^ x2 ;
  assign n3391 = n3384 ^ n3383 ;
  assign n3385 = n3384 ^ n17 ;
  assign n3386 = n3385 ^ n3383 ;
  assign n3387 = n3384 ^ n2512 ;
  assign n3388 = n3387 ^ n17 ;
  assign n3389 = n3388 ^ n3386 ;
  assign n3390 = n3386 & n3389 ;
  assign n3392 = n3391 ^ n3390 ;
  assign n3393 = n3392 ^ n3386 ;
  assign n3394 = n3383 ^ n1948 ;
  assign n3395 = n3390 ^ n3386 ;
  assign n3396 = n3394 & n3395 ;
  assign n3397 = n3396 ^ n3383 ;
  assign n3398 = ~n3393 & ~n3397 ;
  assign n3399 = n3398 ^ n3383 ;
  assign n3400 = n3399 ^ x13 ;
  assign n3401 = n3400 ^ n3383 ;
  assign n3402 = n3382 & ~n3401 ;
  assign n3403 = x5 & n2575 ;
  assign n3404 = n2678 & n3403 ;
  assign n3405 = n1146 & n3404 ;
  assign n3406 = ~n3402 & ~n3405 ;
  assign n3407 = n796 & ~n3406 ;
  assign n3408 = x12 & n2653 ;
  assign n3409 = n418 & n3408 ;
  assign n3410 = n180 & n3009 ;
  assign n3411 = ~n3409 & ~n3410 ;
  assign n3412 = n242 & n2587 ;
  assign n3413 = ~n3411 & n3412 ;
  assign n3414 = n712 & n2910 ;
  assign n3415 = n2023 & n3414 ;
  assign n3416 = n2569 & n3415 ;
  assign n3417 = ~n3413 & ~n3416 ;
  assign n3418 = x12 & n524 ;
  assign n3419 = n430 & n2870 ;
  assign n3420 = x8 & n26 ;
  assign n3421 = n2811 & n3420 ;
  assign n3422 = ~n3419 & ~n3421 ;
  assign n3423 = n3263 & ~n3422 ;
  assign n3424 = ~x8 & n2678 ;
  assign n3425 = x6 & n795 ;
  assign n3426 = n3424 & n3425 ;
  assign n3427 = x2 & ~x6 ;
  assign n3428 = n106 & n3427 ;
  assign n3429 = n2558 & n3428 ;
  assign n3430 = ~x5 & n3429 ;
  assign n3431 = ~n3426 & ~n3430 ;
  assign n3432 = ~n3423 & n3431 ;
  assign n3433 = n3418 & ~n3432 ;
  assign n3434 = n3417 & ~n3433 ;
  assign n3435 = ~n3407 & n3434 ;
  assign n3436 = ~n3381 & n3435 ;
  assign n3437 = n3436 ^ x0 ;
  assign n3438 = n3437 ^ n3436 ;
  assign n3439 = n3438 ^ n3359 ;
  assign n3440 = n2557 & n3094 ;
  assign n3441 = n862 & n2669 ;
  assign n3442 = ~x13 & n3441 ;
  assign n3443 = ~n3440 & ~n3442 ;
  assign n3444 = n292 & ~n3443 ;
  assign n3445 = ~n226 & n3444 ;
  assign n3446 = n151 & n3147 ;
  assign n3447 = n1226 & n3446 ;
  assign n3448 = ~n3445 & ~n3447 ;
  assign n3449 = n3448 ^ x10 ;
  assign n3450 = ~n3448 & ~n3449 ;
  assign n3451 = n3450 ^ n3436 ;
  assign n3452 = n3451 ^ n3448 ;
  assign n3453 = ~n3439 & n3452 ;
  assign n3454 = n3453 ^ n3450 ;
  assign n3455 = n3454 ^ n3448 ;
  assign n3456 = ~n3359 & ~n3455 ;
  assign n3457 = n3456 ^ n3359 ;
  assign n3458 = n3457 ^ x14 ;
  assign n3459 = n3458 ^ n3457 ;
  assign n3460 = n3459 ^ n3329 ;
  assign n3461 = n1671 & n3259 ;
  assign n3462 = n889 & n1226 ;
  assign n3463 = n3147 & n3462 ;
  assign n3464 = ~n3461 & ~n3463 ;
  assign n3465 = ~n3305 & ~n3464 ;
  assign n3466 = ~x7 & n2875 ;
  assign n3467 = ~x4 & ~n2902 ;
  assign n3468 = n2827 & n3467 ;
  assign n3469 = ~x6 & n3468 ;
  assign n3470 = ~n3466 & ~n3469 ;
  assign n3471 = n406 & ~n3470 ;
  assign n3472 = ~x0 & n3471 ;
  assign n3473 = ~n3465 & ~n3472 ;
  assign n3474 = n3473 ^ x2 ;
  assign n3475 = x2 & ~n3474 ;
  assign n3476 = n3475 ^ n3457 ;
  assign n3477 = n3476 ^ x2 ;
  assign n3478 = ~n3460 & n3477 ;
  assign n3479 = n3478 ^ n3475 ;
  assign n3480 = n3479 ^ x2 ;
  assign n3481 = ~n3329 & n3480 ;
  assign n3482 = n3481 ^ n3329 ;
  assign n3483 = n3482 ^ x9 ;
  assign n3484 = n3483 ^ n3482 ;
  assign n3485 = ~n948 & ~n1217 ;
  assign n3486 = ~n1136 & n3485 ;
  assign n3487 = n213 & n2509 ;
  assign n3488 = n3486 & n3487 ;
  assign n3489 = n1165 & ~n2902 ;
  assign n3490 = ~x5 & x10 ;
  assign n3491 = n920 & n3490 ;
  assign n3492 = ~n3489 & ~n3491 ;
  assign n3493 = n3287 & ~n3492 ;
  assign n3494 = ~n2910 & ~n3186 ;
  assign n3495 = n866 & ~n3494 ;
  assign n3496 = x6 & n1078 ;
  assign n3497 = ~n3495 & ~n3496 ;
  assign n3498 = n1435 & ~n3497 ;
  assign n3499 = ~n2690 & ~n2861 ;
  assign n3500 = n175 & ~n3499 ;
  assign n3501 = ~n3498 & ~n3500 ;
  assign n3502 = n3263 & ~n3501 ;
  assign n3503 = ~n3493 & ~n3502 ;
  assign n3504 = ~n3488 & n3503 ;
  assign n3505 = n2646 & ~n3504 ;
  assign n3506 = x6 & n786 ;
  assign n3507 = n3283 & n3506 ;
  assign n3508 = n740 & ~n2902 ;
  assign n3509 = n3507 & n3508 ;
  assign n3510 = ~n44 & ~n3318 ;
  assign n3511 = n2509 & ~n3510 ;
  assign n3512 = ~n954 & n3196 ;
  assign n3513 = n3511 & n3512 ;
  assign n3514 = n418 & n3513 ;
  assign n3515 = ~n3509 & ~n3514 ;
  assign n3516 = x4 & ~n3515 ;
  assign n3517 = x10 & ~n2600 ;
  assign n3518 = x6 & n1165 ;
  assign n3519 = ~n3517 & ~n3518 ;
  assign n3520 = n673 & n2901 ;
  assign n3521 = ~n3519 & n3520 ;
  assign n3522 = n625 & n2816 ;
  assign n3523 = n2561 & n2853 ;
  assign n3524 = ~n3522 & ~n3523 ;
  assign n3525 = ~n3521 & n3524 ;
  assign n3526 = n1536 & ~n3525 ;
  assign n3527 = ~n3516 & ~n3526 ;
  assign n3528 = ~n3505 & n3527 ;
  assign n3529 = ~x12 & ~n3528 ;
  assign n3530 = ~x0 & n2608 ;
  assign n3531 = n1327 & n3530 ;
  assign n3532 = x5 & n2271 ;
  assign n3533 = n2535 & n3532 ;
  assign n3534 = ~n3531 & ~n3533 ;
  assign n3535 = x7 & ~n467 ;
  assign n3536 = ~n3534 & n3535 ;
  assign n3537 = ~n3130 & n3188 ;
  assign n3538 = n1002 & n3537 ;
  assign n3539 = ~n3536 & ~n3538 ;
  assign n3540 = ~x0 & n2557 ;
  assign n3541 = n3188 ^ x5 ;
  assign n3542 = n3541 ^ n3188 ;
  assign n3543 = n3542 ^ n3540 ;
  assign n3544 = n3540 ^ n2823 ;
  assign n3545 = n1407 & ~n3544 ;
  assign n3546 = n3545 ^ n3188 ;
  assign n3547 = ~n3543 & n3546 ;
  assign n3548 = n3547 ^ n3545 ;
  assign n3549 = ~n3540 & n3548 ;
  assign n3550 = n3549 ^ n3545 ;
  assign n3551 = n3550 ^ n3547 ;
  assign n3552 = n3539 & ~n3551 ;
  assign n3553 = ~x14 & n226 ;
  assign n3554 = ~n3552 & n3553 ;
  assign n3555 = ~x13 & n779 ;
  assign n3556 = n175 & n1363 ;
  assign n3557 = n3555 & n3556 ;
  assign n3558 = n2877 & n3557 ;
  assign n3559 = n17 & n3558 ;
  assign n3560 = x14 ^ x11 ;
  assign n3561 = ~x12 & n198 ;
  assign n3562 = n1499 & n2558 ;
  assign n3563 = n3561 & n3562 ;
  assign n3564 = ~x2 & n2608 ;
  assign n3565 = ~x8 & n3564 ;
  assign n3566 = ~n3428 & ~n3565 ;
  assign n3567 = n3540 & ~n3566 ;
  assign n3568 = ~x2 & ~x7 ;
  assign n3569 = n430 & n2608 ;
  assign n3570 = n3568 & n3569 ;
  assign n3571 = ~n3429 & ~n3570 ;
  assign n3572 = n1683 & ~n3571 ;
  assign n3573 = ~n3567 & ~n3572 ;
  assign n3574 = ~n3563 & n3573 ;
  assign n3575 = n3206 & ~n3574 ;
  assign n3576 = n2811 & n3279 ;
  assign n3577 = x12 ^ x7 ;
  assign n3578 = x4 ^ x0 ;
  assign n3579 = x12 ^ x4 ;
  assign n3580 = n3578 & n3579 ;
  assign n3581 = n3580 ^ x4 ;
  assign n3582 = ~n3577 & ~n3581 ;
  assign n3583 = n3576 & n3582 ;
  assign n3584 = n3583 ^ n2036 ;
  assign n3585 = n3584 ^ n3583 ;
  assign n3586 = ~n34 & ~n2562 ;
  assign n3587 = n3467 & ~n3586 ;
  assign n3588 = ~x6 & n2849 ;
  assign n3589 = ~n3587 & ~n3588 ;
  assign n3590 = n784 & ~n3589 ;
  assign n3591 = n3590 ^ n3583 ;
  assign n3592 = n3591 ^ n3583 ;
  assign n3593 = n3585 & n3592 ;
  assign n3594 = n3593 ^ n3583 ;
  assign n3595 = ~x8 & n3594 ;
  assign n3596 = n3595 ^ n3583 ;
  assign n3597 = ~n3575 & ~n3596 ;
  assign n3598 = n3597 ^ x14 ;
  assign n3599 = n3598 ^ n3597 ;
  assign n3600 = n3599 ^ n3560 ;
  assign n3601 = n740 & ~n955 ;
  assign n3602 = n2975 & n3601 ;
  assign n3603 = ~n778 & n1113 ;
  assign n3604 = n3603 ^ x8 ;
  assign n3605 = n3604 ^ n3603 ;
  assign n3606 = n3603 ^ n740 ;
  assign n3607 = n3606 ^ n3603 ;
  assign n3608 = n3605 & n3607 ;
  assign n3609 = n3608 ^ n3603 ;
  assign n3610 = ~x7 & n3609 ;
  assign n3611 = n3610 ^ n3603 ;
  assign n3612 = n2613 & n3611 ;
  assign n3613 = ~n3602 & ~n3612 ;
  assign n3614 = x5 & ~n3613 ;
  assign n3615 = ~n2678 & n2823 ;
  assign n3616 = ~x8 & n3615 ;
  assign n3617 = n827 & n2955 ;
  assign n3618 = ~n3616 & ~n3617 ;
  assign n3619 = n3261 & ~n3618 ;
  assign n3620 = ~n3614 & ~n3619 ;
  assign n3621 = n3620 ^ x12 ;
  assign n3622 = x12 & ~n3621 ;
  assign n3623 = n3622 ^ n3597 ;
  assign n3624 = n3623 ^ x12 ;
  assign n3625 = ~n3600 & ~n3624 ;
  assign n3626 = n3625 ^ n3622 ;
  assign n3627 = n3626 ^ x12 ;
  assign n3628 = n3560 & n3627 ;
  assign n3629 = ~n3559 & ~n3628 ;
  assign n3630 = ~n3554 & n3629 ;
  assign n3631 = ~n3529 & n3630 ;
  assign n3632 = n3631 ^ n3482 ;
  assign n3633 = ~n3484 & ~n3632 ;
  assign n3634 = n3633 ^ n3482 ;
  assign n3635 = n3304 & ~n3634 ;
  assign n3636 = ~n3277 & n3635 ;
  assign n3637 = n55 & ~n3636 ;
  assign n3638 = x8 & n633 ;
  assign n3639 = ~n3464 & n3638 ;
  assign n3640 = n282 & n889 ;
  assign n3641 = n465 & n642 ;
  assign n3642 = ~n3640 & ~n3641 ;
  assign n3643 = n2721 & ~n3642 ;
  assign n3644 = n2466 & n3643 ;
  assign n3645 = ~n3639 & ~n3644 ;
  assign n3646 = ~n230 & n3440 ;
  assign n3647 = n2668 & n3165 ;
  assign n3648 = ~n105 & ~n242 ;
  assign n3649 = n3647 & n3648 ;
  assign n3650 = ~n3646 & ~n3649 ;
  assign n3651 = x10 & ~n3650 ;
  assign n3652 = n2225 & n3258 ;
  assign n3653 = ~n3651 & ~n3652 ;
  assign n3654 = n3653 ^ x5 ;
  assign n3655 = n3654 ^ n3653 ;
  assign n3656 = n3655 ^ n656 ;
  assign n3657 = n248 & n948 ;
  assign n3658 = n230 ^ n105 ;
  assign n3659 = n230 ^ x7 ;
  assign n3660 = n3659 ^ n230 ;
  assign n3661 = n3658 & n3660 ;
  assign n3662 = n3661 ^ n230 ;
  assign n3663 = ~x6 & n3662 ;
  assign n3664 = ~n3657 & ~n3663 ;
  assign n3665 = n2799 & ~n3664 ;
  assign n3666 = x4 & n2806 ;
  assign n3667 = n2957 & n3666 ;
  assign n3668 = n3667 ^ n3665 ;
  assign n3669 = ~n3665 & n3668 ;
  assign n3670 = n3669 ^ n3653 ;
  assign n3671 = n3670 ^ n3665 ;
  assign n3672 = n3656 & ~n3671 ;
  assign n3673 = n3672 ^ n3669 ;
  assign n3674 = n3673 ^ n3665 ;
  assign n3675 = n656 & ~n3674 ;
  assign n3676 = n3675 ^ n656 ;
  assign n3677 = n3645 & ~n3676 ;
  assign n3678 = n742 & ~n3677 ;
  assign n3679 = ~n3637 & ~n3678 ;
  assign n3680 = n981 & n1327 ;
  assign n3681 = n1912 & n3680 ;
  assign n3682 = ~x10 & n2653 ;
  assign n3683 = n1226 & n3682 ;
  assign n3684 = n24 & n3683 ;
  assign n3685 = ~n3681 & ~n3684 ;
  assign n3686 = ~x0 & n318 ;
  assign n3687 = n1581 & n2910 ;
  assign n3688 = n3687 ^ x6 ;
  assign n3689 = n3688 ^ n3687 ;
  assign n3690 = n3687 ^ n1898 ;
  assign n3691 = n3690 ^ n3687 ;
  assign n3692 = ~n3689 & n3691 ;
  assign n3693 = n3692 ^ n3687 ;
  assign n3694 = ~x9 & n3693 ;
  assign n3695 = n3694 ^ n3687 ;
  assign n3696 = n3686 & n3695 ;
  assign n3697 = ~x1 & n224 ;
  assign n3698 = n3564 & n3697 ;
  assign n3699 = n282 & n3698 ;
  assign n3700 = ~n3696 & ~n3699 ;
  assign n3701 = ~n3685 & ~n3700 ;
  assign n3702 = ~x10 & n2959 ;
  assign n3703 = x8 & n1658 ;
  assign n3704 = ~n1407 & ~n2224 ;
  assign n3705 = n2535 & n3704 ;
  assign n3706 = ~n3703 & n3705 ;
  assign n3707 = ~n3702 & ~n3706 ;
  assign n3708 = n3081 & ~n3707 ;
  assign n3709 = n2822 & n3708 ;
  assign n3861 = n3420 ^ n2684 ;
  assign n3862 = n1025 & n1226 ;
  assign n3863 = n489 & n3862 ;
  assign n3864 = n3863 ^ n3861 ;
  assign n3865 = n3864 ^ n3420 ;
  assign n3866 = n3865 ^ n3864 ;
  assign n3867 = n34 & n1010 ;
  assign n3868 = n1255 & n3867 ;
  assign n3869 = n104 & n1226 ;
  assign n3870 = n90 & n3869 ;
  assign n3871 = ~n3868 & ~n3870 ;
  assign n3872 = n3871 ^ n3864 ;
  assign n3873 = n3872 ^ n3861 ;
  assign n3874 = n3866 & n3873 ;
  assign n3875 = n3874 ^ n3871 ;
  assign n3876 = n866 & ~n1703 ;
  assign n3877 = n555 & n3876 ;
  assign n3878 = ~x0 & n1973 ;
  assign n3879 = ~n3877 & ~n3878 ;
  assign n3880 = n3871 & n3879 ;
  assign n3881 = n3880 ^ n3861 ;
  assign n3882 = n3875 & ~n3881 ;
  assign n3883 = n3882 ^ n3880 ;
  assign n3884 = ~n3861 & n3883 ;
  assign n3885 = n3884 ^ n3874 ;
  assign n3886 = n3885 ^ n2684 ;
  assign n3887 = n3886 ^ n3871 ;
  assign n3888 = n24 & n3887 ;
  assign n3889 = n554 & n622 ;
  assign n3890 = n3123 & n3889 ;
  assign n3891 = n1880 & n2708 ;
  assign n3892 = n26 ^ x7 ;
  assign n3893 = n3892 ^ n26 ;
  assign n3894 = ~x5 & ~x6 ;
  assign n3895 = n3894 ^ n26 ;
  assign n3896 = n3893 & n3895 ;
  assign n3897 = n3896 ^ n26 ;
  assign n3898 = n471 & n3897 ;
  assign n3899 = ~n3891 & ~n3898 ;
  assign n3900 = n607 & ~n3899 ;
  assign n3901 = ~n3890 & ~n3900 ;
  assign n3902 = x12 & ~n3901 ;
  assign n3903 = ~x9 & n524 ;
  assign n3904 = ~n2213 & ~n3903 ;
  assign n3905 = n1683 & ~n3904 ;
  assign n3906 = n3147 & n3905 ;
  assign n3907 = n2901 & n3326 ;
  assign n3908 = ~n1618 & ~n2279 ;
  assign n3909 = n2848 & ~n3908 ;
  assign n3910 = ~n3907 & ~n3909 ;
  assign n3911 = n2736 & ~n3910 ;
  assign n3912 = x11 & n3911 ;
  assign n3913 = ~n3906 & ~n3912 ;
  assign n3914 = ~x10 & n1683 ;
  assign n3798 = ~x4 & ~x7 ;
  assign n3915 = n1155 & n3798 ;
  assign n3916 = n3915 ^ x5 ;
  assign n3917 = n3916 ^ n3915 ;
  assign n3918 = n3917 ^ n3914 ;
  assign n3919 = x9 ^ x7 ;
  assign n3920 = x11 & ~n3919 ;
  assign n3921 = n496 ^ x8 ;
  assign n3922 = x9 ^ x6 ;
  assign n3923 = n3922 ^ x8 ;
  assign n3924 = n3923 ^ n3920 ;
  assign n3925 = n3921 & n3924 ;
  assign n3926 = n3925 ^ n496 ;
  assign n3927 = n3920 & n3926 ;
  assign n3928 = n1896 & n3258 ;
  assign n3929 = n3928 ^ n3927 ;
  assign n3930 = ~n3927 & n3929 ;
  assign n3931 = n3930 ^ n3915 ;
  assign n3932 = n3931 ^ n3927 ;
  assign n3933 = ~n3918 & n3932 ;
  assign n3934 = n3933 ^ n3930 ;
  assign n3935 = n3934 ^ n3927 ;
  assign n3936 = n3914 & ~n3935 ;
  assign n3937 = n3936 ^ n3914 ;
  assign n3938 = n3913 & ~n3937 ;
  assign n3939 = ~n3902 & n3938 ;
  assign n3940 = n673 & ~n3939 ;
  assign n3941 = ~n3888 & ~n3940 ;
  assign n3728 = ~x5 & x9 ;
  assign n3751 = n557 & n3165 ;
  assign n3752 = x13 ^ x8 ;
  assign n3753 = n981 & ~n3752 ;
  assign n3754 = ~n3751 & ~n3753 ;
  assign n3755 = n3728 & ~n3754 ;
  assign n3756 = n557 & n948 ;
  assign n3757 = ~n956 & ~n3756 ;
  assign n3758 = n526 & ~n3757 ;
  assign n3759 = ~n3755 & ~n3758 ;
  assign n3760 = n3530 & ~n3759 ;
  assign n3761 = x6 & ~x13 ;
  assign n3762 = ~x7 & ~n3761 ;
  assign n3763 = ~n557 & ~n3762 ;
  assign n3764 = n795 & ~n2693 ;
  assign n3765 = ~n3763 & n3764 ;
  assign n3766 = x8 & n3765 ;
  assign n3767 = ~n473 & ~n2279 ;
  assign n3768 = ~n2557 & ~n2881 ;
  assign n3769 = ~n2684 & n3768 ;
  assign n3770 = ~n3767 & n3769 ;
  assign n3771 = ~n3615 & ~n3770 ;
  assign n3772 = n365 & ~n3771 ;
  assign n3773 = n557 & n3196 ;
  assign n3774 = x10 & ~n3375 ;
  assign n3775 = ~n3773 & ~n3774 ;
  assign n3776 = n2624 & ~n3775 ;
  assign n3777 = n2608 & n2653 ;
  assign n3778 = n889 & n3777 ;
  assign n3779 = ~n3776 & ~n3778 ;
  assign n3780 = ~n3772 & n3779 ;
  assign n3781 = ~n3766 & n3780 ;
  assign n3782 = n2747 & ~n3781 ;
  assign n3783 = n2569 & ~n3490 ;
  assign n3784 = ~n3361 & ~n3783 ;
  assign n3785 = ~x8 & n817 ;
  assign n3786 = n843 & n3783 ;
  assign n3787 = ~n889 & ~n3786 ;
  assign n3788 = n3785 & ~n3787 ;
  assign n3789 = ~n3784 & n3788 ;
  assign n3790 = ~n3782 & ~n3789 ;
  assign n3791 = ~n3760 & n3790 ;
  assign n3792 = n1555 & ~n3791 ;
  assign n3710 = ~x0 & n2560 ;
  assign n3711 = n105 & n2653 ;
  assign n3712 = n151 & ~n2902 ;
  assign n3713 = ~n3711 & ~n3712 ;
  assign n3714 = ~x9 & ~n3713 ;
  assign n3715 = ~x5 & n3657 ;
  assign n3716 = ~n3714 & ~n3715 ;
  assign n3717 = n3710 & ~n3716 ;
  assign n3718 = n24 & n104 ;
  assign n3719 = n2822 & n3718 ;
  assign n3720 = ~x7 & n1920 ;
  assign n3721 = n1905 & n3720 ;
  assign n3722 = n1113 & n3721 ;
  assign n3723 = n817 & n3306 ;
  assign n3724 = ~x14 & n3723 ;
  assign n3725 = ~n3722 & ~n3724 ;
  assign n3726 = ~n3719 & n3725 ;
  assign n3727 = n406 & ~n3726 ;
  assign n3729 = ~n858 & ~n1025 ;
  assign n3730 = x5 & ~n3729 ;
  assign n3731 = ~n3728 & ~n3730 ;
  assign n3732 = x10 & ~n3731 ;
  assign n3733 = n2480 & n3206 ;
  assign n3734 = ~n3732 & ~n3733 ;
  assign n3735 = n151 & n787 ;
  assign n3736 = ~x14 & n3735 ;
  assign n3737 = ~n3734 & n3736 ;
  assign n3738 = ~n3727 & ~n3737 ;
  assign n3739 = ~n3717 & n3738 ;
  assign n3740 = n2608 & ~n3739 ;
  assign n3741 = n106 & n3089 ;
  assign n3742 = ~n3274 & ~n3741 ;
  assign n3743 = x0 & n3490 ;
  assign n3744 = ~n3742 & n3743 ;
  assign n3745 = n497 & n556 ;
  assign n3746 = ~x14 & n1973 ;
  assign n3747 = n3745 & n3746 ;
  assign n3748 = n2633 & n3747 ;
  assign n3749 = ~n3744 & ~n3748 ;
  assign n3750 = ~n3740 & n3749 ;
  assign n3793 = n3792 ^ n3750 ;
  assign n3794 = n3793 ^ n3750 ;
  assign n3795 = ~n45 & ~n2557 ;
  assign n3796 = ~n2599 & ~n2881 ;
  assign n3797 = n3795 & ~n3796 ;
  assign n3799 = n2559 & n2562 ;
  assign n3800 = ~n3798 & n3799 ;
  assign n3801 = ~n3797 & ~n3800 ;
  assign n3802 = n3728 & ~n3801 ;
  assign n3803 = ~n195 & ~n1476 ;
  assign n3804 = ~x9 & ~n2599 ;
  assign n3805 = ~n3803 & ~n3804 ;
  assign n3806 = n1038 & n2848 ;
  assign n3807 = n3805 & n3806 ;
  assign n3808 = ~x9 & n2608 ;
  assign n3809 = n34 & n3808 ;
  assign n3810 = ~n955 & n3809 ;
  assign n3811 = ~n3807 & ~n3810 ;
  assign n3812 = ~n3802 & n3811 ;
  assign n3813 = n466 & ~n3812 ;
  assign n3814 = n2654 & n3530 ;
  assign n3815 = ~n3196 & n3785 ;
  assign n3816 = ~n2703 & n3815 ;
  assign n3817 = ~n3814 & ~n3816 ;
  assign n3818 = n888 & ~n3817 ;
  assign n3819 = n2569 & ~n3130 ;
  assign n3820 = n3819 ^ x13 ;
  assign n3821 = n3819 ^ x6 ;
  assign n3822 = n3821 ^ x6 ;
  assign n3823 = n3361 ^ x6 ;
  assign n3824 = ~n3822 & ~n3823 ;
  assign n3825 = n3824 ^ x6 ;
  assign n3826 = ~n3820 & n3825 ;
  assign n3827 = n3826 ^ x13 ;
  assign n3828 = n1078 & ~n3827 ;
  assign n3829 = ~x9 & n3828 ;
  assign n3830 = ~n3818 & ~n3829 ;
  assign n3831 = ~n3813 & n3830 ;
  assign n3832 = n3307 & ~n3831 ;
  assign n3833 = n299 & n3530 ;
  assign n3834 = ~n2902 & n3833 ;
  assign n3835 = ~x6 & ~x9 ;
  assign n3836 = x5 ^ x0 ;
  assign n3837 = n3836 ^ x7 ;
  assign n3838 = n467 ^ x5 ;
  assign n3839 = ~x5 & n3838 ;
  assign n3840 = n3839 ^ n463 ;
  assign n3841 = n3840 ^ x5 ;
  assign n3842 = n463 ^ x7 ;
  assign n3843 = n3842 ^ x5 ;
  assign n3844 = n3843 ^ n463 ;
  assign n3845 = n3844 ^ n3837 ;
  assign n3846 = ~n3841 & ~n3845 ;
  assign n3847 = n3846 ^ n3839 ;
  assign n3848 = n3847 ^ x5 ;
  assign n3849 = n3837 & ~n3848 ;
  assign n3850 = n3835 & n3849 ;
  assign n3851 = ~x4 & n3850 ;
  assign n3852 = ~n3834 & ~n3851 ;
  assign n3853 = n334 & ~n3852 ;
  assign n3854 = ~n3832 & ~n3853 ;
  assign n3855 = n3854 ^ n3750 ;
  assign n3856 = n3855 ^ n3750 ;
  assign n3857 = ~n3794 & n3856 ;
  assign n3858 = n3857 ^ n3750 ;
  assign n3859 = x12 & n3858 ;
  assign n3860 = n3859 ^ n3750 ;
  assign n3942 = n3941 ^ n3860 ;
  assign n3943 = n3942 ^ n3941 ;
  assign n3944 = n1991 & n2508 ;
  assign n3945 = ~n1136 & n3944 ;
  assign n3946 = n3666 & n3945 ;
  assign n3947 = n1264 & n3946 ;
  assign n3948 = n3947 ^ n3941 ;
  assign n3949 = n3948 ^ n3941 ;
  assign n3950 = n3943 & ~n3949 ;
  assign n3951 = n3950 ^ n3941 ;
  assign n3952 = ~x2 & n3951 ;
  assign n3953 = n3952 ^ n3941 ;
  assign n3954 = ~n3709 & n3953 ;
  assign n3955 = n348 & ~n3954 ;
  assign n3956 = ~n3701 & ~n3955 ;
  assign n3957 = n3679 & n3956 ;
  assign n3958 = ~n3255 & n3957 ;
  assign n3959 = ~x15 & ~n3958 ;
  assign n3960 = ~x14 & ~x15 ;
  assign n3961 = n164 & n2637 ;
  assign n3962 = n828 & n3961 ;
  assign n3963 = ~x7 & n57 ;
  assign n3964 = n1920 & n3963 ;
  assign n3965 = ~n3962 & ~n3964 ;
  assign n3966 = n1104 & ~n3965 ;
  assign n3972 = n2036 & n3196 ;
  assign n3967 = ~x9 & n2458 ;
  assign n3968 = n3490 & n3967 ;
  assign n3969 = n57 & n3968 ;
  assign n3973 = n3972 ^ n3969 ;
  assign n3974 = n3973 ^ n3969 ;
  assign n3970 = n3969 ^ n1169 ;
  assign n3971 = n3970 ^ n3969 ;
  assign n3975 = n3974 ^ n3971 ;
  assign n3976 = n3969 ^ x0 ;
  assign n3977 = n3976 ^ n3969 ;
  assign n3978 = n3977 ^ n3974 ;
  assign n3979 = n3974 & ~n3978 ;
  assign n3980 = n3979 ^ n3974 ;
  assign n3981 = n3975 & n3980 ;
  assign n3982 = n3981 ^ n3979 ;
  assign n3983 = n3982 ^ n3969 ;
  assign n3984 = n3983 ^ n3974 ;
  assign n3985 = x11 & n3984 ;
  assign n3986 = n3985 ^ n3969 ;
  assign n3987 = ~n3966 & ~n3986 ;
  assign n3988 = ~n3960 & ~n3987 ;
  assign n3989 = ~n1382 & n2286 ;
  assign n3990 = ~n19 & ~n863 ;
  assign n3991 = n3989 & n3990 ;
  assign n3992 = ~n306 & ~n874 ;
  assign n3993 = n311 & n3992 ;
  assign n3994 = ~n126 & ~n3993 ;
  assign n3995 = n2564 & ~n3994 ;
  assign n3996 = ~n3991 & ~n3995 ;
  assign n3997 = n311 & n2564 ;
  assign n3998 = ~n19 & n3997 ;
  assign n3999 = ~x0 & ~n3998 ;
  assign n4000 = n3682 & ~n3999 ;
  assign n4001 = ~n3996 & n4000 ;
  assign n4002 = x5 & n363 ;
  assign n4003 = n261 & n4002 ;
  assign n4004 = n833 & n4003 ;
  assign n4005 = n1284 & ~n1327 ;
  assign n4006 = n261 & n4005 ;
  assign n4007 = ~x0 & n700 ;
  assign n4008 = n1214 & n4007 ;
  assign n4009 = ~n4006 & ~n4008 ;
  assign n4010 = n329 & ~n4009 ;
  assign n4011 = n2480 & n4010 ;
  assign n4012 = ~n4004 & ~n4011 ;
  assign n4013 = ~x1 & n2653 ;
  assign n4014 = x1 & ~x7 ;
  assign n4015 = ~x5 & x15 ;
  assign n4016 = n4014 & n4015 ;
  assign n4017 = ~n4013 & ~n4016 ;
  assign n4018 = n3914 & ~n4017 ;
  assign n4019 = ~x1 & n1423 ;
  assign n4020 = n34 & n4019 ;
  assign n4021 = ~n4018 & ~n4020 ;
  assign n4022 = n1565 & ~n4021 ;
  assign n4023 = n1270 & n1682 ;
  assign n4024 = n104 & n4023 ;
  assign n4025 = n4013 & n4024 ;
  assign n4026 = ~x14 & n1241 ;
  assign n4027 = ~x0 & n568 ;
  assign n4028 = n4026 & n4027 ;
  assign n4029 = n3294 & n4028 ;
  assign n4030 = ~n4025 & ~n4029 ;
  assign n4031 = ~n4022 & n4030 ;
  assign n4032 = ~n869 & ~n4031 ;
  assign n4033 = ~x11 & n1214 ;
  assign n4034 = ~n1955 & n4033 ;
  assign n4035 = ~x12 & n311 ;
  assign n4036 = n109 & n4035 ;
  assign n4037 = ~n1113 & n4036 ;
  assign n4038 = ~n4034 & ~n4037 ;
  assign n4039 = n2675 & ~n4038 ;
  assign n4040 = x12 & n3196 ;
  assign n4041 = ~n395 & n978 ;
  assign n4042 = n4041 ^ n700 ;
  assign n4043 = n4042 ^ n4040 ;
  assign n4044 = n1952 ^ n19 ;
  assign n4045 = n4044 ^ n4042 ;
  assign n4046 = ~n4041 & ~n4045 ;
  assign n4047 = n4046 ^ n19 ;
  assign n4048 = n4047 ^ n4041 ;
  assign n4049 = n4048 ^ n4042 ;
  assign n4050 = n4049 ^ n4040 ;
  assign n4051 = n4043 & n4050 ;
  assign n4052 = n4051 ^ n4046 ;
  assign n4053 = n4052 ^ n19 ;
  assign n4054 = n4053 ^ n4042 ;
  assign n4055 = n4040 & ~n4054 ;
  assign n4056 = n4055 ^ n4040 ;
  assign n4057 = n4056 ^ n4040 ;
  assign n4058 = ~n4039 & ~n4057 ;
  assign n4059 = ~x10 & ~n4058 ;
  assign n4060 = ~n4032 & ~n4059 ;
  assign n4061 = n4012 & n4060 ;
  assign n4062 = ~n4001 & n4061 ;
  assign n4063 = ~n3988 & n4062 ;
  assign n4064 = ~x3 & ~n4063 ;
  assign n4065 = n306 & n3294 ;
  assign n4066 = n66 & n2675 ;
  assign n4067 = ~n4065 & ~n4066 ;
  assign n4068 = n1240 & ~n4067 ;
  assign n4069 = x7 & n89 ;
  assign n4070 = n2389 & n4069 ;
  assign n4071 = n4070 ^ n4068 ;
  assign n4072 = n45 & n2654 ;
  assign n4073 = ~x7 & n571 ;
  assign n4074 = ~n438 & ~n870 ;
  assign n4075 = n4073 & ~n4074 ;
  assign n4076 = ~n105 & ~n346 ;
  assign n4077 = n2822 & ~n4076 ;
  assign n4078 = ~n4075 & ~n4077 ;
  assign n4079 = ~n4072 & n4078 ;
  assign n4080 = n700 & ~n4079 ;
  assign n4081 = ~n396 & n2282 ;
  assign n4082 = n248 & n4081 ;
  assign n4083 = n3196 & n4082 ;
  assign n4084 = ~n4080 & ~n4083 ;
  assign n4085 = n4084 ^ x12 ;
  assign n4086 = n4085 ^ n4084 ;
  assign n4087 = n240 & n1270 ;
  assign n4088 = ~n2738 & ~n4087 ;
  assign n4089 = n4088 ^ n555 ;
  assign n4090 = n4089 ^ n555 ;
  assign n4091 = n555 ^ x5 ;
  assign n4092 = n4091 ^ n555 ;
  assign n4093 = ~n4090 & n4092 ;
  assign n4094 = n4093 ^ n555 ;
  assign n4095 = ~x0 & ~n4094 ;
  assign n4096 = n4095 ^ n555 ;
  assign n4097 = n1042 & ~n4096 ;
  assign n4098 = x13 & ~n1270 ;
  assign n4099 = x11 & n4098 ;
  assign n4100 = n396 & ~n4099 ;
  assign n4101 = n3196 & ~n4100 ;
  assign n4102 = ~x14 & ~n290 ;
  assign n4103 = n2329 & ~n4102 ;
  assign n4104 = n240 & ~n395 ;
  assign n4105 = ~n4103 & ~n4104 ;
  assign n4106 = n4105 ^ n197 ;
  assign n4107 = n4105 ^ x0 ;
  assign n4108 = n4107 ^ n4105 ;
  assign n4109 = n4108 ^ n4101 ;
  assign n4110 = n4109 ^ n4100 ;
  assign n4111 = ~n4106 & ~n4110 ;
  assign n4112 = n4111 ^ n4105 ;
  assign n4113 = n4101 & ~n4112 ;
  assign n4114 = n4113 ^ n4101 ;
  assign n4115 = n4114 ^ n3196 ;
  assign n4116 = x0 & n749 ;
  assign n4117 = n3728 & n4116 ;
  assign n4118 = n159 & n2633 ;
  assign n4119 = n4118 ^ x11 ;
  assign n4120 = n4119 ^ n4118 ;
  assign n4121 = n4120 ^ n4117 ;
  assign n4122 = n858 ^ n89 ;
  assign n4123 = n858 & n4122 ;
  assign n4124 = n4123 ^ n4118 ;
  assign n4125 = n4124 ^ n858 ;
  assign n4126 = n4121 & n4125 ;
  assign n4127 = n4126 ^ n4123 ;
  assign n4128 = n4127 ^ n858 ;
  assign n4129 = ~n4117 & n4128 ;
  assign n4130 = n4129 ^ n4117 ;
  assign n4131 = ~n4115 & ~n4130 ;
  assign n4132 = ~n4097 & n4131 ;
  assign n4133 = n4132 ^ n4084 ;
  assign n4134 = n4086 & n4133 ;
  assign n4135 = n4134 ^ n4084 ;
  assign n4136 = n4135 ^ n4068 ;
  assign n4137 = n4071 & ~n4136 ;
  assign n4138 = n4137 ^ n4134 ;
  assign n4139 = n4138 ^ n4084 ;
  assign n4140 = n4139 ^ n4070 ;
  assign n4141 = ~n4068 & ~n4140 ;
  assign n4142 = n4141 ^ n4068 ;
  assign n4143 = n529 & n4142 ;
  assign n4144 = ~n4064 & ~n4143 ;
  assign n4145 = n306 & n845 ;
  assign n4146 = n66 & n524 ;
  assign n4147 = ~n4145 & ~n4146 ;
  assign n4148 = ~n870 & ~n4147 ;
  assign n4149 = n489 & n530 ;
  assign n4150 = n748 & n4149 ;
  assign n4151 = ~n4148 & ~n4150 ;
  assign n4152 = n3408 & ~n4151 ;
  assign n4153 = ~x12 & n524 ;
  assign n4154 = ~n4033 & ~n4153 ;
  assign n4155 = ~n473 & ~n4154 ;
  assign n4156 = ~n633 & ~n2508 ;
  assign n4157 = ~x0 & n4156 ;
  assign n4158 = n196 & n1042 ;
  assign n4159 = ~n817 & n1270 ;
  assign n4160 = ~n274 & ~n4159 ;
  assign n4161 = n4158 & ~n4160 ;
  assign n4162 = ~n4157 & n4161 ;
  assign n4163 = n395 & n2653 ;
  assign n4164 = ~n68 & ~n2991 ;
  assign n4165 = n4163 & n4164 ;
  assign n4166 = ~x7 & x15 ;
  assign n4167 = ~x5 & n4166 ;
  assign n4168 = n348 & n434 ;
  assign n4169 = ~x14 & n4168 ;
  assign n4170 = ~n60 & ~n2568 ;
  assign n4171 = x9 & ~n4170 ;
  assign n4172 = ~n56 & n4171 ;
  assign n4173 = ~n4169 & ~n4172 ;
  assign n4174 = n4167 & ~n4173 ;
  assign n4175 = ~n4165 & ~n4174 ;
  assign n4176 = ~n4162 & n4175 ;
  assign n4177 = n4155 & ~n4176 ;
  assign n4178 = ~n4152 & ~n4177 ;
  assign n4179 = n889 & n1282 ;
  assign n4180 = n1954 & n4179 ;
  assign n4181 = n489 & n1977 ;
  assign n4182 = x12 & n371 ;
  assign n4183 = n76 & n3914 ;
  assign n4184 = ~n4182 & ~n4183 ;
  assign n4185 = ~n4181 & n4184 ;
  assign n4186 = n109 & ~n4185 ;
  assign n4187 = ~n4180 & ~n4186 ;
  assign n4188 = n3196 & ~n4187 ;
  assign n4189 = n4013 & n4179 ;
  assign n4190 = ~n19 & ~n462 ;
  assign n4191 = ~n2607 & ~n4190 ;
  assign n4192 = ~n28 & n1010 ;
  assign n4193 = n4040 & ~n4192 ;
  assign n4194 = n4191 & n4193 ;
  assign n4195 = n1010 & n3196 ;
  assign n4196 = ~x1 & n1282 ;
  assign n4197 = n4195 & n4196 ;
  assign n4198 = ~n4194 & ~n4197 ;
  assign n4199 = ~n4189 & n4198 ;
  assign n4200 = n2747 & ~n4199 ;
  assign n4201 = ~n2607 & ~n3960 ;
  assign n4202 = n109 & n4201 ;
  assign n4203 = x14 & n568 ;
  assign n4204 = ~x11 & n4203 ;
  assign n4205 = ~n4202 & ~n4204 ;
  assign n4206 = ~x9 & n727 ;
  assign n4207 = n4040 & n4206 ;
  assign n4208 = ~n4205 & n4207 ;
  assign n4209 = ~n4200 & ~n4208 ;
  assign n4210 = ~n4188 & n4209 ;
  assign n4211 = n2653 & n3418 ;
  assign n4212 = n4211 ^ x1 ;
  assign n4213 = n4211 ^ x13 ;
  assign n4214 = n4213 ^ x13 ;
  assign n4215 = ~n1423 & ~n2312 ;
  assign n4216 = n3196 & ~n4215 ;
  assign n4217 = n4216 ^ x13 ;
  assign n4218 = ~n4214 & ~n4217 ;
  assign n4219 = n4218 ^ x13 ;
  assign n4220 = n4212 & n4219 ;
  assign n4221 = n4220 ^ x1 ;
  assign n4222 = ~x10 & n260 ;
  assign n4223 = n126 & n3196 ;
  assign n4224 = n4222 & n4223 ;
  assign n4225 = ~n1656 & ~n2607 ;
  assign n4226 = ~x1 & n3196 ;
  assign n4227 = n4225 & n4226 ;
  assign n4228 = n1423 ^ x1 ;
  assign n4229 = n1423 ^ x14 ;
  assign n4230 = n4229 ^ x14 ;
  assign n4231 = n511 & n1282 ;
  assign n4232 = n4231 ^ x14 ;
  assign n4233 = ~n4230 & ~n4232 ;
  assign n4234 = n4233 ^ x14 ;
  assign n4235 = n4228 & n4234 ;
  assign n4236 = n4235 ^ x1 ;
  assign n4237 = n4236 ^ x13 ;
  assign n4238 = n4237 ^ n4236 ;
  assign n4239 = n4238 ^ n2653 ;
  assign n4240 = ~n1656 & ~n2466 ;
  assign n4241 = n568 & ~n3030 ;
  assign n4242 = n4241 ^ n4240 ;
  assign n4243 = n4240 & ~n4242 ;
  assign n4244 = n4243 ^ n4236 ;
  assign n4245 = n4244 ^ n4240 ;
  assign n4246 = ~n4239 & n4245 ;
  assign n4247 = n4246 ^ n4243 ;
  assign n4248 = n4247 ^ n4240 ;
  assign n4249 = n2653 & n4248 ;
  assign n4250 = ~n4227 & ~n4249 ;
  assign n4251 = n4250 ^ x11 ;
  assign n4252 = n4251 ^ n4250 ;
  assign n4253 = ~x1 & ~x7 ;
  assign n4254 = n889 & n4253 ;
  assign n4255 = n2873 & n4254 ;
  assign n4256 = n4255 ^ n4250 ;
  assign n4257 = n4252 & ~n4256 ;
  assign n4258 = n4257 ^ n4250 ;
  assign n4259 = ~n4224 & n4258 ;
  assign n4260 = ~n4221 & n4259 ;
  assign n4261 = n434 & ~n4260 ;
  assign n4262 = ~x1 & n845 ;
  assign n4263 = n3030 & n4262 ;
  assign n4264 = n2654 & n4263 ;
  assign n4265 = ~n4261 & ~n4264 ;
  assign n4266 = n4210 & n4265 ;
  assign n4267 = x3 & ~n4266 ;
  assign n4295 = n311 & n557 ;
  assign n4296 = ~n4182 & ~n4295 ;
  assign n4268 = n828 & n978 ;
  assign n4269 = n489 & n1247 ;
  assign n4270 = ~n4268 & ~n4269 ;
  assign n4271 = ~n240 & ~n1226 ;
  assign n4272 = ~n863 & ~n4271 ;
  assign n4273 = ~n525 & ~n4272 ;
  assign n4274 = n60 & ~n4273 ;
  assign n4275 = ~n1062 & ~n1328 ;
  assign n4276 = n414 & n1671 ;
  assign n4277 = n4275 & ~n4276 ;
  assign n4278 = n2282 & ~n4277 ;
  assign n4279 = ~n4274 & ~n4278 ;
  assign n4280 = x10 & ~n2290 ;
  assign n4281 = x0 & n4280 ;
  assign n4282 = n762 & n1214 ;
  assign n4283 = ~n4281 & ~n4282 ;
  assign n4284 = n4279 & n4283 ;
  assign n4285 = n4270 & n4284 ;
  assign n4297 = n4296 ^ n4285 ;
  assign n4286 = ~x12 & n1905 ;
  assign n4287 = ~n986 & n4286 ;
  assign n4288 = ~n24 & n1423 ;
  assign n4289 = ~n4287 & ~n4288 ;
  assign n4290 = x0 & ~n4289 ;
  assign n4291 = ~n381 & ~n473 ;
  assign n4292 = n4035 & ~n4291 ;
  assign n4293 = ~n4290 & ~n4292 ;
  assign n4294 = n4293 ^ n4285 ;
  assign n4298 = n4297 ^ n4294 ;
  assign n4299 = n4294 ^ x11 ;
  assign n4300 = n4299 ^ n4294 ;
  assign n4301 = n4298 & n4300 ;
  assign n4302 = n4301 ^ n4294 ;
  assign n4303 = ~x1 & n4302 ;
  assign n4304 = n4303 ^ n4285 ;
  assign n4305 = n2653 & ~n4304 ;
  assign n4306 = n122 & n4288 ;
  assign n4307 = n900 & n4023 ;
  assign n4308 = ~n869 & n4307 ;
  assign n4309 = n700 & n1683 ;
  assign n4310 = n2735 & n4309 ;
  assign n4311 = ~n4308 & ~n4310 ;
  assign n4312 = n66 & n3462 ;
  assign n4313 = ~x10 & n57 ;
  assign n4314 = ~x11 & n2282 ;
  assign n4315 = n4313 & n4314 ;
  assign n4316 = ~n4312 & ~n4315 ;
  assign n4317 = n311 & n828 ;
  assign n4318 = ~n1214 & ~n4317 ;
  assign n4319 = n4145 & ~n4318 ;
  assign n4320 = n4316 & ~n4319 ;
  assign n4321 = n4311 & n4320 ;
  assign n4322 = ~n4306 & n4321 ;
  assign n4323 = n3196 & ~n4322 ;
  assign n4324 = ~n4305 & ~n4323 ;
  assign n4325 = n375 & ~n4324 ;
  assign n4326 = ~n4267 & ~n4325 ;
  assign n4327 = n4178 & n4326 ;
  assign n4328 = n4144 & n4327 ;
  assign n4329 = n111 & ~n4328 ;
  assign n4330 = ~x2 & n1233 ;
  assign n4331 = ~x5 & n981 ;
  assign n4332 = n105 & n558 ;
  assign n4333 = ~n348 & ~n442 ;
  assign n4334 = n788 & n4333 ;
  assign n4335 = ~n4332 & ~n4334 ;
  assign n4336 = n4331 & ~n4335 ;
  assign n4337 = x14 & n4336 ;
  assign n4338 = ~x3 & x7 ;
  assign n4339 = ~x1 & x15 ;
  assign n4340 = ~x1 & ~n4339 ;
  assign n4341 = n75 & ~n4340 ;
  assign n4342 = n623 & n4341 ;
  assign n4343 = n4338 & n4342 ;
  assign n4344 = ~x3 & n2653 ;
  assign n4345 = x1 & ~x15 ;
  assign n4346 = ~n700 & ~n4345 ;
  assign n4347 = n4344 & n4346 ;
  assign n4348 = n978 & n4347 ;
  assign n4349 = ~x11 & n3196 ;
  assign n4350 = x1 & x15 ;
  assign n4351 = ~x14 & n4350 ;
  assign n4352 = ~n261 & ~n4351 ;
  assign n4353 = n4349 & ~n4352 ;
  assign n4354 = ~x3 & n4353 ;
  assign n4355 = ~n4348 & ~n4354 ;
  assign n4356 = n38 & n2653 ;
  assign n4357 = n623 & n4356 ;
  assign n4358 = n363 & n2280 ;
  assign n4359 = ~x7 & n561 ;
  assign n4360 = ~n4358 & ~n4359 ;
  assign n4361 = n4116 & ~n4360 ;
  assign n4362 = ~n4357 & ~n4361 ;
  assign n4363 = n4355 & n4362 ;
  assign n4364 = ~n4343 & n4363 ;
  assign n4365 = ~x13 & ~n4364 ;
  assign n4366 = n1611 & n3091 ;
  assign n4367 = n462 & n4366 ;
  assign n4368 = ~x5 & n2467 ;
  assign n4369 = n55 & n4368 ;
  assign n4370 = n3196 ^ n2653 ;
  assign n4371 = n2653 ^ x11 ;
  assign n4372 = n4371 ^ n2653 ;
  assign n4373 = n4370 & n4372 ;
  assign n4374 = n4373 ^ n2653 ;
  assign n4375 = ~n1149 & n4374 ;
  assign n4376 = ~x1 & n4375 ;
  assign n4377 = ~n4369 & ~n4376 ;
  assign n4378 = n4377 ^ n2568 ;
  assign n4379 = n4377 ^ n60 ;
  assign n4380 = n4379 ^ n60 ;
  assign n4381 = n4380 ^ n4378 ;
  assign n4382 = n4349 ^ n348 ;
  assign n4383 = n4349 & n4382 ;
  assign n4384 = n4383 ^ n60 ;
  assign n4385 = n4384 ^ n4349 ;
  assign n4386 = ~n4381 & ~n4385 ;
  assign n4387 = n4386 ^ n4383 ;
  assign n4388 = n4387 ^ n4349 ;
  assign n4389 = ~n4378 & n4388 ;
  assign n4390 = n4389 ^ n4377 ;
  assign n4391 = n145 & ~n4390 ;
  assign n4392 = x7 & n1435 ;
  assign n4393 = n3092 ^ x3 ;
  assign n4394 = n4393 ^ n3092 ;
  assign n4395 = n4394 ^ n4392 ;
  assign n4396 = n4368 ^ x13 ;
  assign n4397 = n4368 & n4396 ;
  assign n4398 = n4397 ^ n3092 ;
  assign n4399 = n4398 ^ n4368 ;
  assign n4400 = ~n4395 & n4399 ;
  assign n4401 = n4400 ^ n4397 ;
  assign n4402 = n4401 ^ n4368 ;
  assign n4403 = ~n4392 & n4402 ;
  assign n4404 = n4403 ^ n4392 ;
  assign n4405 = n306 & n4404 ;
  assign n4406 = ~n4391 & ~n4405 ;
  assign n4407 = ~n4367 & n4406 ;
  assign n4408 = ~n4365 & n4407 ;
  assign n4409 = x10 & ~n4408 ;
  assign n4410 = x3 & n2282 ;
  assign n4411 = ~x11 & n2653 ;
  assign n4412 = ~n3773 & ~n4411 ;
  assign n4413 = n4410 & ~n4412 ;
  assign n4414 = ~x1 & n4413 ;
  assign n4415 = n38 & n3196 ;
  assign n4416 = n623 & n874 ;
  assign n4417 = n4415 & n4416 ;
  assign n4418 = n4166 & n4222 ;
  assign n4419 = n1958 & n4418 ;
  assign n4420 = x13 & n4419 ;
  assign n4421 = n66 & n652 ;
  assign n4422 = ~n29 & ~n690 ;
  assign n4423 = n978 & ~n4422 ;
  assign n4424 = ~n4007 & ~n4423 ;
  assign n4425 = ~x3 & ~n4424 ;
  assign n4426 = ~n4421 & ~n4425 ;
  assign n4427 = n511 & ~n4426 ;
  assign n4428 = n348 & n866 ;
  assign n4429 = n4428 ^ x10 ;
  assign n4430 = n4429 ^ x11 ;
  assign n4437 = n4430 ^ n4429 ;
  assign n4432 = n749 & n1172 ;
  assign n4431 = n4430 ^ n4428 ;
  assign n4433 = n4432 ^ n4431 ;
  assign n4434 = n4432 ^ n4430 ;
  assign n4435 = n4434 ^ n4429 ;
  assign n4436 = ~n4433 & n4435 ;
  assign n4438 = n4437 ^ n4436 ;
  assign n4439 = ~n306 & n4333 ;
  assign n4440 = n4439 ^ n4430 ;
  assign n4441 = ~n4437 & ~n4440 ;
  assign n4442 = n4441 ^ n4439 ;
  assign n4443 = ~n4438 & n4442 ;
  assign n4444 = n4443 ^ n4436 ;
  assign n4445 = n4444 ^ n4430 ;
  assign n4446 = n4445 ^ x10 ;
  assign n4447 = n4446 ^ n4429 ;
  assign n4448 = ~n4427 & n4447 ;
  assign n4449 = n3306 & ~n4448 ;
  assign n4450 = ~n4420 & ~n4449 ;
  assign n4451 = ~n4417 & n4450 ;
  assign n4452 = ~n4414 & n4451 ;
  assign n4453 = ~n4409 & n4452 ;
  assign n4454 = n4453 ^ x9 ;
  assign n4455 = n4454 ^ n4453 ;
  assign n4456 = n4455 ^ n4337 ;
  assign n4457 = n524 & n3196 ;
  assign n4458 = n442 & n4457 ;
  assign n4459 = n1227 & n4458 ;
  assign n4460 = n405 & n4392 ;
  assign n4461 = x7 & n168 ;
  assign n4462 = ~x7 & n1464 ;
  assign n4463 = n511 & n4462 ;
  assign n4464 = ~n4461 & ~n4463 ;
  assign n4465 = n260 & ~n4464 ;
  assign n4466 = ~n4460 & ~n4465 ;
  assign n4467 = n126 & ~n4466 ;
  assign n4468 = n28 & n2803 ;
  assign n4469 = n4331 & n4468 ;
  assign n4470 = ~x7 & ~x10 ;
  assign n4471 = ~x11 & n4470 ;
  assign n4472 = n4471 ^ n4412 ;
  assign n4473 = n4472 ^ n4412 ;
  assign n4474 = n4412 ^ x5 ;
  assign n4475 = n4474 ^ n4412 ;
  assign n4476 = n4473 & ~n4475 ;
  assign n4477 = n4476 ^ n4412 ;
  assign n4478 = x3 & ~n4477 ;
  assign n4479 = n4478 ^ n4412 ;
  assign n4480 = n690 & ~n4479 ;
  assign n4481 = ~n4469 & ~n4480 ;
  assign n4482 = ~n4467 & n4481 ;
  assign n4483 = ~n4459 & n4482 ;
  assign n4484 = n4483 ^ x0 ;
  assign n4485 = ~n4483 & ~n4484 ;
  assign n4486 = n4485 ^ n4453 ;
  assign n4487 = n4486 ^ n4483 ;
  assign n4488 = ~n4456 & n4487 ;
  assign n4489 = n4488 ^ n4485 ;
  assign n4490 = n4489 ^ n4483 ;
  assign n4491 = ~n4337 & ~n4490 ;
  assign n4492 = n4491 ^ n4337 ;
  assign n4493 = n4330 & n4492 ;
  assign n4494 = x13 & n623 ;
  assign n4495 = n55 & n2675 ;
  assign n4496 = n4494 & n4495 ;
  assign n4497 = ~x9 & n4087 ;
  assign n4498 = n38 & ~n919 ;
  assign n4499 = n4497 & n4498 ;
  assign n4500 = n2902 & n4499 ;
  assign n4501 = ~n4496 & ~n4500 ;
  assign n4502 = ~n3305 & ~n4501 ;
  assign n4503 = n240 & n4158 ;
  assign n4504 = n2467 & n4015 ;
  assign n4505 = n673 & n4504 ;
  assign n4506 = n76 & n4411 ;
  assign n4507 = ~n4505 & ~n4506 ;
  assign n4508 = n4333 & ~n4507 ;
  assign n4509 = ~n4503 & ~n4508 ;
  assign n4510 = n269 & ~n4509 ;
  assign n4511 = ~x9 & n4510 ;
  assign n4512 = ~n4502 & ~n4511 ;
  assign n4513 = ~x2 & n798 ;
  assign n4514 = ~n4411 & ~n4504 ;
  assign n4515 = n55 & ~n4514 ;
  assign n4516 = n414 & n4356 ;
  assign n4517 = ~n4515 & ~n4516 ;
  assign n4518 = n4517 ^ x13 ;
  assign n4519 = n4518 ^ n4517 ;
  assign n4520 = n4519 ^ n4513 ;
  assign n4521 = n55 & n2653 ;
  assign n4522 = n4513 ^ n427 ;
  assign n4523 = n4521 & ~n4522 ;
  assign n4524 = n4523 ^ n4517 ;
  assign n4525 = ~n4520 & ~n4524 ;
  assign n4526 = n4525 ^ n4523 ;
  assign n4527 = ~n4513 & n4526 ;
  assign n4528 = n4527 ^ n4523 ;
  assign n4529 = n4528 ^ n4525 ;
  assign n4530 = n105 & n3196 ;
  assign n4531 = ~x11 & n2841 ;
  assign n4532 = ~n4530 & ~n4531 ;
  assign n4533 = n702 & ~n4532 ;
  assign n4534 = n217 & n497 ;
  assign n4535 = ~n142 & n4534 ;
  assign n4536 = x7 & n4535 ;
  assign n4537 = ~n4533 & ~n4536 ;
  assign n4538 = n274 & ~n4537 ;
  assign n4539 = n4538 ^ x8 ;
  assign n4540 = n4539 ^ n4538 ;
  assign n4541 = n4540 ^ n4529 ;
  assign n4542 = x15 & n105 ;
  assign n4543 = n1990 & n4542 ;
  assign n4544 = n65 & n788 ;
  assign n4545 = n240 & n306 ;
  assign n4546 = n38 & n4542 ;
  assign n4547 = ~n4545 & ~n4546 ;
  assign n4548 = ~x2 & ~n4547 ;
  assign n4549 = ~n4544 & ~n4548 ;
  assign n4550 = ~n4543 & n4549 ;
  assign n4551 = n4550 ^ n2653 ;
  assign n4552 = ~n4550 & ~n4551 ;
  assign n4553 = n4552 ^ n4538 ;
  assign n4554 = n4553 ^ n4550 ;
  assign n4555 = ~n4541 & ~n4554 ;
  assign n4556 = n4555 ^ n4552 ;
  assign n4557 = n4556 ^ n4550 ;
  assign n4558 = ~n4529 & ~n4557 ;
  assign n4559 = n4558 ^ n4529 ;
  assign n4560 = n633 & n4559 ;
  assign n4561 = ~x7 & n79 ;
  assign n4562 = ~n4002 & ~n4561 ;
  assign n4563 = n3686 & ~n4562 ;
  assign n4564 = n240 & n4563 ;
  assign n4565 = x1 & n928 ;
  assign n4566 = ~n644 & n4565 ;
  assign n4567 = ~n650 & ~n659 ;
  assign n4568 = n4002 & n4567 ;
  assign n4569 = n4566 & n4568 ;
  assign n4570 = n25 & n311 ;
  assign n4571 = n4530 & n4570 ;
  assign n4572 = ~x15 & n25 ;
  assign n4573 = n4002 & ~n4572 ;
  assign n4574 = n224 & n3196 ;
  assign n4575 = ~n4573 & ~n4574 ;
  assign n4576 = n240 & ~n4575 ;
  assign n4577 = ~n4571 & ~n4576 ;
  assign n4578 = n74 & ~n4577 ;
  assign n4579 = ~n4569 & ~n4578 ;
  assign n4580 = ~n4564 & n4579 ;
  assign n4581 = n263 & ~n4580 ;
  assign n4582 = ~x5 & n948 ;
  assign n4583 = n4582 ^ x14 ;
  assign n4584 = n4583 ^ n4088 ;
  assign n4585 = n4584 ^ n4582 ;
  assign n4586 = n4585 ^ n4584 ;
  assign n4587 = n503 & n4392 ;
  assign n4588 = ~x8 & n2653 ;
  assign n4589 = ~n986 & n4588 ;
  assign n4590 = ~n2739 & n4589 ;
  assign n4591 = ~n4587 & ~n4590 ;
  assign n4592 = n4591 ^ n4584 ;
  assign n4593 = n4592 ^ n4583 ;
  assign n4594 = n4586 & ~n4593 ;
  assign n4595 = n4594 ^ n4591 ;
  assign n4596 = ~n1949 & n4591 ;
  assign n4597 = n4596 ^ n4583 ;
  assign n4598 = n4595 & ~n4597 ;
  assign n4599 = n4598 ^ n4596 ;
  assign n4600 = ~n4583 & n4599 ;
  assign n4601 = n4600 ^ n4594 ;
  assign n4602 = n4601 ^ x14 ;
  assign n4603 = n4602 ^ n4591 ;
  assign n4604 = n742 & n4603 ;
  assign n4605 = n517 & n718 ;
  assign n4606 = n4356 & n4605 ;
  assign n4607 = ~n75 & n2902 ;
  assign n4608 = n270 & n4087 ;
  assign n4609 = n4607 & n4608 ;
  assign n4610 = ~n4606 & ~n4609 ;
  assign n4611 = ~n850 & ~n4610 ;
  assign n4612 = ~x8 & n442 ;
  assign n4613 = n145 & n4002 ;
  assign n4614 = n4613 ^ x0 ;
  assign n4615 = n4614 ^ n517 ;
  assign n4616 = n213 & n2678 ;
  assign n4617 = n4616 ^ x2 ;
  assign n4618 = x0 & ~n4617 ;
  assign n4619 = n4618 ^ x2 ;
  assign n4620 = n4615 & n4619 ;
  assign n4621 = n4620 ^ n4618 ;
  assign n4622 = n4621 ^ x2 ;
  assign n4623 = n4622 ^ x0 ;
  assign n4624 = n517 & n4623 ;
  assign n4625 = n4612 & n4624 ;
  assign n4626 = ~n4611 & ~n4625 ;
  assign n4627 = n442 & ~n741 ;
  assign n4628 = x8 & n2653 ;
  assign n4629 = ~n4088 & n4628 ;
  assign n4630 = ~n4087 & ~n4494 ;
  assign n4631 = n3294 & ~n4630 ;
  assign n4632 = n3256 & n3728 ;
  assign n4633 = n105 & n4632 ;
  assign n4634 = n4166 & n4633 ;
  assign n4635 = ~n4631 & ~n4634 ;
  assign n4636 = ~n4629 & n4635 ;
  assign n4637 = n4627 & ~n4636 ;
  assign n4638 = n4626 & ~n4637 ;
  assign n4639 = ~n4604 & n4638 ;
  assign n4640 = ~n4581 & n4639 ;
  assign n4641 = ~n4560 & n4640 ;
  assign n4642 = n4512 & n4641 ;
  assign n4643 = ~n1658 & ~n4642 ;
  assign n4644 = ~x2 & n1909 ;
  assign n4645 = n38 & n290 ;
  assign n4646 = n525 & n4645 ;
  assign n4647 = ~x9 & n442 ;
  assign n4648 = n474 & n4647 ;
  assign n4649 = ~n427 & ~n524 ;
  assign n4650 = n348 & n404 ;
  assign n4651 = ~n4649 & n4650 ;
  assign n4652 = ~n4648 & ~n4651 ;
  assign n4653 = x0 & ~n4652 ;
  assign n4654 = ~n4646 & ~n4653 ;
  assign n4655 = n2653 & ~n4654 ;
  assign n4656 = ~x12 & x15 ;
  assign n4657 = n196 & n858 ;
  assign n4658 = n462 & n875 ;
  assign n4659 = n371 ^ n19 ;
  assign n4660 = n4659 ^ n19 ;
  assign n4661 = n4660 ^ x11 ;
  assign n4662 = n381 ^ x1 ;
  assign n4663 = x1 & ~n4662 ;
  assign n4664 = n4663 ^ n19 ;
  assign n4665 = n4664 ^ x1 ;
  assign n4666 = ~n4661 & n4665 ;
  assign n4667 = n4666 ^ n4663 ;
  assign n4668 = n4667 ^ x1 ;
  assign n4669 = x11 & n4668 ;
  assign n4670 = ~n4658 & ~n4669 ;
  assign n4671 = n4657 & ~n4670 ;
  assign n4672 = ~n284 & ~n492 ;
  assign n4673 = n524 & n1002 ;
  assign n4674 = n159 & n4673 ;
  assign n4675 = n2653 & n4145 ;
  assign n4676 = n568 & n1113 ;
  assign n4677 = n4368 & n4676 ;
  assign n4678 = ~n4675 & ~n4677 ;
  assign n4679 = ~n4674 & n4678 ;
  assign n4680 = ~n4672 & ~n4679 ;
  assign n4681 = ~n4671 & ~n4680 ;
  assign n4682 = n4656 & ~n4681 ;
  assign n4683 = n1201 & n4158 ;
  assign n4684 = ~x11 & n1169 ;
  assign n4685 = ~n28 & ~n197 ;
  assign n4686 = ~n1038 & ~n4685 ;
  assign n4687 = ~n4684 & ~n4686 ;
  assign n4688 = n4359 & ~n4687 ;
  assign n4689 = ~n4683 & ~n4688 ;
  assign n4690 = n2631 & ~n4689 ;
  assign n4691 = n474 & n2480 ;
  assign n4692 = n1958 & n4691 ;
  assign n4693 = ~n4690 & ~n4692 ;
  assign n4694 = ~n4682 & n4693 ;
  assign n4695 = ~n4655 & n4694 ;
  assign n4696 = n4644 & ~n4695 ;
  assign n4697 = ~x10 & n311 ;
  assign n4698 = x0 & n4697 ;
  assign n4699 = ~n780 & ~n2631 ;
  assign n4700 = ~n4698 & n4699 ;
  assign n4701 = n720 & n2637 ;
  assign n4702 = n55 & n248 ;
  assign n4703 = n4701 & n4702 ;
  assign n4704 = ~n4700 & n4703 ;
  assign n4730 = ~x11 & n311 ;
  assign n4731 = n1327 & n4730 ;
  assign n4732 = ~n2117 & ~n4731 ;
  assign n4733 = x9 & ~n4732 ;
  assign n4734 = ~n830 & ~n4733 ;
  assign n4735 = ~x3 & n568 ;
  assign n4736 = n2653 & n4735 ;
  assign n4737 = ~n4734 & n4736 ;
  assign n4738 = x11 & ~n673 ;
  assign n4739 = n4495 & n4738 ;
  assign n4740 = n4415 & n4497 ;
  assign n4741 = ~n4739 & ~n4740 ;
  assign n4742 = n3914 & ~n4741 ;
  assign n4743 = n1226 & n2480 ;
  assign n4744 = ~n1136 & n2343 ;
  assign n4745 = n4743 & n4744 ;
  assign n4746 = ~n4742 & ~n4745 ;
  assign n4747 = n1226 ^ n605 ;
  assign n4748 = ~x9 & n4747 ;
  assign n4749 = n4748 ^ n605 ;
  assign n4750 = n700 & n4749 ;
  assign n4751 = ~x1 & n1263 ;
  assign n4752 = n105 & n4751 ;
  assign n4753 = ~n4750 & ~n4752 ;
  assign n4754 = n381 & n4344 ;
  assign n4755 = ~n4753 & n4754 ;
  assign n4756 = n4746 & ~n4755 ;
  assign n4757 = ~n4737 & n4756 ;
  assign n4705 = n3718 & n4415 ;
  assign n4706 = n363 & n1459 ;
  assign n4707 = ~n4705 & ~n4706 ;
  assign n4708 = n787 & ~n4707 ;
  assign n4709 = x15 & n4708 ;
  assign n4710 = ~x7 & n104 ;
  assign n4711 = n2343 & n4710 ;
  assign n4712 = ~n888 & ~n1905 ;
  assign n4713 = n4495 & ~n4712 ;
  assign n4714 = ~n4711 & ~n4713 ;
  assign n4715 = n978 & ~n4714 ;
  assign n4716 = ~x3 & n4392 ;
  assign n4717 = x14 & n899 ;
  assign n4718 = ~n1105 & ~n4717 ;
  assign n4719 = n4718 ^ n306 ;
  assign n4720 = n4719 ^ n4718 ;
  assign n4721 = n4718 ^ n4712 ;
  assign n4722 = n4721 ^ n4718 ;
  assign n4723 = n4720 & ~n4722 ;
  assign n4724 = n4723 ^ n4718 ;
  assign n4725 = ~x9 & ~n4724 ;
  assign n4726 = n4725 ^ n4718 ;
  assign n4727 = n4716 & ~n4726 ;
  assign n4728 = ~n4715 & ~n4727 ;
  assign n4729 = ~n4709 & n4728 ;
  assign n4758 = n4757 ^ n4729 ;
  assign n4759 = n4758 ^ n4757 ;
  assign n4760 = n4757 ^ x12 ;
  assign n4761 = n4760 ^ n4757 ;
  assign n4762 = ~n4759 & n4761 ;
  assign n4763 = n4762 ^ n4757 ;
  assign n4764 = ~x8 & ~n4763 ;
  assign n4765 = n4764 ^ n4757 ;
  assign n4766 = ~n4704 & n4765 ;
  assign n4767 = ~n4696 & n4766 ;
  assign n4768 = ~n4643 & n4767 ;
  assign n4769 = x8 & n946 ;
  assign n4770 = n329 & n1025 ;
  assign n4771 = ~n530 & n4411 ;
  assign n4772 = ~n4770 & ~n4771 ;
  assign n4773 = n4769 & ~n4772 ;
  assign n4774 = ~x13 & n198 ;
  assign n4775 = ~x9 & ~n778 ;
  assign n4776 = ~n4774 & n4775 ;
  assign n4777 = ~n1123 & ~n4776 ;
  assign n4778 = n4411 & ~n4777 ;
  assign n4779 = ~n430 & ~n4775 ;
  assign n4780 = ~n503 & n4392 ;
  assign n4781 = ~n4779 & n4780 ;
  assign n4782 = n180 & n2678 ;
  assign n4783 = n282 & n4782 ;
  assign n4784 = ~x11 & n4783 ;
  assign n4785 = ~n4781 & ~n4784 ;
  assign n4786 = ~n4778 & n4785 ;
  assign n4787 = x10 & ~n4786 ;
  assign n4788 = ~n4773 & ~n4787 ;
  assign n4789 = n1682 & ~n4788 ;
  assign n4793 = ~x5 & n3263 ;
  assign n4794 = ~x8 & n1263 ;
  assign n4795 = ~n3009 & ~n4794 ;
  assign n4796 = n4793 & ~n4795 ;
  assign n4797 = ~x12 & n530 ;
  assign n4798 = n4628 & n4797 ;
  assign n4799 = ~n4796 & ~n4798 ;
  assign n4800 = n471 & ~n4799 ;
  assign n4801 = n3462 & n4701 ;
  assign n4802 = ~n4800 & ~n4801 ;
  assign n4790 = ~x9 & n2841 ;
  assign n4791 = ~n4530 & ~n4790 ;
  assign n4792 = n463 & ~n4791 ;
  assign n4803 = n4802 ^ n4792 ;
  assign n4804 = n4803 ^ n4802 ;
  assign n4805 = n4802 ^ n364 ;
  assign n4806 = n4805 ^ n4802 ;
  assign n4807 = n4804 & n4806 ;
  assign n4808 = n4807 ^ n4802 ;
  assign n4809 = ~x0 & ~n4808 ;
  assign n4810 = n4809 ^ n4802 ;
  assign n4811 = ~n4789 & n4810 ;
  assign n4812 = ~x14 & ~n4811 ;
  assign n4813 = n828 & n845 ;
  assign n4814 = n3257 & n4813 ;
  assign n4815 = ~n787 & ~n1683 ;
  assign n4816 = n2735 & ~n4815 ;
  assign n4817 = ~n2952 & ~n4816 ;
  assign n4818 = n112 & ~n4817 ;
  assign n4819 = n2949 ^ n2119 ;
  assign n4820 = ~x8 & n4819 ;
  assign n4821 = n4820 ^ n2119 ;
  assign n4822 = n928 & ~n4821 ;
  assign n4823 = ~n4818 & ~n4822 ;
  assign n4824 = ~x9 & ~n4823 ;
  assign n4825 = ~n4814 & ~n4824 ;
  assign n4826 = n3092 & ~n4825 ;
  assign n4827 = ~n4812 & ~n4826 ;
  assign n4828 = n55 & ~n4827 ;
  assign n4829 = ~x1 & ~x14 ;
  assign n4830 = x10 ^ x2 ;
  assign n4831 = n1327 & n1440 ;
  assign n4832 = ~n828 & ~n1214 ;
  assign n4833 = n283 & ~n4832 ;
  assign n4834 = ~n4831 & ~n4833 ;
  assign n4835 = n4834 ^ x10 ;
  assign n4836 = n4835 ^ n4834 ;
  assign n4837 = n4836 ^ n4830 ;
  assign n4838 = n4795 ^ x3 ;
  assign n4839 = ~n4795 & ~n4838 ;
  assign n4840 = n4839 ^ n4834 ;
  assign n4841 = n4840 ^ n4795 ;
  assign n4842 = n4837 & n4841 ;
  assign n4843 = n4842 ^ n4839 ;
  assign n4844 = n4843 ^ n4795 ;
  assign n4845 = n4830 & ~n4844 ;
  assign n4846 = x11 & n4845 ;
  assign n4847 = ~n1667 & ~n2824 ;
  assign n4848 = ~n284 & n471 ;
  assign n4849 = ~n850 & n4848 ;
  assign n4850 = ~n4847 & n4849 ;
  assign n4851 = ~x10 & n2803 ;
  assign n4852 = ~n405 & ~n4851 ;
  assign n4853 = n112 & n4797 ;
  assign n4854 = ~n4852 & n4853 ;
  assign n4855 = ~n4850 & ~n4854 ;
  assign n4856 = ~n4846 & n4855 ;
  assign n4857 = n4073 & ~n4856 ;
  assign n4858 = ~n555 & n2036 ;
  assign n4859 = x3 & ~n1563 ;
  assign n4860 = ~n850 & n4859 ;
  assign n4861 = n4858 & n4860 ;
  assign n4862 = n318 & n2540 ;
  assign n4863 = n248 & n264 ;
  assign n4864 = ~n4862 & ~n4863 ;
  assign n4865 = n4864 ^ x12 ;
  assign n4866 = n4865 ^ n4864 ;
  assign n4867 = n4866 ^ n4861 ;
  assign n4868 = n392 & n1515 ;
  assign n4869 = n4868 ^ x2 ;
  assign n4870 = x2 & n4869 ;
  assign n4871 = n4870 ^ n4864 ;
  assign n4872 = n4871 ^ x2 ;
  assign n4873 = n4867 & ~n4872 ;
  assign n4874 = n4873 ^ n4870 ;
  assign n4875 = n4874 ^ x2 ;
  assign n4876 = ~n4861 & n4875 ;
  assign n4877 = n4876 ^ n4861 ;
  assign n4878 = n866 & n4877 ;
  assign n4879 = n392 & n1708 ;
  assign n4880 = ~x2 & ~x12 ;
  assign n4881 = ~n650 & ~n2326 ;
  assign n4882 = n4880 & ~n4881 ;
  assign n4883 = n217 & n1739 ;
  assign n4884 = ~n4882 & ~n4883 ;
  assign n4885 = ~n4879 & n4884 ;
  assign n4886 = n1217 & ~n4885 ;
  assign n4887 = n1226 & n1514 ;
  assign n4888 = ~x3 & n1739 ;
  assign n4889 = ~n4887 & ~n4888 ;
  assign n4890 = n175 & ~n4889 ;
  assign n4891 = ~n1708 & ~n1739 ;
  assign n4892 = n798 & ~n4891 ;
  assign n4893 = ~n105 & n4892 ;
  assign n4894 = ~n4890 & ~n4893 ;
  assign n4895 = ~n4886 & n4894 ;
  assign n4896 = n104 & ~n4895 ;
  assign n4897 = n248 & n4330 ;
  assign n4898 = x8 & n226 ;
  assign n4899 = n1327 & n4898 ;
  assign n4900 = ~n4897 & ~n4899 ;
  assign n4901 = n68 & ~n4900 ;
  assign n4902 = n240 & ~n850 ;
  assign n4903 = ~x2 & n1265 ;
  assign n4904 = ~n4902 & ~n4903 ;
  assign n4905 = n1667 & ~n4904 ;
  assign n4906 = ~n4901 & ~n4905 ;
  assign n4907 = n18 & ~n4906 ;
  assign n4908 = ~x10 & ~n1667 ;
  assign n4909 = ~n105 & ~n1246 ;
  assign n4910 = n848 & ~n4909 ;
  assign n4911 = n4908 & n4910 ;
  assign n4912 = ~n650 & n4911 ;
  assign n4913 = ~n4907 & ~n4912 ;
  assign n4914 = ~n4896 & n4913 ;
  assign n4915 = ~n4878 & n4914 ;
  assign n4916 = n2653 & ~n4915 ;
  assign n4917 = ~n4857 & ~n4916 ;
  assign n4918 = n4829 & ~n4917 ;
  assign n4919 = n588 & n2957 ;
  assign n4920 = n3640 & n4887 ;
  assign n4921 = ~n4919 & ~n4920 ;
  assign n4922 = n2822 & n4422 ;
  assign n4923 = ~n4003 & ~n4922 ;
  assign n4924 = ~n4921 & ~n4923 ;
  assign n4925 = n718 & n2822 ;
  assign n4926 = n845 & n4925 ;
  assign n4927 = n1977 & n4368 ;
  assign n4928 = n3021 & n4411 ;
  assign n4929 = ~n4927 & ~n4928 ;
  assign n4930 = n866 & ~n4929 ;
  assign n4931 = n86 & n3286 ;
  assign n4932 = n2653 & n3212 ;
  assign n4933 = ~n4931 & ~n4932 ;
  assign n4934 = n248 & ~n4933 ;
  assign n4935 = ~n4930 & ~n4934 ;
  assign n4936 = ~n4926 & n4935 ;
  assign n4937 = n4936 ^ x1 ;
  assign n4938 = n4937 ^ n4936 ;
  assign n4939 = n489 & n2653 ;
  assign n4940 = n2165 & n4939 ;
  assign n4941 = n1683 & ~n3040 ;
  assign n4942 = x11 & n489 ;
  assign n4943 = n3021 & n4942 ;
  assign n4944 = ~n4941 & ~n4943 ;
  assign n4945 = n3196 & ~n4944 ;
  assign n4946 = ~n4940 & ~n4945 ;
  assign n4947 = n4946 ^ n4936 ;
  assign n4948 = n4938 & n4947 ;
  assign n4949 = n4948 ^ n4936 ;
  assign n4950 = ~n1517 & ~n4949 ;
  assign n4951 = n240 & n3196 ;
  assign n4952 = x14 & n1117 ;
  assign n4953 = n310 & n4952 ;
  assign n4954 = n66 & n262 ;
  assign n4958 = n4954 ^ n3010 ;
  assign n4959 = n4958 ^ n4954 ;
  assign n4955 = ~x8 & ~x14 ;
  assign n4956 = n4955 ^ n4954 ;
  assign n4957 = n4956 ^ n4954 ;
  assign n4960 = n4959 ^ n4957 ;
  assign n4961 = n4954 ^ n1874 ;
  assign n4962 = n4961 ^ n4954 ;
  assign n4963 = n4962 ^ n4959 ;
  assign n4964 = ~n4959 & ~n4963 ;
  assign n4965 = n4964 ^ n4959 ;
  assign n4966 = n4960 & ~n4965 ;
  assign n4967 = n4966 ^ n4964 ;
  assign n4968 = n4967 ^ n4954 ;
  assign n4969 = n4968 ^ n4959 ;
  assign n4970 = ~n786 & ~n4969 ;
  assign n4971 = n4970 ^ n4954 ;
  assign n4972 = ~n4953 & ~n4971 ;
  assign n4973 = n4951 & ~n4972 ;
  assign n4974 = n348 & n2653 ;
  assign n4975 = ~x14 & ~n406 ;
  assign n4976 = n4974 & n4975 ;
  assign n4977 = ~n642 & n4976 ;
  assign n4978 = n442 & n3196 ;
  assign n4979 = ~x11 & n200 ;
  assign n4980 = n4978 & n4979 ;
  assign n4981 = ~n4977 & ~n4980 ;
  assign n4982 = n929 & ~n4981 ;
  assign n4983 = ~n4973 & ~n4982 ;
  assign n4984 = n4983 ^ x9 ;
  assign n4985 = n4984 ^ n4983 ;
  assign n4986 = n4985 ^ n1658 ;
  assign n4987 = ~x7 & n180 ;
  assign n4988 = n334 & n4987 ;
  assign n4989 = n3256 & n3711 ;
  assign n4990 = ~n4988 & ~n4989 ;
  assign n4991 = n1990 & ~n4990 ;
  assign n4992 = ~x3 & n306 ;
  assign n4993 = n3308 & n4992 ;
  assign n4994 = ~x8 & n4993 ;
  assign n4995 = ~n4991 & ~n4994 ;
  assign n4996 = ~n850 & n3308 ;
  assign n4997 = n47 & n2601 ;
  assign n4998 = ~n4996 & ~n4997 ;
  assign n4999 = n38 & ~n4998 ;
  assign n5000 = n4999 ^ n4995 ;
  assign n5001 = n4995 & ~n5000 ;
  assign n5002 = n5001 ^ n4983 ;
  assign n5003 = n5002 ^ n4995 ;
  assign n5004 = ~n4986 & n5003 ;
  assign n5005 = n5004 ^ n5001 ;
  assign n5006 = n5005 ^ n4995 ;
  assign n5007 = ~n1658 & n5006 ;
  assign n5008 = n5007 ^ n1658 ;
  assign n5009 = ~n4950 & n5008 ;
  assign n5010 = ~n4924 & n5009 ;
  assign n5011 = ~n4918 & n5010 ;
  assign n5012 = n344 & n3091 ;
  assign n5013 = ~x9 & n1117 ;
  assign n5014 = n58 & n2946 ;
  assign n5015 = n20 & ~n2119 ;
  assign n5016 = n928 & ~n2949 ;
  assign n5017 = ~n5015 & ~n5016 ;
  assign n5018 = ~n5014 & n5017 ;
  assign n5019 = n5013 & ~n5018 ;
  assign n5020 = n224 & n557 ;
  assign n5021 = ~n198 & n1364 ;
  assign n5022 = ~x11 & n5021 ;
  assign n5023 = n5020 & n5022 ;
  assign n5024 = ~n5019 & ~n5023 ;
  assign n5025 = n265 & n828 ;
  assign n5026 = n318 & n1104 ;
  assign n5027 = n5025 & n5026 ;
  assign n5028 = n1605 & n2735 ;
  assign n5029 = n465 & n828 ;
  assign n5030 = n346 & n5029 ;
  assign n5031 = n1201 & ~n3704 ;
  assign n5032 = ~n5030 & ~n5031 ;
  assign n5033 = ~n5028 & n5032 ;
  assign n5034 = n3686 & ~n5033 ;
  assign n5035 = ~n5027 & ~n5034 ;
  assign n5040 = n818 & n828 ;
  assign n5041 = ~n555 & n874 ;
  assign n5042 = x10 & ~n1703 ;
  assign n5043 = n5041 & ~n5042 ;
  assign n5044 = ~x0 & n2036 ;
  assign n5045 = n555 & n5044 ;
  assign n5046 = ~n354 & n5045 ;
  assign n5047 = ~n5043 & ~n5046 ;
  assign n5048 = ~n5040 & n5047 ;
  assign n5036 = n554 & n2700 ;
  assign n5037 = n866 & ~n2662 ;
  assign n5038 = ~n643 & n5037 ;
  assign n5039 = ~n5036 & ~n5038 ;
  assign n5049 = n5048 ^ n5039 ;
  assign n5050 = n5049 ^ n5048 ;
  assign n5051 = n5048 ^ x12 ;
  assign n5052 = n5051 ^ n5048 ;
  assign n5053 = ~n5050 & ~n5052 ;
  assign n5054 = n5053 ^ n5048 ;
  assign n5055 = x8 & ~n5054 ;
  assign n5056 = n5055 ^ n5048 ;
  assign n5057 = n262 & ~n5056 ;
  assign n5058 = n5035 & ~n5057 ;
  assign n5059 = n5024 & n5058 ;
  assign n5060 = n5012 & ~n5059 ;
  assign n5061 = n364 & n3283 ;
  assign n5062 = ~x11 & n2036 ;
  assign n5063 = n784 & n5062 ;
  assign n5064 = ~n5061 & ~n5063 ;
  assign n5065 = n656 & ~n5064 ;
  assign n5066 = ~n850 & ~n4275 ;
  assign n5067 = ~n525 & ~n4033 ;
  assign n5068 = n778 & ~n5067 ;
  assign n5069 = ~n5066 & ~n5068 ;
  assign n5070 = n2508 & ~n5069 ;
  assign n5071 = ~n5065 & ~n5070 ;
  assign n5072 = n4069 & ~n5071 ;
  assign n5073 = ~n1807 & ~n3146 ;
  assign n5074 = n176 & ~n5073 ;
  assign n5075 = n885 & n1247 ;
  assign n5076 = ~n5074 & ~n5075 ;
  assign n5077 = n2653 & ~n5076 ;
  assign n5078 = n1095 & n3196 ;
  assign n5079 = n2761 & n5078 ;
  assign n5080 = ~n5077 & ~n5079 ;
  assign n5081 = n3710 & ~n5080 ;
  assign n5082 = ~n5072 & ~n5081 ;
  assign n5083 = n2290 & n3721 ;
  assign n5084 = ~n947 & n3307 ;
  assign n5085 = n2675 & n5084 ;
  assign n5086 = ~n5083 & ~n5085 ;
  assign n5087 = n151 & ~n5086 ;
  assign n5088 = n673 & n757 ;
  assign n5089 = n1233 & n5088 ;
  assign n5090 = n4411 & n5089 ;
  assign n5091 = n2625 & n4987 ;
  assign n5092 = n104 & n3196 ;
  assign n5093 = ~x11 & n2675 ;
  assign n5094 = ~n5092 & ~n5093 ;
  assign n5095 = n1214 & n1524 ;
  assign n5096 = ~n1739 & ~n5095 ;
  assign n5097 = ~n5094 & ~n5096 ;
  assign n5098 = ~n5091 & ~n5097 ;
  assign n5099 = n3256 & ~n5098 ;
  assign n5100 = ~n5090 & ~n5099 ;
  assign n5101 = ~n5087 & n5100 ;
  assign n5102 = ~x0 & ~n5101 ;
  assign n5103 = n5082 & ~n5102 ;
  assign n5104 = n348 & ~n5103 ;
  assign n5105 = ~n5060 & ~n5104 ;
  assign n5106 = n5011 & n5105 ;
  assign n5107 = ~n4828 & n5106 ;
  assign n5108 = ~x15 & ~n5107 ;
  assign n5109 = n4768 & ~n5108 ;
  assign n5110 = ~n4493 & n5109 ;
  assign n5111 = ~n371 & ~n1214 ;
  assign n5112 = ~n1173 & ~n5111 ;
  assign n5113 = n4279 & ~n5112 ;
  assign n5114 = ~n4268 & n5113 ;
  assign n5115 = n348 & ~n5114 ;
  assign n5116 = x14 & n2827 ;
  assign n5117 = ~n3418 & ~n5116 ;
  assign n5118 = n5117 ^ n306 ;
  assign n5119 = n5117 ^ n874 ;
  assign n5120 = n5119 ^ n874 ;
  assign n5121 = ~x11 & n4287 ;
  assign n5122 = n5121 ^ n874 ;
  assign n5123 = n5120 & ~n5122 ;
  assign n5124 = n5123 ^ n874 ;
  assign n5125 = ~n5118 & n5124 ;
  assign n5126 = n5125 ^ n306 ;
  assign n5127 = ~n4263 & ~n5126 ;
  assign n5128 = ~x3 & ~n5127 ;
  assign n5129 = ~x12 & n145 ;
  assign n5130 = n4222 & n5129 ;
  assign n5131 = n5117 & ~n5130 ;
  assign n5132 = n3697 & ~n5131 ;
  assign n5133 = ~x0 & n2290 ;
  assign n5134 = ~n248 & ~n5133 ;
  assign n5135 = n38 & n4697 ;
  assign n5136 = ~n5134 & n5135 ;
  assign n5137 = ~n5132 & ~n5136 ;
  assign n5138 = ~n5128 & n5137 ;
  assign n5139 = ~n5115 & n5138 ;
  assign n5140 = n4701 & ~n5139 ;
  assign n5141 = ~n162 & ~n1440 ;
  assign n5142 = n1227 & n1743 ;
  assign n5143 = n306 & n828 ;
  assign n5144 = ~n3960 & n5143 ;
  assign n5145 = ~n5142 & ~n5144 ;
  assign n5146 = n845 & ~n5145 ;
  assign n5147 = n491 & n3225 ;
  assign n5148 = ~n5146 & ~n5147 ;
  assign n5149 = n2654 & ~n5148 ;
  assign n5150 = n395 & n866 ;
  assign n5151 = n828 & n4358 ;
  assign n5152 = n5150 & n5151 ;
  assign n5153 = n817 & n4286 ;
  assign n5154 = n642 & n4561 ;
  assign n5155 = n5153 & n5154 ;
  assign n5156 = ~n5152 & ~n5155 ;
  assign n5157 = ~n5149 & n5156 ;
  assign n5158 = n5141 & ~n5157 ;
  assign n5159 = n858 & n1108 ;
  assign n5160 = n489 & n2213 ;
  assign n5161 = ~n5159 & ~n5160 ;
  assign n5162 = n38 & ~n5161 ;
  assign n5163 = x0 & n4333 ;
  assign n5164 = n263 & n845 ;
  assign n5165 = n5163 & n5164 ;
  assign n5166 = n517 & n1906 ;
  assign n5167 = n900 & n5166 ;
  assign n5168 = ~n5165 & ~n5167 ;
  assign n5169 = ~n5162 & n5168 ;
  assign n5170 = n1630 & ~n5169 ;
  assign n5171 = ~n5158 & ~n5170 ;
  assign n5172 = ~x10 & n1226 ;
  assign n5173 = n817 & n5172 ;
  assign n5174 = x8 & n5173 ;
  assign n5175 = ~x8 & n2154 ;
  assign n5176 = n200 & n1364 ;
  assign n5177 = ~n5175 & ~n5176 ;
  assign n5178 = n762 & ~n5177 ;
  assign n5179 = n1682 & n2213 ;
  assign n5180 = ~x0 & n1515 ;
  assign n5181 = n1246 & n5180 ;
  assign n5182 = ~n5179 & ~n5181 ;
  assign n5183 = ~n5178 & n5182 ;
  assign n5184 = x10 & ~n5183 ;
  assign n5185 = ~n5174 & ~n5184 ;
  assign n5186 = n442 & ~n5185 ;
  assign n5187 = x7 & n5186 ;
  assign n5188 = n282 & n4356 ;
  assign n5189 = x3 & ~x7 ;
  assign n5190 = n3728 & n5189 ;
  assign n5191 = ~n4657 & ~n5190 ;
  assign n5192 = ~x1 & ~n5191 ;
  assign n5193 = ~x9 & n348 ;
  assign n5194 = n3196 & n5193 ;
  assign n5195 = ~n5192 & ~n5194 ;
  assign n5196 = ~n4170 & ~n5195 ;
  assign n5197 = n2991 & n4065 ;
  assign n5198 = ~n5196 & ~n5197 ;
  assign n5199 = n456 & ~n5198 ;
  assign n5200 = n3256 & n4333 ;
  assign n5201 = n290 & n2822 ;
  assign n5202 = n5200 & n5201 ;
  assign n5203 = ~n5199 & ~n5202 ;
  assign n5204 = ~n5188 & n5203 ;
  assign n5205 = n4155 & ~n5204 ;
  assign n5206 = n981 & n1282 ;
  assign n5207 = n329 & n5206 ;
  assign n5208 = ~n3683 & ~n5207 ;
  assign n5209 = n126 & ~n5208 ;
  assign n5210 = n900 & n2653 ;
  assign n5211 = n2312 & n5210 ;
  assign n5212 = ~n5209 & ~n5211 ;
  assign n5213 = n265 & ~n5212 ;
  assign n5214 = n845 & n1270 ;
  assign n5215 = ~x13 & n5214 ;
  assign n5216 = n2527 & n5215 ;
  assign n5217 = n4163 & n5216 ;
  assign n5218 = ~n5213 & ~n5217 ;
  assign n5219 = ~n25 & ~n224 ;
  assign n5220 = ~n5218 & n5219 ;
  assign n5221 = n1328 & n5150 ;
  assign n5222 = n4582 & n5221 ;
  assign n5223 = n997 & n1423 ;
  assign n5224 = n595 & n5223 ;
  assign n5225 = n858 & n2280 ;
  assign n5226 = ~n4770 & ~n5225 ;
  assign n5227 = n3914 & ~n5226 ;
  assign n5228 = x8 & n5227 ;
  assign n5229 = ~n5224 & ~n5228 ;
  assign n5230 = n19 & ~n5229 ;
  assign n5231 = ~n1233 & ~n2527 ;
  assign n5232 = n3903 & ~n5231 ;
  assign n5233 = ~x7 & n624 ;
  assign n5234 = n1954 & n5233 ;
  assign n5235 = n5232 & n5234 ;
  assign n5236 = ~n5230 & ~n5235 ;
  assign n5237 = ~n5222 & n5236 ;
  assign n5238 = x3 & ~x15 ;
  assign n5239 = ~n652 & ~n5238 ;
  assign n5240 = ~n5237 & n5239 ;
  assign n5241 = ~n5220 & ~n5240 ;
  assign n5242 = ~n5205 & n5241 ;
  assign n5243 = ~n5187 & n5242 ;
  assign n5244 = n2478 & n4013 ;
  assign n5245 = n396 & n456 ;
  assign n5246 = ~n1287 & ~n5245 ;
  assign n5247 = n4073 & ~n5246 ;
  assign n5248 = ~n79 & ~n4015 ;
  assign n5249 = n948 & n1855 ;
  assign n5250 = ~n5248 & n5249 ;
  assign n5251 = ~n5247 & ~n5250 ;
  assign n5252 = ~n5244 & n5251 ;
  assign n5253 = x3 & n4286 ;
  assign n5254 = ~n5252 & n5253 ;
  assign n5255 = n265 & n4002 ;
  assign n5256 = ~x14 & n290 ;
  assign n5257 = n4582 & n5256 ;
  assign n5258 = ~n5255 & ~n5257 ;
  assign n5259 = n306 & ~n5258 ;
  assign n5260 = n786 & n4163 ;
  assign n5261 = ~n5259 & ~n5260 ;
  assign n5262 = ~x3 & n1671 ;
  assign n5263 = ~n5261 & n5262 ;
  assign n5264 = n4024 & n4588 ;
  assign n5265 = n442 & n5264 ;
  assign n5266 = ~n5263 & ~n5265 ;
  assign n5267 = ~n5254 & n5266 ;
  assign n5268 = n642 & ~n5267 ;
  assign n5269 = n5243 & ~n5268 ;
  assign n5270 = n5171 & n5269 ;
  assign n5271 = ~n5140 & n5270 ;
  assign n5272 = n2868 & ~n4732 ;
  assign n5273 = n2803 & n4182 ;
  assign n5274 = n45 & n311 ;
  assign n5275 = ~n673 & n1683 ;
  assign n5276 = ~n5274 & ~n5275 ;
  assign n5277 = x11 & n1679 ;
  assign n5278 = ~n5276 & n5277 ;
  assign n5279 = ~n5273 & ~n5278 ;
  assign n5280 = ~n5272 & n5279 ;
  assign n5281 = n858 & ~n5280 ;
  assign n5282 = x1 & n5281 ;
  assign n5283 = n748 & n1263 ;
  assign n5284 = ~x7 & n866 ;
  assign n5285 = n5283 & n5284 ;
  assign n5286 = ~x11 & ~n3729 ;
  assign n5287 = ~x7 & n217 ;
  assign n5288 = ~n5286 & ~n5287 ;
  assign n5289 = n900 & ~n5288 ;
  assign n5290 = n392 & n492 ;
  assign n5291 = x11 & ~n126 ;
  assign n5292 = ~n375 & ~n659 ;
  assign n5293 = ~n5291 & ~n5292 ;
  assign n5294 = ~n870 & n5293 ;
  assign n5295 = ~n5290 & ~n5294 ;
  assign n5296 = n622 & ~n5295 ;
  assign n5297 = ~n5289 & ~n5296 ;
  assign n5298 = n1682 & ~n5297 ;
  assign n5299 = ~x9 & ~n1282 ;
  assign n5300 = ~n503 & n1679 ;
  assign n5301 = ~n5299 & n5300 ;
  assign n5302 = n5301 ^ n1202 ;
  assign n5303 = n5302 ^ x1 ;
  assign n5310 = n5303 ^ n5302 ;
  assign n5304 = n5303 ^ n698 ;
  assign n5305 = n5304 ^ n5302 ;
  assign n5306 = n5303 ^ n5301 ;
  assign n5307 = n5306 ^ n698 ;
  assign n5308 = n5307 ^ n5305 ;
  assign n5309 = n5305 & ~n5308 ;
  assign n5311 = n5310 ^ n5309 ;
  assign n5312 = n5311 ^ n5305 ;
  assign n5313 = n5302 ^ x9 ;
  assign n5314 = n5309 ^ n5305 ;
  assign n5315 = ~n5313 & n5314 ;
  assign n5316 = n5315 ^ n5302 ;
  assign n5317 = ~n5312 & n5316 ;
  assign n5318 = n5317 ^ n5302 ;
  assign n5319 = n5318 ^ n1202 ;
  assign n5320 = n5319 ^ n5302 ;
  assign n5321 = ~n2116 & n5320 ;
  assign n5322 = n284 & n1010 ;
  assign n5323 = ~n1327 & n5322 ;
  assign n5324 = ~x1 & n5323 ;
  assign n5325 = n1169 & n5172 ;
  assign n5326 = ~n5324 & ~n5325 ;
  assign n5327 = n845 & n5193 ;
  assign n5328 = n260 & n1202 ;
  assign n5329 = n2824 & n5328 ;
  assign n5330 = ~n5327 & ~n5329 ;
  assign n5331 = n5326 & n5330 ;
  assign n5332 = n396 & n1336 ;
  assign n5333 = n5332 ^ x1 ;
  assign n5334 = x11 ^ x9 ;
  assign n5335 = n1327 ^ x11 ;
  assign n5336 = n5334 & n5335 ;
  assign n5337 = n5336 ^ x11 ;
  assign n5338 = n5337 ^ n5332 ;
  assign n5339 = n5333 & n5338 ;
  assign n5340 = n5339 ^ n5336 ;
  assign n5341 = n5340 ^ x11 ;
  assign n5342 = n5341 ^ x1 ;
  assign n5343 = ~n5332 & n5342 ;
  assign n5344 = n5343 ^ n5332 ;
  assign n5345 = n5344 ^ n5332 ;
  assign n5346 = n529 & ~n5345 ;
  assign n5347 = n5331 & ~n5346 ;
  assign n5348 = ~n5321 & n5347 ;
  assign n5349 = n884 & ~n5348 ;
  assign n5350 = ~n5298 & ~n5349 ;
  assign n5351 = ~n5285 & n5350 ;
  assign n5352 = n24 & n2803 ;
  assign n5353 = x9 & ~n5352 ;
  assign n5354 = ~n383 & n5353 ;
  assign n5355 = n163 ^ x11 ;
  assign n5356 = n5355 ^ x11 ;
  assign n5357 = n5356 ^ x9 ;
  assign n5358 = n1555 ^ n110 ;
  assign n5359 = ~n110 & ~n5358 ;
  assign n5360 = n5359 ^ x11 ;
  assign n5361 = n5360 ^ n110 ;
  assign n5362 = n5357 & ~n5361 ;
  assign n5363 = n5362 ^ n5359 ;
  assign n5364 = n5363 ^ n110 ;
  assign n5365 = ~x9 & ~n5364 ;
  assign n5366 = n5365 ^ x9 ;
  assign n5367 = ~n5354 & n5366 ;
  assign n5368 = n17 & ~n5367 ;
  assign n5369 = n4027 & n5368 ;
  assign n5370 = ~n428 & n1627 ;
  assign n5371 = ~n4672 & n5370 ;
  assign n5372 = ~x3 & n503 ;
  assign n5373 = ~x15 & ~n375 ;
  assign n5374 = ~n276 & n828 ;
  assign n5375 = ~n5373 & n5374 ;
  assign n5376 = ~n5372 & ~n5375 ;
  assign n5377 = n748 & ~n5376 ;
  assign n5378 = n1627 & n4542 ;
  assign n5379 = ~n587 & ~n5378 ;
  assign n5380 = n375 & ~n5379 ;
  assign n5381 = ~n5377 & ~n5380 ;
  assign n5382 = ~n5371 & n5381 ;
  assign n5383 = n1905 & ~n5382 ;
  assign n5384 = ~x11 & n1349 ;
  assign n5385 = n888 & n5384 ;
  assign n5386 = n462 & n828 ;
  assign n5387 = ~n2398 & ~n5386 ;
  assign n5388 = ~n5385 & n5387 ;
  assign n5389 = n375 & ~n5388 ;
  assign n5390 = x13 & n375 ;
  assign n5391 = ~x11 & n5390 ;
  assign n5392 = ~n1642 & ~n5391 ;
  assign n5393 = n749 & n1282 ;
  assign n5394 = ~n5392 & n5393 ;
  assign n5395 = ~n5389 & ~n5394 ;
  assign n5396 = ~n5383 & n5395 ;
  assign n5397 = n1002 & ~n5396 ;
  assign n5398 = ~n5369 & ~n5397 ;
  assign n5399 = n5351 & n5398 ;
  assign n5400 = n524 ^ x9 ;
  assign n5401 = n5400 ^ n1042 ;
  assign n5402 = n5400 & n5401 ;
  assign n5403 = n5402 ^ x9 ;
  assign n5404 = n5403 ^ n5400 ;
  assign n5410 = ~x12 & n471 ;
  assign n5411 = ~n673 & n5410 ;
  assign n5412 = ~n405 & ~n5411 ;
  assign n5413 = n5412 ^ x3 ;
  assign n5405 = n524 ^ x3 ;
  assign n5406 = n5405 ^ x9 ;
  assign n5407 = n5406 ^ n5400 ;
  assign n5408 = x9 & ~n5407 ;
  assign n5409 = n5408 ^ n5405 ;
  assign n5414 = n5413 ^ n5409 ;
  assign n5415 = n5405 ^ n145 ;
  assign n5416 = n5415 ^ n5413 ;
  assign n5417 = ~n145 & ~n5416 ;
  assign n5418 = n5417 ^ x9 ;
  assign n5419 = n5414 & n5418 ;
  assign n5420 = n5419 ^ n5405 ;
  assign n5421 = n5420 ^ n5400 ;
  assign n5422 = n5421 ^ n1042 ;
  assign n5423 = n5404 & ~n5422 ;
  assign n5424 = n5423 ^ n5408 ;
  assign n5425 = n5424 ^ n5419 ;
  assign n5426 = n5425 ^ x9 ;
  assign n5427 = n5399 & ~n5426 ;
  assign n5428 = n5427 ^ x8 ;
  assign n5429 = n5428 ^ n5427 ;
  assign n5430 = n5429 ^ n5282 ;
  assign n5431 = ~x3 & n1423 ;
  assign n5432 = n105 & n5431 ;
  assign n5433 = n511 & n2358 ;
  assign n5434 = ~n846 & ~n5433 ;
  assign n5435 = x1 & ~n5434 ;
  assign n5436 = n110 ^ x10 ;
  assign n5437 = ~n57 & ~n1667 ;
  assign n5438 = n5437 ^ n110 ;
  assign n5439 = n5438 ^ n5437 ;
  assign n5440 = n5439 ^ n5436 ;
  assign n5441 = n1283 ^ x1 ;
  assign n5442 = ~n1283 & n5441 ;
  assign n5443 = n5442 ^ n5437 ;
  assign n5444 = n5443 ^ n1283 ;
  assign n5445 = n5440 & n5444 ;
  assign n5446 = n5445 ^ n5442 ;
  assign n5447 = n5446 ^ n1283 ;
  assign n5448 = n5436 & ~n5447 ;
  assign n5449 = ~n5435 & ~n5448 ;
  assign n5450 = n260 & ~n5449 ;
  assign n5451 = ~x1 & n5433 ;
  assign n5452 = ~x3 & n2827 ;
  assign n5453 = ~n5451 & ~n5452 ;
  assign n5454 = n623 & ~n5453 ;
  assign n5455 = ~n1214 & ~n1246 ;
  assign n5456 = ~n2329 & n5455 ;
  assign n5457 = n405 & ~n5456 ;
  assign n5458 = ~n5454 & ~n5457 ;
  assign n5459 = ~n5450 & n5458 ;
  assign n5460 = ~n5432 & n5459 ;
  assign n5461 = n1002 & ~n5460 ;
  assign n5462 = n1214 & n1679 ;
  assign n5463 = ~x12 & n473 ;
  assign n5464 = ~n1656 & ~n5463 ;
  assign n5465 = n328 & ~n5464 ;
  assign n5466 = ~n5462 & ~n5465 ;
  assign n5467 = x7 & n109 ;
  assign n5468 = ~n5466 & n5467 ;
  assign n5469 = n718 & n1665 ;
  assign n5470 = n1050 & n5469 ;
  assign n5471 = n2512 & ~n2803 ;
  assign n5472 = ~n197 & n5471 ;
  assign n5473 = ~n5470 & ~n5472 ;
  assign n5474 = n371 & ~n5473 ;
  assign n5475 = ~n5468 & ~n5474 ;
  assign n5478 = ~x12 & ~n392 ;
  assign n5479 = n348 & ~n5478 ;
  assign n5480 = ~n328 & ~n1667 ;
  assign n5481 = n1950 & ~n5480 ;
  assign n5482 = n869 & n4035 ;
  assign n5483 = ~n56 & n5482 ;
  assign n5484 = ~n5481 & ~n5483 ;
  assign n5485 = ~n5479 & n5484 ;
  assign n5476 = ~x3 & n749 ;
  assign n5477 = ~n5384 & ~n5476 ;
  assign n5486 = n5485 ^ n5477 ;
  assign n5487 = n5485 ^ x10 ;
  assign n5488 = n5487 ^ n5485 ;
  assign n5489 = n5488 ^ n884 ;
  assign n5490 = ~n5486 & n5489 ;
  assign n5491 = n5490 ^ n5477 ;
  assign n5492 = n884 & n5491 ;
  assign n5493 = n5475 & ~n5492 ;
  assign n5494 = ~n5461 & n5493 ;
  assign n5495 = n5494 ^ x9 ;
  assign n5496 = ~n5494 & n5495 ;
  assign n5497 = n5496 ^ n5427 ;
  assign n5498 = n5497 ^ n5494 ;
  assign n5499 = n5430 & n5498 ;
  assign n5500 = n5499 ^ n5496 ;
  assign n5501 = n5500 ^ n5494 ;
  assign n5502 = ~n5282 & ~n5501 ;
  assign n5503 = n5502 ^ n5282 ;
  assign n5504 = n5503 ^ x5 ;
  assign n5505 = n5504 ^ n5503 ;
  assign n5506 = n5505 ^ n5271 ;
  assign n5507 = ~x3 & n66 ;
  assign n5508 = n2625 & n5507 ;
  assign n5509 = n2605 & n4333 ;
  assign n5510 = n60 & ~n1795 ;
  assign n5511 = ~n846 & n5510 ;
  assign n5512 = ~x3 & n19 ;
  assign n5513 = n348 & n1227 ;
  assign n5514 = ~n5512 & ~n5513 ;
  assign n5515 = n1682 & ~n5514 ;
  assign n5516 = ~n145 & ~n718 ;
  assign n5517 = n5507 & ~n5516 ;
  assign n5518 = ~n5515 & ~n5517 ;
  assign n5519 = ~n5511 & n5518 ;
  assign n5520 = n346 & ~n5519 ;
  assign n5521 = ~n2116 & ~n2466 ;
  assign n5522 = n4168 & n5521 ;
  assign n5523 = ~n5520 & ~n5522 ;
  assign n5524 = ~n5509 & n5523 ;
  assign n5525 = ~n467 & ~n5524 ;
  assign n5526 = ~x10 & n462 ;
  assign n5527 = n4672 & n5526 ;
  assign n5528 = x8 & n5527 ;
  assign n5529 = ~n373 & n5528 ;
  assign n5530 = n25 & n1515 ;
  assign n5531 = n109 & n5530 ;
  assign n5532 = n558 & ~n2541 ;
  assign n5533 = ~n5531 & ~n5532 ;
  assign n5534 = ~n5529 & n5533 ;
  assign n5535 = n4005 & ~n5534 ;
  assign n5536 = ~n5525 & ~n5535 ;
  assign n5537 = ~n633 & ~n1949 ;
  assign n5538 = n405 & ~n5537 ;
  assign n5539 = n404 & n2395 ;
  assign n5540 = ~n5538 & ~n5539 ;
  assign n5541 = n1682 & ~n5540 ;
  assign n5542 = ~n871 & n1682 ;
  assign n5543 = n866 & ~n1704 ;
  assign n5544 = ~n2036 & n5543 ;
  assign n5545 = ~n5542 & ~n5544 ;
  assign n5546 = n328 & ~n5545 ;
  assign n5547 = ~n1263 & n4410 ;
  assign n5548 = ~n1423 & n5547 ;
  assign n5549 = ~n1038 & n5548 ;
  assign n5550 = n473 & ~n4672 ;
  assign n5551 = ~n1642 & ~n5550 ;
  assign n5552 = n4023 & ~n5551 ;
  assign n5553 = n473 & n1683 ;
  assign n5554 = n276 & n5553 ;
  assign n5555 = ~n5552 & ~n5554 ;
  assign n5556 = ~n5549 & n5555 ;
  assign n5557 = ~n5546 & n5556 ;
  assign n5558 = x11 & ~n5557 ;
  assign n5559 = ~n5541 & ~n5558 ;
  assign n5560 = n206 & ~n5559 ;
  assign n5561 = n5560 ^ n5536 ;
  assign n5562 = n1946 & n2471 ;
  assign n5563 = n56 & ~n370 ;
  assign n5564 = n1104 & ~n5563 ;
  assign n5565 = ~n284 & n900 ;
  assign n5566 = x1 & ~n529 ;
  assign n5567 = ~n375 & n5566 ;
  assign n5568 = ~n5565 & ~n5567 ;
  assign n5569 = n122 & ~n5568 ;
  assign n5570 = ~n5564 & ~n5569 ;
  assign n5571 = ~x13 & ~n5570 ;
  assign n5572 = ~n512 & ~n1169 ;
  assign n5573 = ~x0 & n2326 ;
  assign n5574 = ~n453 & n5573 ;
  assign n5575 = ~n5572 & n5574 ;
  assign n5576 = ~n5571 & ~n5575 ;
  assign n5577 = ~n5562 & n5576 ;
  assign n5578 = n1282 & ~n5577 ;
  assign n5579 = ~n4147 & n5390 ;
  assign n5580 = ~x12 & n5579 ;
  assign n5581 = ~n1555 & n1682 ;
  assign n5582 = ~n2477 & n5581 ;
  assign n5583 = n38 & n5582 ;
  assign n5584 = ~n55 & ~n395 ;
  assign n5585 = x3 & ~n517 ;
  assign n5586 = n5584 & ~n5585 ;
  assign n5587 = ~n405 & ~n5586 ;
  assign n5588 = n5587 ^ x0 ;
  assign n5589 = n5588 ^ n5587 ;
  assign n5590 = x12 & n348 ;
  assign n5591 = ~n104 & ~n1131 ;
  assign n5592 = n5590 & ~n5591 ;
  assign n5593 = ~n404 & n462 ;
  assign n5594 = ~x3 & ~n2607 ;
  assign n5595 = n5593 & n5594 ;
  assign n5596 = ~n1031 & n5595 ;
  assign n5597 = ~n5592 & ~n5596 ;
  assign n5598 = n529 & n1382 ;
  assign n5599 = x11 & n5598 ;
  assign n5600 = n5597 & ~n5599 ;
  assign n5601 = n5600 ^ n5587 ;
  assign n5602 = ~n5589 & n5601 ;
  assign n5603 = n5602 ^ n5587 ;
  assign n5604 = ~n5583 & n5603 ;
  assign n5605 = ~n5580 & n5604 ;
  assign n5606 = ~n5578 & n5605 ;
  assign n5607 = n5606 ^ x8 ;
  assign n5608 = n5607 ^ n5606 ;
  assign n5609 = ~n656 & n978 ;
  assign n5610 = n1031 & n5609 ;
  assign n5611 = n1667 & n5610 ;
  assign n5612 = ~n890 & n1683 ;
  assign n5613 = ~n2037 & ~n5612 ;
  assign n5614 = n554 & ~n5613 ;
  assign n5615 = ~x13 & n1364 ;
  assign n5616 = n489 & n5615 ;
  assign n5617 = ~n5614 & ~n5616 ;
  assign n5618 = n652 & ~n5617 ;
  assign n5619 = ~x13 & n1683 ;
  assign n5620 = n104 & n5619 ;
  assign n5621 = n1247 & n2747 ;
  assign n5622 = ~n5040 & ~n5621 ;
  assign n5623 = ~n5620 & n5622 ;
  assign n5624 = n328 & ~n5623 ;
  assign n5625 = n25 & n524 ;
  assign n5626 = n656 & n1214 ;
  assign n5627 = n5625 & n5626 ;
  assign n5628 = n224 & n1030 ;
  assign n5629 = n2291 & n5628 ;
  assign n5630 = ~n5627 & ~n5629 ;
  assign n5631 = x15 & ~n5630 ;
  assign n5632 = ~n5624 & ~n5631 ;
  assign n5633 = ~x3 & n3869 ;
  assign n5634 = ~n642 & n1682 ;
  assign n5635 = ~n2350 & ~n5634 ;
  assign n5636 = x10 & n284 ;
  assign n5637 = ~n5635 & n5636 ;
  assign n5638 = ~n5633 & ~n5637 ;
  assign n5639 = n1682 & ~n4074 ;
  assign n5640 = ~n5041 & ~n5639 ;
  assign n5641 = n2395 & ~n5640 ;
  assign n5642 = n5638 & ~n5641 ;
  assign n5643 = n5632 & n5642 ;
  assign n5644 = ~n5618 & n5643 ;
  assign n5645 = n5644 ^ x1 ;
  assign n5646 = n5645 ^ n5644 ;
  assign n5647 = n5646 ^ n5611 ;
  assign n5648 = ~n503 & ~n1364 ;
  assign n5649 = n5328 & ~n5648 ;
  assign n5650 = ~n828 & ~n4098 ;
  assign n5651 = n346 & n5650 ;
  assign n5652 = ~n1010 & ~n5651 ;
  assign n5653 = n5652 ^ x3 ;
  assign n5654 = n5653 ^ n5652 ;
  assign n5655 = n5654 ^ n5649 ;
  assign n5656 = n104 & n828 ;
  assign n5657 = ~n1131 & ~n5656 ;
  assign n5658 = n5657 ^ x14 ;
  assign n5659 = ~n5657 & ~n5658 ;
  assign n5660 = n5659 ^ n5652 ;
  assign n5661 = n5660 ^ n5657 ;
  assign n5662 = ~n5655 & n5661 ;
  assign n5663 = n5662 ^ n5659 ;
  assign n5664 = n5663 ^ n5657 ;
  assign n5665 = ~n5649 & ~n5664 ;
  assign n5666 = n5665 ^ n5649 ;
  assign n5667 = n5666 ^ x0 ;
  assign n5668 = x0 & n5667 ;
  assign n5669 = n5668 ^ n5644 ;
  assign n5670 = n5669 ^ x0 ;
  assign n5671 = n5647 & ~n5670 ;
  assign n5672 = n5671 ^ n5668 ;
  assign n5673 = n5672 ^ x0 ;
  assign n5674 = ~n5611 & n5673 ;
  assign n5675 = n5674 ^ n5611 ;
  assign n5676 = n5675 ^ n5606 ;
  assign n5677 = ~n5608 & ~n5676 ;
  assign n5678 = n5677 ^ n5606 ;
  assign n5679 = n5678 ^ n5536 ;
  assign n5680 = ~n5561 & n5679 ;
  assign n5681 = n5680 ^ n5677 ;
  assign n5682 = n5681 ^ n5606 ;
  assign n5683 = n5682 ^ n5560 ;
  assign n5684 = n5536 & ~n5683 ;
  assign n5685 = n5684 ^ n5536 ;
  assign n5686 = ~n5508 & n5685 ;
  assign n5687 = n5686 ^ x7 ;
  assign n5688 = ~n5686 & n5687 ;
  assign n5689 = n5688 ^ n5503 ;
  assign n5690 = n5689 ^ n5686 ;
  assign n5691 = ~n5506 & ~n5690 ;
  assign n5692 = n5691 ^ n5688 ;
  assign n5693 = n5692 ^ n5686 ;
  assign n5694 = n5271 & ~n5693 ;
  assign n5695 = n5694 ^ n5271 ;
  assign n5696 = n5695 ^ x2 ;
  assign n5697 = n5696 ^ n5695 ;
  assign n5698 = ~x13 & x15 ;
  assign n5699 = n3903 & n5698 ;
  assign n5700 = n393 & n1241 ;
  assign n5701 = ~n5699 & ~n5700 ;
  assign n5702 = n4974 & ~n5701 ;
  assign n5703 = ~x11 & ~n56 ;
  assign n5704 = ~x7 & n531 ;
  assign n5705 = ~n2654 & ~n5704 ;
  assign n5706 = n5703 & ~n5705 ;
  assign n5707 = n1435 & n5193 ;
  assign n5708 = n955 & n5707 ;
  assign n5709 = ~n5706 & ~n5708 ;
  assign n5710 = n1423 & ~n5709 ;
  assign n5711 = ~n5702 & ~n5710 ;
  assign n5712 = n60 & ~n5711 ;
  assign n5713 = ~n1062 & ~n3172 ;
  assign n5714 = x15 & n348 ;
  assign n5715 = ~n5713 & n5714 ;
  assign n5716 = n846 & n1124 ;
  assign n5717 = ~n5715 & ~n5716 ;
  assign n5718 = n633 & n4069 ;
  assign n5719 = ~n5717 & n5718 ;
  assign n5720 = ~n5712 & ~n5719 ;
  assign n5721 = ~x9 & n2036 ;
  assign n5722 = n227 & n524 ;
  assign n5723 = n5721 & n5722 ;
  assign n5724 = n4574 & n5723 ;
  assign n5725 = ~x1 & n554 ;
  assign n5726 = n2754 & n5725 ;
  assign n5727 = n4073 & n5726 ;
  assign n5728 = n2478 ^ n900 ;
  assign n5729 = ~x13 & n164 ;
  assign n5730 = n827 & n2116 ;
  assign n5731 = n5729 & n5730 ;
  assign n5732 = n5731 ^ n5728 ;
  assign n5733 = n5732 ^ n2478 ;
  assign n5734 = n5733 ^ n5732 ;
  assign n5735 = n404 & n1226 ;
  assign n5736 = n2822 & n5735 ;
  assign n5737 = n1002 & n1435 ;
  assign n5738 = n1275 & n5737 ;
  assign n5739 = ~n5736 & ~n5738 ;
  assign n5740 = n5739 ^ n5732 ;
  assign n5741 = n5740 ^ n5728 ;
  assign n5742 = n5734 & n5741 ;
  assign n5743 = n5742 ^ n5739 ;
  assign n5744 = x13 & n4349 ;
  assign n5745 = ~n2842 & ~n5744 ;
  assign n5746 = n5739 & n5745 ;
  assign n5747 = n5746 ^ n5728 ;
  assign n5748 = n5743 & ~n5747 ;
  assign n5749 = n5748 ^ n5746 ;
  assign n5750 = ~n5728 & n5749 ;
  assign n5751 = n5750 ^ n5742 ;
  assign n5752 = n5751 ^ n900 ;
  assign n5753 = n5752 ^ n5739 ;
  assign n5754 = ~n5727 & ~n5753 ;
  assign n5755 = ~x3 & ~n5754 ;
  assign n5756 = ~n5724 & ~n5755 ;
  assign n5757 = ~n3960 & ~n5756 ;
  assign n5758 = n2859 & n4521 ;
  assign n5759 = n1214 & n1565 ;
  assign n5760 = n490 & n4974 ;
  assign n5761 = n4356 & ~n4649 ;
  assign n5762 = ~n3682 & ~n4457 ;
  assign n5763 = n25 & n4339 ;
  assign n5764 = ~n5762 & n5763 ;
  assign n5765 = ~n5761 & ~n5764 ;
  assign n5766 = ~n5760 & n5765 ;
  assign n5767 = n5759 & ~n5766 ;
  assign n5768 = ~n5758 & ~n5767 ;
  assign n5769 = ~x8 & ~n5768 ;
  assign n5770 = n345 & n3862 ;
  assign n5771 = n833 & n4974 ;
  assign n5772 = ~n5770 & ~n5771 ;
  assign n5773 = n371 & ~n5772 ;
  assign n5774 = ~n5769 & ~n5773 ;
  assign n5775 = ~n5757 & n5774 ;
  assign n5776 = n5720 & n5775 ;
  assign n5777 = n5776 ^ n5695 ;
  assign n5778 = ~n5697 & n5777 ;
  assign n5779 = n5778 ^ n5695 ;
  assign n5780 = n5110 & n5779 ;
  assign n5781 = ~n4329 & n5780 ;
  assign n5782 = ~n2702 & ~n5781 ;
  assign n5783 = ~n3959 & ~n5782 ;
  assign n5784 = n2453 & n5783 ;
  assign n5785 = x9 & n2633 ;
  assign n5786 = n659 & ~n4955 ;
  assign n5787 = x12 & n5786 ;
  assign n5788 = n5787 ^ x11 ;
  assign n5789 = n5788 ^ n5787 ;
  assign n5790 = n5787 ^ n5469 ;
  assign n5791 = n5790 ^ n5787 ;
  assign n5792 = n5789 & n5791 ;
  assign n5793 = n5792 ^ n5787 ;
  assign n5794 = ~n467 & n5793 ;
  assign n5795 = n5794 ^ n5787 ;
  assign n5796 = n5785 & n5795 ;
  assign n5797 = n1217 & n5636 ;
  assign n5798 = n1226 & n5797 ;
  assign n5799 = n290 & n5463 ;
  assign n5800 = ~n2783 & ~n5799 ;
  assign n5801 = n5800 ^ n145 ;
  assign n5802 = n5801 ^ n5800 ;
  assign n5803 = n5800 ^ n1263 ;
  assign n5804 = n5803 ^ n5800 ;
  assign n5805 = n5802 & n5804 ;
  assign n5806 = n5805 ^ n5800 ;
  assign n5807 = ~x8 & ~n5806 ;
  assign n5808 = n5807 ^ n5800 ;
  assign n5809 = n373 & ~n5808 ;
  assign n5810 = ~x11 & ~n5809 ;
  assign n5811 = n283 & n1601 ;
  assign n5812 = x0 & n5811 ;
  assign n5813 = n275 & n1656 ;
  assign n5814 = ~n1665 & ~n5238 ;
  assign n5815 = n299 & n5814 ;
  assign n5816 = ~n5813 & ~n5815 ;
  assign n5817 = n45 & ~n5816 ;
  assign n5818 = n276 & n3009 ;
  assign n5819 = x15 & n404 ;
  assign n5820 = n1117 & n5819 ;
  assign n5821 = ~n5818 & ~n5820 ;
  assign n5822 = n866 & ~n5821 ;
  assign n5823 = x11 & ~n5822 ;
  assign n5824 = ~n5817 & n5823 ;
  assign n5825 = x14 & ~n5824 ;
  assign n5826 = ~n5797 & ~n5825 ;
  assign n5827 = ~n5812 & n5826 ;
  assign n5828 = ~n5810 & ~n5827 ;
  assign n5829 = ~n467 & n651 ;
  assign n5830 = n1682 & n5829 ;
  assign n5831 = ~n5828 & ~n5830 ;
  assign n5832 = ~n5798 & n5831 ;
  assign n5835 = n5832 ^ x9 ;
  assign n5836 = n5835 ^ n5832 ;
  assign n5833 = n5832 ^ n1906 ;
  assign n5834 = n5833 ^ n5832 ;
  assign n5837 = n5836 ^ n5834 ;
  assign n5838 = n1246 & n1905 ;
  assign n5839 = n5838 ^ n5832 ;
  assign n5840 = n5839 ^ n5832 ;
  assign n5841 = n5840 ^ n5836 ;
  assign n5842 = n5836 & n5841 ;
  assign n5843 = n5842 ^ n5836 ;
  assign n5844 = n5837 & n5843 ;
  assign n5845 = n5844 ^ n5842 ;
  assign n5846 = n5845 ^ n5832 ;
  assign n5847 = n5846 ^ n5836 ;
  assign n5848 = ~x7 & ~n5847 ;
  assign n5849 = n5848 ^ n5832 ;
  assign n5850 = ~n5796 & n5849 ;
  assign n5851 = ~x2 & n79 ;
  assign n5852 = ~n5850 & n5851 ;
  assign n5853 = n28 & n4987 ;
  assign n5854 = n2480 & n5729 ;
  assign n5855 = n57 & n2901 ;
  assign n5856 = ~n5854 & ~n5855 ;
  assign n5857 = x2 & ~n5856 ;
  assign n5858 = ~n669 & ~n3730 ;
  assign n5859 = n57 & ~n5858 ;
  assign n5860 = n370 & n3306 ;
  assign n5861 = ~n5859 & ~n5860 ;
  assign n5862 = ~n5857 & n5861 ;
  assign n5863 = ~n5853 & n5862 ;
  assign n5864 = n2395 & ~n5863 ;
  assign n5865 = ~x10 & n1565 ;
  assign n5866 = n176 & n5865 ;
  assign n5867 = n784 & n1169 ;
  assign n5868 = ~x13 & n5867 ;
  assign n5869 = ~n5866 & ~n5868 ;
  assign n5870 = ~n18 & ~n557 ;
  assign n5871 = n5870 ^ x1 ;
  assign n5872 = n5871 ^ n5870 ;
  assign n5873 = n5872 ^ n44 ;
  assign n5874 = n5870 ^ n889 ;
  assign n5875 = n5873 & ~n5874 ;
  assign n5876 = n5875 ^ n889 ;
  assign n5877 = n44 & n5876 ;
  assign n5878 = n5869 & ~n5877 ;
  assign n5879 = n4359 & ~n5878 ;
  assign n5880 = ~n18 & ~n2558 ;
  assign n5881 = x1 & ~n5880 ;
  assign n5882 = ~n2637 & n5881 ;
  assign n5883 = ~n4254 & ~n5882 ;
  assign n5884 = n180 & ~n5883 ;
  assign n5885 = x14 & n5884 ;
  assign n5886 = n2841 ^ x1 ;
  assign n5887 = n5886 ^ n2841 ;
  assign n5888 = ~x2 & x13 ;
  assign n5889 = n2653 & n5888 ;
  assign n5890 = ~n4616 & ~n5889 ;
  assign n5891 = n5890 ^ n2841 ;
  assign n5892 = ~n5887 & ~n5891 ;
  assign n5893 = n5892 ^ n2841 ;
  assign n5894 = n1030 & n5893 ;
  assign n5895 = ~n5885 & ~n5894 ;
  assign n5896 = ~x3 & ~n5895 ;
  assign n5897 = ~n5879 & ~n5896 ;
  assign n5898 = ~n5864 & n5897 ;
  assign n5899 = ~x12 & ~n5898 ;
  assign n5900 = n526 & n919 ;
  assign n5901 = ~n405 & ~n1671 ;
  assign n5902 = n5900 & n5901 ;
  assign n5903 = ~n492 & ~n5189 ;
  assign n5904 = n946 & n1630 ;
  assign n5905 = ~n5903 & n5904 ;
  assign n5906 = ~n5902 & ~n5905 ;
  assign n5907 = ~x1 & ~n5906 ;
  assign n5908 = ~x3 & ~x7 ;
  assign n5909 = n1742 & n3279 ;
  assign n5910 = n5908 & n5909 ;
  assign n5911 = ~n5907 & ~n5910 ;
  assign n5912 = n404 & n3092 ;
  assign n5913 = ~n2654 & ~n5912 ;
  assign n5914 = x3 & ~n5913 ;
  assign n5915 = ~n4462 & ~n5914 ;
  assign n5916 = n1095 & ~n5915 ;
  assign n5917 = ~n4657 & ~n5916 ;
  assign n5918 = n568 & ~n5917 ;
  assign n5919 = n718 & n4462 ;
  assign n5920 = x13 & n4359 ;
  assign n5921 = ~n4344 & ~n5920 ;
  assign n5922 = ~n5919 & n5921 ;
  assign n5923 = n1263 & n1649 ;
  assign n5924 = ~n5922 & n5923 ;
  assign n5925 = ~n5918 & ~n5924 ;
  assign n5926 = n5911 & n5925 ;
  assign n5927 = ~n5899 & n5926 ;
  assign n5928 = x11 & ~n5927 ;
  assign n5929 = ~x3 & n332 ;
  assign n5930 = ~n827 & ~n3196 ;
  assign n5931 = n5929 & ~n5930 ;
  assign n5932 = x9 & ~n3490 ;
  assign n5933 = n5931 & ~n5932 ;
  assign n5934 = n802 & n2653 ;
  assign n5935 = ~n5933 & ~n5934 ;
  assign n5936 = n55 & n5092 ;
  assign n5937 = ~n561 & ~n2848 ;
  assign n5938 = n900 & ~n5937 ;
  assign n5939 = ~n5936 & ~n5938 ;
  assign n5940 = x2 & ~n5939 ;
  assign n5941 = ~x2 & n4338 ;
  assign n5942 = n1920 & n4179 ;
  assign n5943 = n5942 ^ x1 ;
  assign n5944 = n5943 ^ n5942 ;
  assign n5945 = n5944 ^ n5941 ;
  assign n5946 = n526 & ~n1671 ;
  assign n5947 = n1423 & n1920 ;
  assign n5948 = n5947 ^ n5946 ;
  assign n5949 = ~n5946 & n5948 ;
  assign n5950 = n5949 ^ n5942 ;
  assign n5951 = n5950 ^ n5946 ;
  assign n5952 = n5945 & n5951 ;
  assign n5953 = n5952 ^ n5949 ;
  assign n5954 = n5953 ^ n5946 ;
  assign n5955 = n5941 & ~n5954 ;
  assign n5956 = n5955 ^ n5941 ;
  assign n5957 = ~n5940 & ~n5956 ;
  assign n5958 = n5935 & n5957 ;
  assign n5959 = n1169 & n2356 ;
  assign n5960 = x12 & ~n397 ;
  assign n5961 = ~n5959 & ~n5960 ;
  assign n5962 = x2 & n4338 ;
  assign n5963 = ~n5961 & n5962 ;
  assign n5964 = n395 & ~n964 ;
  assign n5965 = ~n32 & n1667 ;
  assign n5966 = ~n5964 & n5965 ;
  assign n5967 = n332 & n4797 ;
  assign n5968 = ~x2 & n718 ;
  assign n5969 = n370 & n5968 ;
  assign n5970 = ~n851 & ~n5969 ;
  assign n5971 = ~n5967 & n5970 ;
  assign n5972 = n5971 ^ x3 ;
  assign n5973 = n5972 ^ n5971 ;
  assign n5974 = n5973 ^ n5966 ;
  assign n5975 = ~n1016 & n3019 ;
  assign n5976 = ~x1 & n1270 ;
  assign n5977 = n1038 & n5976 ;
  assign n5978 = ~n668 & n5977 ;
  assign n5979 = n44 & ~n395 ;
  assign n5980 = ~n126 & n5979 ;
  assign n5981 = ~n5978 & ~n5980 ;
  assign n5982 = ~n5975 & n5981 ;
  assign n5983 = n5982 ^ x12 ;
  assign n5984 = ~x12 & n5983 ;
  assign n5985 = n5984 ^ n5971 ;
  assign n5986 = n5985 ^ x12 ;
  assign n5987 = ~n5974 & n5986 ;
  assign n5988 = n5987 ^ n5984 ;
  assign n5989 = n5988 ^ x12 ;
  assign n5990 = ~n5966 & ~n5989 ;
  assign n5991 = n5990 ^ n5966 ;
  assign n5992 = n3196 & n5991 ;
  assign n5993 = ~n5963 & ~n5992 ;
  assign n5994 = n955 & n1364 ;
  assign n5995 = n33 & n5994 ;
  assign n5996 = x2 & ~n3960 ;
  assign n5997 = n163 & n5996 ;
  assign n5998 = x3 & x15 ;
  assign n5999 = x14 & n5998 ;
  assign n6000 = n5888 & n5999 ;
  assign n6001 = ~n5997 & ~n6000 ;
  assign n6002 = n1627 & ~n6001 ;
  assign n6003 = x12 & n332 ;
  assign n6004 = ~n24 & n1708 ;
  assign n6005 = ~n6003 & ~n6004 ;
  assign n6006 = ~n6002 & n6005 ;
  assign n6007 = n858 & ~n6006 ;
  assign n6008 = ~n1317 & ~n1478 ;
  assign n6009 = n442 & n3091 ;
  assign n6010 = n6008 & n6009 ;
  assign n6011 = n2512 & ~n5584 ;
  assign n6012 = x2 & n6011 ;
  assign n6013 = ~n6010 & ~n6012 ;
  assign n6014 = ~n6007 & n6013 ;
  assign n6015 = ~n5995 & n6014 ;
  assign n6016 = n6015 ^ x5 ;
  assign n6017 = n6016 ^ n6015 ;
  assign n6018 = n6017 ^ n5993 ;
  assign n6019 = n141 & n846 ;
  assign n6020 = ~n1665 & ~n1667 ;
  assign n6021 = ~n1327 & ~n2466 ;
  assign n6022 = n332 & n6021 ;
  assign n6023 = ~n6020 & n6022 ;
  assign n6024 = n301 & n1742 ;
  assign n6025 = ~n6023 & ~n6024 ;
  assign n6026 = ~n6019 & n6025 ;
  assign n6027 = n6026 ^ x9 ;
  assign n6028 = x9 & ~n6027 ;
  assign n6029 = n6028 ^ n6015 ;
  assign n6030 = n6029 ^ x9 ;
  assign n6031 = ~n6018 & ~n6030 ;
  assign n6032 = n6031 ^ n6028 ;
  assign n6033 = n6032 ^ x9 ;
  assign n6034 = n5993 & n6033 ;
  assign n6035 = n6034 ^ n5993 ;
  assign n6036 = n845 & ~n6035 ;
  assign n6037 = x5 & x12 ;
  assign n6038 = n1025 & n6037 ;
  assign n6039 = ~x12 & n870 ;
  assign n6040 = ~n1630 & ~n6039 ;
  assign n6041 = x2 & ~n1920 ;
  assign n6042 = ~n6040 & n6041 ;
  assign n6043 = n5968 ^ n1692 ;
  assign n6044 = n6043 ^ n1692 ;
  assign n6045 = n1692 ^ x5 ;
  assign n6046 = n6045 ^ n1692 ;
  assign n6047 = n6044 & ~n6046 ;
  assign n6048 = n6047 ^ n1692 ;
  assign n6049 = ~x12 & n6048 ;
  assign n6050 = n6049 ^ n1692 ;
  assign n6051 = ~n6042 & ~n6050 ;
  assign n6052 = x7 & ~n6051 ;
  assign n6053 = n885 & n1977 ;
  assign n6054 = x5 & n6053 ;
  assign n6055 = ~n6052 & ~n6054 ;
  assign n6056 = ~n6038 & n6055 ;
  assign n6057 = n55 & ~n6056 ;
  assign n6058 = ~n328 & ~n5189 ;
  assign n6059 = ~n2848 & ~n6058 ;
  assign n6060 = n5615 & n6059 ;
  assign n6061 = n110 & ~n3196 ;
  assign n6062 = ~n526 & n6061 ;
  assign n6063 = ~n4657 & ~n6062 ;
  assign n6064 = n1282 & ~n6063 ;
  assign n6065 = n846 & n2637 ;
  assign n6066 = ~n3720 & ~n6065 ;
  assign n6067 = ~n955 & ~n3091 ;
  assign n6068 = n196 & ~n6067 ;
  assign n6069 = n1364 & n6068 ;
  assign n6070 = n6066 & ~n6069 ;
  assign n6071 = ~n6064 & n6070 ;
  assign n6072 = ~n6060 & n6071 ;
  assign n6073 = n74 & ~n6072 ;
  assign n6074 = ~n1630 & ~n5233 ;
  assign n6075 = n55 & n668 ;
  assign n6076 = ~n6074 & n6075 ;
  assign n6077 = ~n6073 & ~n6076 ;
  assign n6078 = n4793 & n5615 ;
  assign n6079 = ~n657 & n2653 ;
  assign n6080 = ~n3720 & ~n6079 ;
  assign n6081 = ~n3197 & n6080 ;
  assign n6082 = n1095 & ~n6081 ;
  assign n6083 = ~n6078 & ~n6082 ;
  assign n6084 = n348 & ~n6083 ;
  assign n6085 = n4461 & n6039 ;
  assign n6086 = n44 & n6085 ;
  assign n6087 = ~n6084 & ~n6086 ;
  assign n6088 = n6077 & n6087 ;
  assign n6089 = ~n6057 & n6088 ;
  assign n6090 = n1010 & ~n6089 ;
  assign n6091 = ~n6036 & ~n6090 ;
  assign n6092 = n5958 & n6091 ;
  assign n6093 = ~n5928 & n6092 ;
  assign n6094 = n175 & ~n6093 ;
  assign n6095 = n404 & n5976 ;
  assign n6096 = ~x3 & n6095 ;
  assign n6097 = ~x3 & n1270 ;
  assign n6098 = ~n633 & ~n6097 ;
  assign n6099 = n126 & ~n276 ;
  assign n6100 = x8 & n6099 ;
  assign n6101 = ~n6098 & n6100 ;
  assign n6102 = ~n6096 & ~n6101 ;
  assign n6103 = n3196 & ~n6102 ;
  assign n6104 = x13 & n196 ;
  assign n6105 = n1042 & n6104 ;
  assign n6106 = n263 & n6105 ;
  assign n6107 = ~n6103 & ~n6106 ;
  assign n6108 = n845 & ~n6107 ;
  assign n6109 = n348 & n634 ;
  assign n6110 = n3682 & n6109 ;
  assign n6111 = ~x9 & n4738 ;
  assign n6112 = ~n1949 & ~n6111 ;
  assign n6113 = n569 & n4359 ;
  assign n6114 = ~n6112 & n6113 ;
  assign n6115 = ~n6110 & ~n6114 ;
  assign n6116 = ~n6108 & n6115 ;
  assign n6117 = n1685 & ~n6116 ;
  assign n6118 = x11 & ~n1327 ;
  assign n6119 = n568 & ~n1095 ;
  assign n6120 = ~n4313 & ~n6119 ;
  assign n6121 = n6118 & ~n6120 ;
  assign n6122 = n946 & n4033 ;
  assign n6123 = ~n6121 & ~n6122 ;
  assign n6124 = ~x0 & n6123 ;
  assign n6125 = ~n226 & ~n2117 ;
  assign n6126 = n866 & n6125 ;
  assign n6127 = ~n261 & ~n6126 ;
  assign n6128 = ~n6124 & n6127 ;
  assign n6129 = ~x1 & n524 ;
  assign n6130 = x2 & n6129 ;
  assign n6131 = ~n6128 & ~n6130 ;
  assign n6132 = n4344 & ~n6131 ;
  assign n6133 = ~n4358 & ~n4368 ;
  assign n6134 = n2271 & ~n6133 ;
  assign n6135 = n2116 & n2653 ;
  assign n6136 = ~n978 & n1282 ;
  assign n6137 = x7 & ~n34 ;
  assign n6138 = n6136 & ~n6137 ;
  assign n6139 = ~n6135 & ~n6138 ;
  assign n6140 = ~n6134 & n6139 ;
  assign n6141 = n889 & ~n6140 ;
  assign n6142 = ~n1113 & n2512 ;
  assign n6143 = n85 & n6142 ;
  assign n6144 = ~n489 & n6143 ;
  assign n6145 = n2413 & n6144 ;
  assign n6146 = ~x7 & n1656 ;
  assign n6147 = ~n4286 & ~n6146 ;
  assign n6148 = n6147 ^ x5 ;
  assign n6149 = n6148 ^ n6147 ;
  assign n6150 = ~x7 & n1282 ;
  assign n6151 = n6150 ^ n6147 ;
  assign n6152 = n6149 & ~n6151 ;
  assign n6153 = n6152 ^ n6147 ;
  assign n6154 = n1114 & ~n6153 ;
  assign n6155 = ~n6145 & ~n6154 ;
  assign n6156 = ~n6141 & n6155 ;
  assign n6157 = n38 & ~n6156 ;
  assign n6158 = n828 & n4314 ;
  assign n6159 = ~n371 & ~n6158 ;
  assign n6160 = ~n759 & ~n1247 ;
  assign n6161 = ~n2291 & n6160 ;
  assign n6162 = ~n6159 & ~n6161 ;
  assign n6163 = n60 & n1226 ;
  assign n6164 = n889 & n6163 ;
  assign n6165 = ~n6162 & ~n6164 ;
  assign n6166 = n4561 & ~n6165 ;
  assign n6167 = x3 & n6166 ;
  assign n6168 = x5 & n462 ;
  assign n6169 = ~n2510 & ~n5206 ;
  assign n6170 = x13 & ~n2510 ;
  assign n6171 = ~n6169 & ~n6170 ;
  assign n6172 = n6168 & n6171 ;
  assign n6173 = n2312 & n2901 ;
  assign n6174 = n900 & n6173 ;
  assign n6175 = ~n6172 & ~n6174 ;
  assign n6176 = n6175 ^ n1246 ;
  assign n6177 = n6176 ^ n6175 ;
  assign n6178 = n6175 ^ n5210 ;
  assign n6179 = n6178 ^ n6175 ;
  assign n6180 = n6177 & n6179 ;
  assign n6181 = n6180 ^ n6175 ;
  assign n6182 = ~x0 & ~n6181 ;
  assign n6183 = n6182 ^ n6175 ;
  assign n6184 = ~n6167 & n6183 ;
  assign n6185 = ~n6157 & n6184 ;
  assign n6186 = n6185 ^ x5 ;
  assign n6187 = n6186 ^ n6185 ;
  assign n6188 = ~x13 & n5189 ;
  assign n6189 = ~x12 & n749 ;
  assign n6190 = ~n2398 & ~n6189 ;
  assign n6191 = n6188 & ~n6190 ;
  assign n6192 = n1042 & n3172 ;
  assign n6193 = ~n6191 & ~n6192 ;
  assign n6194 = n60 & ~n6193 ;
  assign n6195 = x1 & n224 ;
  assign n6196 = n2601 & n6195 ;
  assign n6197 = x12 & n6196 ;
  assign n6198 = ~n6194 & ~n6197 ;
  assign n6199 = n6198 ^ n6185 ;
  assign n6200 = n6199 ^ n6185 ;
  assign n6201 = ~n6187 & ~n6200 ;
  assign n6202 = n6201 ^ n6185 ;
  assign n6203 = x2 & ~n6202 ;
  assign n6204 = n6203 ^ n6185 ;
  assign n6205 = ~n6132 & n6204 ;
  assign n6206 = n282 & ~n6205 ;
  assign n6207 = ~n6117 & ~n6206 ;
  assign n6208 = ~n6094 & n6207 ;
  assign n6209 = n453 & n4002 ;
  assign n6210 = n1478 & n6209 ;
  assign n6242 = n19 & n2653 ;
  assign n6243 = ~n4223 & ~n6242 ;
  assign n6244 = n4201 & ~n6243 ;
  assign n6245 = ~n947 & n6244 ;
  assign n6246 = n28 & n946 ;
  assign n6247 = ~n2583 & n6246 ;
  assign n6248 = n74 & n3091 ;
  assign n6249 = ~x10 & n6248 ;
  assign n6250 = ~n76 & ~n2557 ;
  assign n6251 = n1007 & ~n6250 ;
  assign n6252 = ~n6249 & ~n6251 ;
  assign n6253 = ~n6247 & n6252 ;
  assign n6254 = ~x5 & ~n6253 ;
  assign n6255 = ~n690 & n1061 ;
  assign n6256 = n5889 & ~n6255 ;
  assign n6257 = ~n6254 & ~n6256 ;
  assign n6258 = ~n6245 & n6257 ;
  assign n6211 = ~x2 & n2653 ;
  assign n6212 = ~n4793 & ~n6211 ;
  assign n6213 = n142 & n473 ;
  assign n6214 = ~n6212 & n6213 ;
  assign n6215 = n6214 ^ x14 ;
  assign n6216 = n679 & n2653 ;
  assign n6217 = ~n890 & n6216 ;
  assign n6218 = n213 & ~n622 ;
  assign n6219 = ~n473 & n6218 ;
  assign n6220 = ~n6217 & ~n6219 ;
  assign n6221 = n6220 ^ x1 ;
  assign n6222 = n6221 ^ n6220 ;
  assign n6223 = ~x15 & ~n176 ;
  assign n6224 = n622 & ~n6223 ;
  assign n6225 = n473 & n3568 ;
  assign n6226 = ~n6224 & ~n6225 ;
  assign n6227 = x5 & ~n6226 ;
  assign n6228 = n981 ^ x13 ;
  assign n6229 = n213 & ~n6228 ;
  assign n6230 = ~n6227 & ~n6229 ;
  assign n6231 = n6230 ^ n6220 ;
  assign n6232 = n6222 & n6231 ;
  assign n6233 = n6232 ^ n6220 ;
  assign n6234 = n6233 ^ n6214 ;
  assign n6235 = ~n6215 & n6234 ;
  assign n6236 = n6235 ^ n6232 ;
  assign n6237 = n6236 ^ n6220 ;
  assign n6238 = n6237 ^ x14 ;
  assign n6239 = ~n6214 & ~n6238 ;
  assign n6240 = n6239 ^ n6214 ;
  assign n6241 = n6240 ^ n6214 ;
  assign n6259 = n6258 ^ n6241 ;
  assign n6260 = x0 & n6259 ;
  assign n6261 = n6260 ^ n6241 ;
  assign n6262 = ~n6210 & n6261 ;
  assign n6263 = n1665 & ~n6262 ;
  assign n6264 = ~n489 & ~n4313 ;
  assign n6265 = n1095 & ~n6264 ;
  assign n6266 = n332 & ~n371 ;
  assign n6267 = n381 & ~n1327 ;
  assign n6268 = n6266 & ~n6267 ;
  assign n6269 = ~n6265 & ~n6268 ;
  assign n6270 = n4461 & ~n6269 ;
  assign n6271 = n4470 & n6037 ;
  assign n6272 = n1645 & n6271 ;
  assign n6273 = x11 & ~n6272 ;
  assign n6274 = ~n6270 & n6273 ;
  assign n6275 = ~n6263 & n6274 ;
  assign n6276 = ~x2 & n827 ;
  assign n6277 = n2356 & n6276 ;
  assign n6278 = ~x10 & n1146 ;
  assign n6279 = ~n6277 & ~n6278 ;
  assign n6280 = n261 & ~n6279 ;
  assign n6281 = n6280 ^ x7 ;
  assign n6282 = n3019 & n4313 ;
  assign n6283 = ~n673 & n1380 ;
  assign n6284 = ~n557 & n6283 ;
  assign n6285 = n28 & n4201 ;
  assign n6286 = x10 & ~n5516 ;
  assign n6287 = ~n29 & n6286 ;
  assign n6288 = ~n6285 & ~n6287 ;
  assign n6289 = n364 & ~n6288 ;
  assign n6290 = ~n6284 & ~n6289 ;
  assign n6291 = ~n6282 & n6290 ;
  assign n6292 = n6291 ^ x0 ;
  assign n6293 = n6292 ^ n6291 ;
  assign n6294 = ~n828 & ~n1282 ;
  assign n6295 = ~n28 & ~n6294 ;
  assign n6296 = n946 & n6295 ;
  assign n6297 = n6283 ^ x2 ;
  assign n6298 = n6297 ^ n6283 ;
  assign n6299 = n6283 ^ n1977 ;
  assign n6300 = n6299 ^ n6283 ;
  assign n6301 = ~n6298 & n6300 ;
  assign n6302 = n6301 ^ n6283 ;
  assign n6303 = x10 & n6302 ;
  assign n6304 = n6303 ^ n6283 ;
  assign n6305 = ~n6296 & ~n6304 ;
  assign n6306 = n6305 ^ n6291 ;
  assign n6307 = n6293 & n6306 ;
  assign n6308 = n6307 ^ n6291 ;
  assign n6309 = n6308 ^ n6280 ;
  assign n6310 = n6281 & n6309 ;
  assign n6311 = n6310 ^ n6307 ;
  assign n6312 = n6311 ^ n6291 ;
  assign n6313 = n6312 ^ x7 ;
  assign n6314 = ~n6280 & n6313 ;
  assign n6315 = n6314 ^ n6280 ;
  assign n6316 = n6315 ^ n6280 ;
  assign n6317 = n561 & ~n6316 ;
  assign n6318 = n57 & n1702 ;
  assign n6319 = x0 & ~n79 ;
  assign n6320 = ~n1349 & n6319 ;
  assign n6321 = ~n6318 & ~n6320 ;
  assign n6322 = n6276 & ~n6321 ;
  assign n6323 = x1 & n5233 ;
  assign n6324 = ~n3306 & ~n6323 ;
  assign n6325 = n1682 & ~n6324 ;
  assign n6326 = n60 & n4253 ;
  assign n6327 = n497 & n6326 ;
  assign n6328 = ~n164 & ~n4253 ;
  assign n6329 = n2271 & n6328 ;
  assign n6330 = ~n6327 & ~n6329 ;
  assign n6331 = ~n6325 & n6330 ;
  assign n6332 = n946 & ~n6331 ;
  assign n6333 = n20 & n1060 ;
  assign n6334 = n3197 & n6333 ;
  assign n6335 = n827 & n1617 ;
  assign n6336 = n1383 & n3490 ;
  assign n6337 = ~n6335 & ~n6336 ;
  assign n6338 = ~n6334 & n6337 ;
  assign n6339 = ~n6332 & n6338 ;
  assign n6340 = ~n6322 & n6339 ;
  assign n6341 = ~x3 & ~n6340 ;
  assign n6342 = ~n6317 & ~n6341 ;
  assign n6343 = n6275 & n6342 ;
  assign n6344 = n328 & n5284 ;
  assign n6345 = ~n750 & n1002 ;
  assign n6346 = x10 & n6345 ;
  assign n6347 = ~n6344 & ~n6346 ;
  assign n6348 = ~x2 & n6037 ;
  assign n6349 = ~n6347 & n6348 ;
  assign n6350 = n39 & n3263 ;
  assign n6351 = n314 & n6350 ;
  assign n6352 = n232 & n363 ;
  assign n6353 = n163 & n6352 ;
  assign n6354 = ~n6351 & ~n6353 ;
  assign n6355 = x15 & n3914 ;
  assign n6356 = ~n6354 & n6355 ;
  assign n6357 = n561 & n6150 ;
  assign n6358 = n2873 & ~n6250 ;
  assign n6359 = ~n828 & ~n2466 ;
  assign n6360 = x7 & ~n1641 ;
  assign n6361 = n6359 & n6360 ;
  assign n6362 = ~n6358 & ~n6361 ;
  assign n6363 = ~x3 & ~n6362 ;
  assign n6364 = ~n6357 & ~n6363 ;
  assign n6365 = n3330 & ~n6364 ;
  assign n6366 = ~n3306 & ~n6188 ;
  assign n6367 = ~n168 & ~n1658 ;
  assign n6368 = ~n6366 & n6367 ;
  assign n6369 = x10 & n4344 ;
  assign n6370 = n6021 & n6369 ;
  assign n6371 = ~x5 & n846 ;
  assign n6372 = n1905 & n6371 ;
  assign n6373 = x12 & n168 ;
  assign n6374 = n981 & n6373 ;
  assign n6375 = ~n6372 & ~n6374 ;
  assign n6376 = ~n6370 & n6375 ;
  assign n6377 = ~n6368 & n6376 ;
  assign n6378 = n20 & ~n6377 ;
  assign n6379 = ~n6365 & ~n6378 ;
  assign n6380 = n3092 ^ x12 ;
  assign n6381 = n3092 ^ x10 ;
  assign n6382 = n6381 ^ x10 ;
  assign n6383 = n3682 ^ x10 ;
  assign n6384 = ~n6382 & n6383 ;
  assign n6385 = n6384 ^ x10 ;
  assign n6386 = ~n6380 & ~n6385 ;
  assign n6387 = n6386 ^ x12 ;
  assign n6388 = n110 & ~n6387 ;
  assign n6389 = x7 & n5431 ;
  assign n6390 = ~n6388 & ~n6389 ;
  assign n6391 = n740 & ~n6390 ;
  assign n6392 = n196 & n928 ;
  assign n6393 = n1270 & n6392 ;
  assign n6394 = n2876 & n6393 ;
  assign n6395 = n1682 & n4782 ;
  assign n6396 = n405 & n6395 ;
  assign n6397 = ~n6394 & ~n6396 ;
  assign n6398 = ~n6391 & n6397 ;
  assign n6399 = n6379 & n6398 ;
  assign n6400 = ~n6356 & n6399 ;
  assign n6401 = n6400 ^ x1 ;
  assign n6402 = n6401 ^ n6400 ;
  assign n6447 = n712 & n955 ;
  assign n6448 = ~n314 & ~n328 ;
  assign n6449 = n4656 & ~n6448 ;
  assign n6450 = ~n1667 & ~n6449 ;
  assign n6451 = n6447 & ~n6450 ;
  assign n6452 = n311 & n1214 ;
  assign n6453 = n5941 & n6452 ;
  assign n6454 = n2512 & n3019 ;
  assign n6455 = ~n6453 & ~n6454 ;
  assign n6456 = n6455 ^ x5 ;
  assign n6457 = n6456 ^ n6455 ;
  assign n6458 = n6457 ^ n6451 ;
  assign n6459 = ~x7 & n1353 ;
  assign n6460 = ~n3019 & ~n6459 ;
  assign n6461 = n6460 ^ n1667 ;
  assign n6462 = ~n6460 & ~n6461 ;
  assign n6463 = n6462 ^ n6455 ;
  assign n6464 = n6463 ^ n6460 ;
  assign n6465 = n6458 & n6464 ;
  assign n6466 = n6465 ^ n6462 ;
  assign n6467 = n6466 ^ n6460 ;
  assign n6468 = ~n6451 & ~n6467 ;
  assign n6469 = n6468 ^ n6451 ;
  assign n6403 = ~n24 & n1686 ;
  assign n6404 = ~n561 & ~n650 ;
  assign n6405 = x7 & n6404 ;
  assign n6406 = n6403 & n6405 ;
  assign n6407 = n6037 ^ x0 ;
  assign n6408 = n6407 ^ n919 ;
  assign n6409 = n2362 ^ n328 ;
  assign n6410 = x0 & ~n6409 ;
  assign n6411 = n6410 ^ n328 ;
  assign n6412 = n6408 & n6411 ;
  assign n6413 = n6412 ^ n6410 ;
  assign n6414 = n6413 ^ n328 ;
  assign n6415 = n6414 ^ x0 ;
  assign n6416 = n919 & n6415 ;
  assign n6417 = ~n6406 & ~n6416 ;
  assign n6418 = x2 ^ x0 ;
  assign n6419 = n6418 ^ x2 ;
  assign n6420 = n4005 ^ x2 ;
  assign n6421 = ~n6419 & ~n6420 ;
  assign n6422 = n6421 ^ x2 ;
  assign n6423 = ~x2 & n1282 ;
  assign n6424 = n6423 ^ n4359 ;
  assign n6425 = ~n6422 & n6424 ;
  assign n6426 = n6425 ^ n6423 ;
  assign n6427 = n4359 & n6426 ;
  assign n6428 = n6427 ^ n4359 ;
  assign n6429 = n6428 ^ n4359 ;
  assign n6430 = n6417 & ~n6429 ;
  assign n6470 = n6469 ^ n6430 ;
  assign n6431 = n561 & ~n6250 ;
  assign n6432 = x13 & n4461 ;
  assign n6433 = ~n3192 & ~n6432 ;
  assign n6434 = ~n6431 & n6433 ;
  assign n6435 = n364 & ~n6434 ;
  assign n6436 = ~x2 & n3030 ;
  assign n6437 = ~n311 & ~n5996 ;
  assign n6438 = n1978 & ~n6437 ;
  assign n6439 = ~n6436 & ~n6438 ;
  assign n6440 = n4338 & ~n6439 ;
  assign n6441 = n1667 & n3196 ;
  assign n6442 = n1271 & n4359 ;
  assign n6443 = ~n6441 & ~n6442 ;
  assign n6444 = ~n6440 & n6443 ;
  assign n6445 = ~n6435 & n6444 ;
  assign n6446 = n6445 ^ n6430 ;
  assign n6471 = n6470 ^ n6446 ;
  assign n6472 = n6446 ^ x0 ;
  assign n6473 = n6472 ^ n6446 ;
  assign n6474 = ~n6471 & ~n6473 ;
  assign n6475 = n6474 ^ n6446 ;
  assign n6476 = ~x10 & n6475 ;
  assign n6477 = n6476 ^ n6430 ;
  assign n6478 = n6477 ^ n6400 ;
  assign n6479 = ~n6402 & n6478 ;
  assign n6480 = n6479 ^ n6400 ;
  assign n6481 = ~n6349 & n6480 ;
  assign n6482 = ~x11 & n6481 ;
  assign n6483 = ~n6343 & ~n6482 ;
  assign n6514 = n712 & n1002 ;
  assign n6515 = x0 & ~n6212 ;
  assign n6516 = ~n6514 & ~n6515 ;
  assign n6517 = n5590 & ~n6516 ;
  assign n6484 = ~x0 & n65 ;
  assign n6485 = n828 & n5012 ;
  assign n6486 = x1 & n2902 ;
  assign n6487 = ~n2873 & n6486 ;
  assign n6488 = ~n6485 & ~n6487 ;
  assign n6489 = n6484 & ~n6488 ;
  assign n6490 = x3 & n58 ;
  assign n6491 = ~n1672 & ~n6490 ;
  assign n6492 = ~n348 & ~n6491 ;
  assign n6493 = n6492 ^ x5 ;
  assign n6494 = n6493 ^ n6492 ;
  assign n6495 = n6494 ^ n6489 ;
  assign n6496 = ~x2 & ~n2362 ;
  assign n6497 = n4253 & ~n6496 ;
  assign n6498 = n141 ^ x3 ;
  assign n6499 = n6498 ^ n141 ;
  assign n6500 = n142 ^ n141 ;
  assign n6501 = n6499 & n6500 ;
  assign n6502 = n6501 ^ n141 ;
  assign n6503 = x7 & n6502 ;
  assign n6504 = ~n6497 & ~n6503 ;
  assign n6505 = n6504 ^ x0 ;
  assign n6506 = ~n6504 & ~n6505 ;
  assign n6507 = n6506 ^ n6492 ;
  assign n6508 = n6507 ^ n6504 ;
  assign n6509 = ~n6495 & ~n6508 ;
  assign n6510 = n6509 ^ n6506 ;
  assign n6511 = n6510 ^ n6504 ;
  assign n6512 = ~n6489 & ~n6511 ;
  assign n6513 = n6512 ^ n6489 ;
  assign n6518 = n6517 ^ n6513 ;
  assign n6519 = ~x10 & n6518 ;
  assign n6520 = n6519 ^ n6513 ;
  assign n6521 = ~n6483 & ~n6520 ;
  assign n6522 = n265 & ~n6521 ;
  assign n6523 = n383 & n885 ;
  assign n6524 = n4628 & n6523 ;
  assign n6525 = n900 & n6524 ;
  assign n6526 = ~n6522 & ~n6525 ;
  assign n6527 = n6208 & n6526 ;
  assign n6528 = n1665 & n4494 ;
  assign n6529 = n3490 & n6528 ;
  assign n6530 = ~n5713 & n5999 ;
  assign n6531 = n1202 & n1247 ;
  assign n6532 = n328 & n3177 ;
  assign n6533 = ~n6531 & ~n6532 ;
  assign n6534 = ~n6530 & n6533 ;
  assign n6535 = n2653 & ~n6534 ;
  assign n6536 = ~n6529 & ~n6535 ;
  assign n6537 = n396 & ~n6536 ;
  assign n6538 = n2329 & n3294 ;
  assign n6539 = n1202 & n6538 ;
  assign n6540 = n3030 & n6539 ;
  assign n6541 = ~n6537 & ~n6540 ;
  assign n6542 = n928 & ~n6541 ;
  assign n6543 = n472 & n848 ;
  assign n6544 = ~n1684 & n4462 ;
  assign n6545 = n6543 & n6544 ;
  assign n6546 = n1762 & ~n5772 ;
  assign n6547 = n2711 & n4710 ;
  assign n6548 = ~n4461 & ~n6547 ;
  assign n6549 = n1672 & ~n6548 ;
  assign n6550 = ~n6546 & ~n6549 ;
  assign n6551 = ~n6545 & n6550 ;
  assign n6552 = n4974 & n6111 ;
  assign n6553 = n290 & n768 ;
  assign n6554 = n4978 & n6553 ;
  assign n6555 = ~n6552 & ~n6554 ;
  assign n6556 = ~x12 & ~n6555 ;
  assign n6557 = ~n5770 & ~n6556 ;
  assign n6558 = ~n947 & ~n6557 ;
  assign n6559 = ~x0 & n6558 ;
  assign n6560 = n6551 & ~n6559 ;
  assign n6561 = ~n6542 & n6560 ;
  assign n6562 = ~x3 & n20 ;
  assign n6563 = x7 & n164 ;
  assign n6564 = n2115 & n6563 ;
  assign n6565 = n2115 & n2653 ;
  assign n6566 = ~n24 & n6565 ;
  assign n6567 = ~n4195 & ~n6566 ;
  assign n6568 = ~x1 & ~n6567 ;
  assign n6569 = ~n6564 & ~n6568 ;
  assign n6570 = n6562 & ~n6569 ;
  assign n6571 = n1010 & n4462 ;
  assign n6572 = n2115 & n4461 ;
  assign n6573 = ~n6571 & ~n6572 ;
  assign n6574 = ~x0 & n332 ;
  assign n6575 = ~n6573 & n6574 ;
  assign n6576 = ~n768 & n2228 ;
  assign n6577 = n529 & n6576 ;
  assign n6578 = n6211 & n6577 ;
  assign n6579 = ~n6575 & ~n6578 ;
  assign n6580 = ~n6570 & n6579 ;
  assign n6581 = ~n987 & ~n2601 ;
  assign n6582 = n141 & ~n6581 ;
  assign n6583 = n1042 & n3283 ;
  assign n6584 = n6583 ^ x2 ;
  assign n6585 = n6584 ^ n6583 ;
  assign n6586 = n6585 ^ n6582 ;
  assign n6587 = n1010 ^ x7 ;
  assign n6588 = n1010 & ~n6587 ;
  assign n6589 = n6588 ^ n6583 ;
  assign n6590 = n6589 ^ n1010 ;
  assign n6591 = n6586 & n6590 ;
  assign n6592 = n6591 ^ n6588 ;
  assign n6593 = n6592 ^ n1010 ;
  assign n6594 = ~n6582 & n6593 ;
  assign n6595 = n6594 ^ n6582 ;
  assign n6596 = n3532 & n6595 ;
  assign n6597 = x11 & ~x15 ;
  assign n6598 = n6447 & ~n6597 ;
  assign n6599 = n176 & n4392 ;
  assign n6600 = ~n6598 & ~n6599 ;
  assign n6601 = n453 & ~n6600 ;
  assign n6602 = ~x5 & n982 ;
  assign n6603 = ~n3682 & ~n6602 ;
  assign n6604 = n197 & ~n6603 ;
  assign n6605 = ~n74 & ~n4253 ;
  assign n6606 = n329 & ~n6605 ;
  assign n6607 = ~n947 & n6606 ;
  assign n6608 = ~n1042 & ~n2848 ;
  assign n6609 = n1524 & ~n6608 ;
  assign n6610 = x10 & n6609 ;
  assign n6611 = ~n6607 & ~n6610 ;
  assign n6612 = ~n6604 & n6611 ;
  assign n6613 = n874 & ~n6612 ;
  assign n6614 = ~n6601 & ~n6613 ;
  assign n6615 = n1282 & ~n6614 ;
  assign n6616 = ~n828 & n1060 ;
  assign n6617 = ~x12 & n1954 ;
  assign n6618 = ~n6616 & ~n6617 ;
  assign n6619 = n4793 & n6618 ;
  assign n6620 = n105 & n1627 ;
  assign n6621 = ~x0 & ~n248 ;
  assign n6622 = ~n6620 & ~n6621 ;
  assign n6623 = ~n1743 & n6622 ;
  assign n6624 = n6619 & n6623 ;
  assign n6625 = ~n471 & n6624 ;
  assign n6626 = ~n6615 & ~n6625 ;
  assign n6627 = ~n6596 & n6626 ;
  assign n6628 = n712 & n2678 ;
  assign n6629 = x11 & n6628 ;
  assign n6630 = ~n1062 & ~n4471 ;
  assign n6631 = n213 & ~n6630 ;
  assign n6632 = n511 & n2280 ;
  assign n6633 = ~n3490 & ~n6632 ;
  assign n6634 = n919 & ~n6633 ;
  assign n6635 = ~n180 & ~n2653 ;
  assign n6636 = n524 & n6635 ;
  assign n6637 = ~n6634 & ~n6636 ;
  assign n6638 = x13 & ~n6637 ;
  assign n6639 = ~n6631 & ~n6638 ;
  assign n6640 = ~n6629 & n6639 ;
  assign n6641 = n1349 & ~n6640 ;
  assign n6642 = ~n2477 & n6350 ;
  assign n6643 = n240 & n862 ;
  assign n6644 = n6643 ^ n3711 ;
  assign n6645 = n6644 ^ n3711 ;
  assign n6646 = n3711 ^ x5 ;
  assign n6647 = n6646 ^ n3711 ;
  assign n6648 = n6645 & n6647 ;
  assign n6649 = n6648 ^ n3711 ;
  assign n6650 = x10 & n6649 ;
  assign n6651 = n6650 ^ n3711 ;
  assign n6652 = ~n6642 & ~n6651 ;
  assign n6653 = n1382 & ~n6652 ;
  assign n6654 = ~n511 & n2653 ;
  assign n6655 = n141 & ~n3490 ;
  assign n6656 = ~n827 & n6655 ;
  assign n6657 = ~n6654 & n6656 ;
  assign n6658 = ~x11 & ~n6657 ;
  assign n6659 = ~n2653 & ~n4253 ;
  assign n6660 = ~n126 & ~n6659 ;
  assign n6661 = ~x12 & ~n471 ;
  assign n6662 = ~n6660 & n6661 ;
  assign n6663 = ~n6658 & n6662 ;
  assign n6664 = n6663 ^ n2653 ;
  assign n6665 = n6664 ^ n6653 ;
  assign n6666 = n1062 & n4350 ;
  assign n6667 = n6666 ^ n176 ;
  assign n6668 = ~n2653 & ~n6667 ;
  assign n6669 = n6668 ^ n6666 ;
  assign n6670 = ~n6665 & ~n6669 ;
  assign n6671 = n6670 ^ n6668 ;
  assign n6672 = n6671 ^ n6666 ;
  assign n6673 = n6672 ^ n2653 ;
  assign n6674 = ~n6653 & n6673 ;
  assign n6675 = ~n6641 & n6674 ;
  assign n6676 = n60 & ~n6675 ;
  assign n6677 = n6627 & ~n6676 ;
  assign n6678 = n492 & ~n6677 ;
  assign n6679 = n6580 & ~n6678 ;
  assign n6680 = n6679 ^ x8 ;
  assign n6681 = n6680 ^ n6679 ;
  assign n6682 = n6681 ^ n6561 ;
  assign n6796 = n1692 & n2115 ;
  assign n6797 = ~n2637 & n3490 ;
  assign n6798 = ~n3720 & ~n6797 ;
  assign n6799 = ~n2653 & n6798 ;
  assign n6800 = ~n6796 & n6799 ;
  assign n6801 = ~x3 & ~n6800 ;
  assign n6802 = ~n5190 & ~n6801 ;
  assign n6785 = n4470 & n6118 ;
  assign n6786 = ~n2480 & ~n6785 ;
  assign n6787 = n561 & ~n6786 ;
  assign n6788 = ~n276 & n2653 ;
  assign n6789 = n471 & ~n1977 ;
  assign n6790 = ~n5191 & ~n6789 ;
  assign n6791 = ~n4462 & ~n6790 ;
  assign n6792 = ~n6788 & n6791 ;
  assign n6793 = ~n6787 & n6792 ;
  assign n6683 = ~n2116 & n3720 ;
  assign n6684 = ~n1464 & ~n2654 ;
  assign n6685 = ~n6683 & n6684 ;
  assign n6686 = n568 & ~n6685 ;
  assign n6687 = n6686 ^ n3961 ;
  assign n6737 = n634 & n3286 ;
  assign n6738 = n1630 & ~n2601 ;
  assign n6739 = ~n2637 & n6738 ;
  assign n6740 = n2290 & ~n2637 ;
  assign n6741 = n85 & ~n2557 ;
  assign n6742 = n6740 & n6741 ;
  assign n6743 = ~n6739 & ~n6742 ;
  assign n6744 = n5286 & n6037 ;
  assign n6745 = n6743 & ~n6744 ;
  assign n6746 = ~n6737 & n6745 ;
  assign n6688 = ~n1382 & n3196 ;
  assign n6689 = ~n126 & n6688 ;
  assign n6690 = ~n6563 & ~n6689 ;
  assign n6691 = n346 & ~n6690 ;
  assign n6692 = ~x5 & n2512 ;
  assign n6693 = ~n673 & n2389 ;
  assign n6694 = ~n462 & ~n1458 ;
  assign n6695 = ~n6693 & n6694 ;
  assign n6696 = n6692 & ~n6695 ;
  assign n6697 = n3091 & ~n3130 ;
  assign n6698 = n1703 & n5291 ;
  assign n6699 = n6697 & n6698 ;
  assign n6700 = ~n6696 & ~n6699 ;
  assign n6701 = ~n6691 & n6700 ;
  assign n6747 = n6746 ^ n6701 ;
  assign n6702 = ~n2374 & ~n2512 ;
  assign n6703 = n1435 & ~n6702 ;
  assign n6704 = n1977 ^ x9 ;
  assign n6705 = n6704 ^ n2901 ;
  assign n6706 = n6705 ^ n1977 ;
  assign n6707 = n6706 ^ n6705 ;
  assign n6708 = n6707 ^ n6704 ;
  assign n6709 = ~n2653 & n6074 ;
  assign n6710 = n6705 ^ n6704 ;
  assign n6711 = n6707 & n6710 ;
  assign n6712 = n6711 ^ n6708 ;
  assign n6713 = n6709 & n6712 ;
  assign n6714 = n6713 ^ n6711 ;
  assign n6715 = n6708 & n6714 ;
  assign n6716 = n6715 ^ n6711 ;
  assign n6717 = n6716 ^ x9 ;
  assign n6721 = n6717 ^ n6250 ;
  assign n6722 = n6721 ^ n6717 ;
  assign n6718 = ~n3192 & ~n3728 ;
  assign n6719 = n6718 ^ n6717 ;
  assign n6720 = n6719 ^ n6717 ;
  assign n6723 = n6722 ^ n6720 ;
  assign n6724 = n6717 ^ x12 ;
  assign n6725 = n6724 ^ n6717 ;
  assign n6726 = n6725 ^ n6722 ;
  assign n6727 = ~n6722 & n6726 ;
  assign n6728 = n6727 ^ n6722 ;
  assign n6729 = n6723 & ~n6728 ;
  assign n6730 = n6729 ^ n6727 ;
  assign n6731 = n6730 ^ n6717 ;
  assign n6732 = n6731 ^ n6722 ;
  assign n6733 = ~x11 & ~n6732 ;
  assign n6734 = n6733 ^ n6717 ;
  assign n6735 = ~n6703 & ~n6734 ;
  assign n6736 = n6735 ^ n6701 ;
  assign n6748 = n6747 ^ n6736 ;
  assign n6749 = n6736 ^ x1 ;
  assign n6750 = n6749 ^ n6736 ;
  assign n6751 = n6748 & n6750 ;
  assign n6752 = n6751 ^ n6736 ;
  assign n6753 = ~x3 & n6752 ;
  assign n6754 = n6753 ^ n6701 ;
  assign n6755 = n6754 ^ x10 ;
  assign n6756 = n6755 ^ n6754 ;
  assign n6759 = n2901 ^ x3 ;
  assign n6760 = n6759 ^ x3 ;
  assign n6757 = n2083 ^ x3 ;
  assign n6758 = n6757 ^ x3 ;
  assign n6761 = n6760 ^ n6758 ;
  assign n6762 = ~n1435 & ~n1978 ;
  assign n6763 = n6762 ^ x3 ;
  assign n6764 = n6763 ^ x3 ;
  assign n6765 = n6764 ^ n6760 ;
  assign n6766 = ~n6760 & ~n6765 ;
  assign n6767 = n6766 ^ n6760 ;
  assign n6768 = ~n6761 & ~n6767 ;
  assign n6769 = n6768 ^ n6766 ;
  assign n6770 = n6769 ^ x3 ;
  assign n6771 = n6770 ^ n6760 ;
  assign n6772 = ~n2848 & n6771 ;
  assign n6773 = n6772 ^ x3 ;
  assign n6774 = ~n1869 & n6773 ;
  assign n6775 = n6774 ^ n6754 ;
  assign n6776 = n6756 & n6775 ;
  assign n6777 = n6776 ^ n6754 ;
  assign n6778 = n6777 ^ n6686 ;
  assign n6779 = n6687 & ~n6778 ;
  assign n6780 = n6779 ^ n6776 ;
  assign n6781 = n6780 ^ n6754 ;
  assign n6782 = n6781 ^ n3961 ;
  assign n6783 = ~n6686 & ~n6782 ;
  assign n6784 = n6783 ^ n6686 ;
  assign n6794 = n6793 ^ n6784 ;
  assign n6795 = n6794 ^ n6793 ;
  assign n6803 = n6802 ^ n6795 ;
  assign n6804 = n6803 ^ n6794 ;
  assign n6805 = n6794 ^ x1 ;
  assign n6806 = n6805 ^ n6794 ;
  assign n6807 = n6804 & n6806 ;
  assign n6808 = n6807 ^ n6794 ;
  assign n6809 = x2 & ~n6808 ;
  assign n6810 = n6809 ^ n6784 ;
  assign n6811 = n6810 ^ x0 ;
  assign n6812 = x0 & n6811 ;
  assign n6813 = n6812 ^ n6679 ;
  assign n6814 = n6813 ^ x0 ;
  assign n6815 = n6682 & ~n6814 ;
  assign n6816 = n6815 ^ n6812 ;
  assign n6817 = n6816 ^ x0 ;
  assign n6818 = n6561 & n6817 ;
  assign n6819 = n6818 ^ n6561 ;
  assign n6820 = n6527 & n6819 ;
  assign n6821 = x4 & ~n6820 ;
  assign n6822 = ~n3561 & ~n4330 ;
  assign n6823 = ~n467 & ~n6822 ;
  assign n6824 = ~x7 & ~x15 ;
  assign n6825 = n1716 & ~n6824 ;
  assign n6826 = n4605 & n6825 ;
  assign n6827 = n1290 & n1806 ;
  assign n6828 = n2678 & n6827 ;
  assign n6829 = ~n6826 & ~n6828 ;
  assign n6830 = ~x0 & ~n6829 ;
  assign n6831 = n1050 & n1559 ;
  assign n6832 = n1509 & n6831 ;
  assign n6833 = ~n6830 & ~n6832 ;
  assign n6834 = n6823 & ~n6833 ;
  assign n6835 = n145 & n1910 ;
  assign n6836 = x8 & n2738 ;
  assign n6837 = ~n6835 & ~n6836 ;
  assign n6838 = ~n1092 & ~n6837 ;
  assign n6839 = n1478 ^ x14 ;
  assign n6840 = n6839 ^ n1478 ;
  assign n6841 = n1478 ^ n964 ;
  assign n6842 = n6841 ^ n1478 ;
  assign n6843 = n6840 & n6842 ;
  assign n6844 = n6843 ^ n1478 ;
  assign n6845 = x0 & n6844 ;
  assign n6846 = n6845 ^ n1478 ;
  assign n6847 = n426 & n6846 ;
  assign n6848 = ~x11 & n6847 ;
  assign n6849 = ~n6838 & ~n6848 ;
  assign n6850 = n3104 & ~n6849 ;
  assign n6851 = n310 & n5189 ;
  assign n6852 = n6835 & n6851 ;
  assign n6853 = x15 & n5180 ;
  assign n6854 = ~n3785 & ~n6853 ;
  assign n6855 = ~x2 & n955 ;
  assign n6856 = n623 & n6855 ;
  assign n6857 = ~n6854 & n6856 ;
  assign n6858 = n348 & n6857 ;
  assign n6859 = ~n6852 & ~n6858 ;
  assign n6860 = ~n6850 & n6859 ;
  assign n6861 = ~x5 & ~n6860 ;
  assign n6862 = ~x4 & n1565 ;
  assign n6863 = n826 & n6862 ;
  assign n6864 = n74 & n6097 ;
  assign n6865 = n1692 & n6864 ;
  assign n6866 = ~n6863 & ~n6865 ;
  assign n6867 = n978 & n3424 ;
  assign n6868 = ~n6866 & n6867 ;
  assign n6869 = ~n6861 & ~n6868 ;
  assign n6870 = ~n1658 & ~n6869 ;
  assign n6871 = n465 & n740 ;
  assign n6872 = n784 & n798 ;
  assign n6873 = ~n6871 & ~n6872 ;
  assign n6874 = n1806 & n4743 ;
  assign n6875 = n348 & n2901 ;
  assign n6876 = n829 & n6875 ;
  assign n6877 = ~n6874 & ~n6876 ;
  assign n6878 = ~n6873 & ~n6877 ;
  assign n6879 = ~n6870 & ~n6878 ;
  assign n6880 = ~n6834 & n6879 ;
  assign n6881 = n1478 & ~n6169 ;
  assign n6882 = n981 & n6436 ;
  assign n6883 = ~n6881 & ~n6882 ;
  assign n6884 = n373 & ~n6883 ;
  assign n6885 = n363 & n1762 ;
  assign n6886 = n846 & n6885 ;
  assign n6887 = ~n6884 & ~n6886 ;
  assign n6888 = ~x8 & ~n6887 ;
  assign n6889 = n1977 & n6871 ;
  assign n6890 = n5189 & n6889 ;
  assign n6891 = ~n6888 & ~n6890 ;
  assign n6892 = n2389 & ~n6891 ;
  assign n6893 = ~x9 & n2581 ;
  assign n6894 = n5838 & n6893 ;
  assign n6895 = n2481 & ~n6740 ;
  assign n6896 = ~n6894 & ~n6895 ;
  assign n6897 = n1874 & ~n6896 ;
  assign n6898 = x2 & n6897 ;
  assign n6899 = ~n6892 & ~n6898 ;
  assign n6900 = ~x5 & ~n6899 ;
  assign n6901 = n6880 & ~n6900 ;
  assign n6902 = ~n6821 & n6901 ;
  assign n6903 = ~n5852 & n6902 ;
  assign n6904 = x6 & ~n6903 ;
  assign n6905 = ~x1 & x6 ;
  assign n6906 = n1226 & n6905 ;
  assign n6907 = ~n1136 & n6906 ;
  assign n6908 = n496 & n6907 ;
  assign n6909 = n462 & n1656 ;
  assign n6910 = n524 & n1349 ;
  assign n6911 = n1742 & n5214 ;
  assign n6912 = ~n6910 & ~n6911 ;
  assign n6913 = ~n6909 & n6912 ;
  assign n6914 = x13 & n3530 ;
  assign n6915 = ~n6913 & n6914 ;
  assign n6916 = x6 & n1581 ;
  assign n6917 = n4271 & n6916 ;
  assign n6918 = ~x6 & n178 ;
  assign n6919 = ~x11 & n3030 ;
  assign n6920 = n6918 & n6919 ;
  assign n6921 = ~n6917 & ~n6920 ;
  assign n6922 = n866 & ~n6921 ;
  assign n6923 = ~x6 & ~x15 ;
  assign n6924 = ~x4 & n261 ;
  assign n6925 = n524 & n3021 ;
  assign n6926 = n6924 & n6925 ;
  assign n6927 = n6923 & n6926 ;
  assign n6928 = ~n6922 & ~n6927 ;
  assign n6929 = ~n6915 & n6928 ;
  assign n6930 = n276 & ~n6929 ;
  assign n6931 = ~n3293 & ~n3914 ;
  assign n6932 = n376 & n2286 ;
  assign n6933 = n6923 & n6932 ;
  assign n6934 = ~n6931 & n6933 ;
  assign n6935 = n2612 & n4309 ;
  assign n6936 = ~x11 & ~x15 ;
  assign n6937 = n381 & n3030 ;
  assign n6938 = ~n1136 & ~n3229 ;
  assign n6939 = ~n3098 & n6938 ;
  assign n6940 = ~n6937 & ~n6939 ;
  assign n6941 = n6940 ^ x1 ;
  assign n6942 = n6941 ^ n6940 ;
  assign n6943 = ~x0 & n2612 ;
  assign n6944 = n3030 & n6943 ;
  assign n6945 = n6944 ^ n6940 ;
  assign n6946 = n6942 & ~n6945 ;
  assign n6947 = n6946 ^ n6940 ;
  assign n6948 = n6936 & ~n6947 ;
  assign n6949 = ~n6935 & ~n6948 ;
  assign n6950 = n3075 & ~n6949 ;
  assign n6951 = ~n1169 & n4286 ;
  assign n6952 = ~x15 & ~n370 ;
  assign n6953 = n787 & ~n6952 ;
  assign n6954 = n6951 & n6953 ;
  assign n6955 = n877 & n2116 ;
  assign n6956 = n1010 & n1627 ;
  assign n6957 = n2747 & n6956 ;
  assign n6958 = n1954 & n2154 ;
  assign n6959 = ~n397 & n1683 ;
  assign n6960 = ~n6958 & ~n6959 ;
  assign n6961 = n845 & ~n6960 ;
  assign n6962 = ~n6957 & ~n6961 ;
  assign n6963 = ~n6955 & n6962 ;
  assign n6964 = ~n3960 & ~n6963 ;
  assign n6965 = ~n6954 & ~n6964 ;
  assign n6966 = n2608 & ~n6965 ;
  assign n6967 = ~n6950 & ~n6966 ;
  assign n6968 = ~n6934 & n6967 ;
  assign n6969 = n163 & ~n6968 ;
  assign n6970 = ~n6930 & ~n6969 ;
  assign n6971 = ~n6908 & n6970 ;
  assign n6972 = n2653 & ~n6971 ;
  assign n6973 = x11 & n371 ;
  assign n6974 = n348 & n2535 ;
  assign n6975 = n6973 & n6974 ;
  assign n6976 = n2831 & n4146 ;
  assign n6977 = ~n6975 & ~n6976 ;
  assign n6978 = ~n1136 & n2608 ;
  assign n6979 = n5703 & n6978 ;
  assign n6980 = ~n568 & n6979 ;
  assign n6981 = n6977 & ~n6980 ;
  assign n6982 = n1263 & ~n6981 ;
  assign n6983 = ~n4024 & ~n5153 ;
  assign n6984 = ~x4 & n4333 ;
  assign n6985 = ~n6983 & n6984 ;
  assign n6986 = x9 & n2358 ;
  assign n6987 = n376 & n6986 ;
  assign n6988 = n1905 & n6987 ;
  assign n6989 = ~n6985 & ~n6988 ;
  assign n6990 = n2806 & ~n6989 ;
  assign n6991 = ~x6 & x15 ;
  assign n6992 = ~x4 & n6991 ;
  assign n6993 = n396 & n846 ;
  assign n6994 = n6992 & n6993 ;
  assign n6995 = n827 & n2568 ;
  assign n6996 = n6994 & n6995 ;
  assign n6997 = n261 & n1494 ;
  assign n6998 = ~x15 & n2466 ;
  assign n6999 = ~x10 & n2686 ;
  assign n7000 = n6998 & n6999 ;
  assign n7001 = n6997 & n7000 ;
  assign n7002 = ~n6996 & ~n7001 ;
  assign n7003 = ~n6990 & n7002 ;
  assign n7004 = ~n869 & ~n7003 ;
  assign n7005 = ~n6982 & ~n7004 ;
  assign n7006 = ~x5 & ~n7005 ;
  assign n7007 = ~n5582 & n6159 ;
  assign n7008 = ~x9 & ~n7007 ;
  assign n7009 = ~n5173 & ~n7008 ;
  assign n7010 = n2831 & ~n7009 ;
  assign n7011 = ~x1 & n7010 ;
  assign n7291 = n261 & n2535 ;
  assign n7292 = n3462 & n7291 ;
  assign n7293 = n779 & n5386 ;
  assign n7294 = n195 & n7293 ;
  assign n7217 = ~x4 & ~x10 ;
  assign n7295 = ~n2466 & ~n7217 ;
  assign n7296 = n4545 & ~n7295 ;
  assign n7297 = n3229 & n3908 ;
  assign n7298 = n7296 & ~n7297 ;
  assign n7299 = ~x1 & n4155 ;
  assign n7300 = n3803 ^ n1499 ;
  assign n7301 = ~x14 & ~n7300 ;
  assign n7302 = n7301 ^ n1499 ;
  assign n7303 = n7299 & n7302 ;
  assign n7304 = ~n7298 & ~n7303 ;
  assign n7305 = x15 & ~n7304 ;
  assign n7306 = n391 & n1742 ;
  assign n7307 = n28 & n1282 ;
  assign n7308 = ~x12 & ~n7307 ;
  assign n7309 = x4 & ~n7308 ;
  assign n7139 = ~n1214 & ~n3030 ;
  assign n7310 = n513 & ~n7139 ;
  assign n7311 = ~n7309 & ~n7310 ;
  assign n7312 = n1104 & ~n7311 ;
  assign n7313 = ~n7306 & ~n7312 ;
  assign n7314 = ~n7305 & n7313 ;
  assign n7315 = ~n7294 & n7314 ;
  assign n7316 = x6 & ~n7315 ;
  assign n7317 = ~n7292 & ~n7316 ;
  assign n7012 = n4351 ^ n1742 ;
  assign n7013 = n7012 ^ n1742 ;
  assign n7014 = n1742 ^ x12 ;
  assign n7015 = n7014 ^ n1742 ;
  assign n7016 = n7013 & ~n7015 ;
  assign n7017 = n7016 ^ n1742 ;
  assign n7018 = x6 & n7017 ;
  assign n7019 = n7018 ^ n1742 ;
  assign n7020 = n2279 & n7019 ;
  assign n7021 = n762 & n7020 ;
  assign n7022 = ~x6 & x14 ;
  assign n7023 = n178 & n7022 ;
  assign n7024 = n2271 & n7023 ;
  assign n7025 = ~x10 & n7024 ;
  assign n7026 = n7025 ^ n7021 ;
  assign n7027 = ~x1 & n6923 ;
  assign n7028 = ~n1684 & n7027 ;
  assign n7029 = x0 & x6 ;
  assign n7030 = ~x15 & ~n7029 ;
  assign n7031 = ~x12 & ~n2815 ;
  assign n7032 = n568 & n7031 ;
  assign n7033 = ~n7030 & n7032 ;
  assign n7034 = ~n7028 & ~n7033 ;
  assign n7035 = n225 & ~n7034 ;
  assign n7036 = n568 & n1270 ;
  assign n7037 = n2538 & n7036 ;
  assign n7038 = ~n7035 & ~n7037 ;
  assign n7039 = n7038 ^ x11 ;
  assign n7040 = n7039 ^ n7038 ;
  assign n7041 = x1 & x6 ;
  assign n7042 = ~n5976 & ~n7041 ;
  assign n7043 = n1476 & ~n7042 ;
  assign n7044 = n2568 & n4339 ;
  assign n7045 = x14 & ~x15 ;
  assign n7046 = ~n7029 & n7045 ;
  assign n7047 = x1 & n7046 ;
  assign n7048 = ~n7044 & ~n7047 ;
  assign n7049 = ~x4 & ~n7048 ;
  assign n7050 = ~n7043 & ~n7049 ;
  assign n7051 = ~n1658 & ~n7050 ;
  assign n7052 = x4 & n7045 ;
  assign n7053 = n1628 & n7052 ;
  assign n7054 = ~n7051 & ~n7053 ;
  assign n7056 = ~x15 & n29 ;
  assign n7057 = n7042 & ~n7056 ;
  assign n7058 = n2799 & ~n7057 ;
  assign n7055 = n1382 & n2613 ;
  assign n7059 = n7058 ^ n7055 ;
  assign n7060 = n7059 ^ n7058 ;
  assign n7061 = n376 & n2607 ;
  assign n7062 = n4656 & n7061 ;
  assign n7063 = n7062 ^ n7058 ;
  assign n7064 = n7063 ^ n7058 ;
  assign n7065 = ~n7060 & ~n7064 ;
  assign n7066 = n7065 ^ n7058 ;
  assign n7067 = x0 & ~n7066 ;
  assign n7068 = n7067 ^ n7058 ;
  assign n7069 = n7054 & ~n7068 ;
  assign n7070 = n7069 ^ n7038 ;
  assign n7071 = ~n7040 & n7070 ;
  assign n7072 = n7071 ^ n7038 ;
  assign n7073 = n7072 ^ n7021 ;
  assign n7074 = n7026 & ~n7073 ;
  assign n7075 = n7074 ^ n7071 ;
  assign n7076 = n7075 ^ n7038 ;
  assign n7077 = n7076 ^ n7025 ;
  assign n7078 = ~n7021 & ~n7077 ;
  assign n7079 = n7078 ^ n7021 ;
  assign n7080 = n870 & n7079 ;
  assign n7081 = n306 & n2587 ;
  assign n7082 = ~n828 & ~n2290 ;
  assign n7083 = n7081 & n7082 ;
  assign n7084 = n1241 & n3098 ;
  assign n7085 = n489 & n7084 ;
  assign n7086 = n1905 & n7029 ;
  assign n7087 = x0 & n4201 ;
  assign n7088 = ~n780 & ~n7087 ;
  assign n7089 = n2668 & ~n7088 ;
  assign n7090 = ~n7086 & ~n7089 ;
  assign n7091 = ~n7085 & n7090 ;
  assign n7092 = n2329 & ~n7091 ;
  assign n7093 = ~n7083 & ~n7092 ;
  assign n7094 = ~x4 & ~n7093 ;
  assign n7095 = n1180 & n2522 ;
  assign n7096 = ~x10 & n7041 ;
  assign n7097 = n1227 & n7096 ;
  assign n7098 = ~n900 & ~n7097 ;
  assign n7099 = n2517 & ~n7098 ;
  assign n7100 = ~n7095 & ~n7099 ;
  assign n7101 = n57 & n60 ;
  assign n7102 = n2916 & n7101 ;
  assign n7103 = n381 & n2608 ;
  assign n7104 = x12 & n145 ;
  assign n7105 = ~n718 & ~n7104 ;
  assign n7106 = n462 & ~n7105 ;
  assign n7107 = n7103 & n7106 ;
  assign n7108 = ~n7102 & ~n7107 ;
  assign n7109 = n489 & n7027 ;
  assign n7110 = ~n1061 & ~n1241 ;
  assign n7111 = n2562 & ~n4339 ;
  assign n7112 = n274 & n7096 ;
  assign n7113 = x12 & n7112 ;
  assign n7114 = ~n7111 & ~n7113 ;
  assign n7115 = ~n7110 & ~n7114 ;
  assign n7116 = ~n7109 & ~n7115 ;
  assign n7117 = n718 & ~n7116 ;
  assign n7118 = n371 & n1282 ;
  assign n7119 = x6 ^ x1 ;
  assign n7120 = n7118 & ~n7119 ;
  assign n7121 = ~n7117 & ~n7120 ;
  assign n7122 = n1880 & ~n7121 ;
  assign n7123 = n7108 & ~n7122 ;
  assign n7124 = n7100 & n7123 ;
  assign n7125 = ~n7094 & n7124 ;
  assign n7126 = n7125 ^ x9 ;
  assign n7127 = n7126 ^ n7125 ;
  assign n7128 = n7127 ^ n7080 ;
  assign n7129 = ~n225 & ~n3288 ;
  assign n7130 = n828 & n4145 ;
  assign n7131 = n66 & n4155 ;
  assign n7132 = ~n7130 & ~n7131 ;
  assign n7133 = ~n7129 & ~n7132 ;
  assign n7134 = n178 & n4155 ;
  assign n7135 = n2568 & n7134 ;
  assign n7136 = ~n7133 & ~n7135 ;
  assign n7137 = x15 & ~n7136 ;
  assign n7138 = n1948 & n3039 ;
  assign n7140 = ~x10 & n7139 ;
  assign n7141 = ~x4 & n2413 ;
  assign n7142 = ~n7140 & n7141 ;
  assign n7143 = ~n7138 & ~n7142 ;
  assign n7144 = n306 & ~n7143 ;
  assign n7145 = ~n7137 & ~n7144 ;
  assign n7146 = n7145 ^ x6 ;
  assign n7147 = x6 & ~n7146 ;
  assign n7148 = n7147 ^ n7125 ;
  assign n7149 = n7148 ^ x6 ;
  assign n7150 = ~n7128 & ~n7149 ;
  assign n7151 = n7150 ^ n7147 ;
  assign n7152 = n7151 ^ x6 ;
  assign n7153 = ~n7080 & n7152 ;
  assign n7154 = n7153 ^ n7080 ;
  assign n7318 = n7317 ^ n7154 ;
  assign n7155 = n726 & n1601 ;
  assign n7156 = n2815 & n7155 ;
  assign n7157 = n1113 & ~n3960 ;
  assign n7158 = ~n5274 & ~n7157 ;
  assign n7159 = n1948 & ~n7158 ;
  assign n7160 = n7159 ^ x4 ;
  assign n7161 = n4318 ^ x0 ;
  assign n7162 = n7161 ^ n4318 ;
  assign n7163 = n718 & n4656 ;
  assign n7164 = n1214 & ~n3960 ;
  assign n7165 = ~n7163 & ~n7164 ;
  assign n7166 = n7165 ^ n4318 ;
  assign n7167 = ~n7162 & n7166 ;
  assign n7168 = n7167 ^ n4318 ;
  assign n7169 = n7168 ^ n7159 ;
  assign n7170 = n7160 & n7169 ;
  assign n7171 = n7170 ^ n7167 ;
  assign n7172 = n7171 ^ n4318 ;
  assign n7173 = n7172 ^ x4 ;
  assign n7174 = ~n7159 & n7173 ;
  assign n7175 = n7174 ^ n7159 ;
  assign n7176 = n7175 ^ n7159 ;
  assign n7177 = n453 & ~n7176 ;
  assign n7178 = ~x10 & ~n7139 ;
  assign n7179 = n1476 & n7178 ;
  assign n7180 = ~x14 & n863 ;
  assign n7181 = ~x12 & ~n7180 ;
  assign n7182 = ~x4 & ~n7181 ;
  assign n7183 = n866 & ~n7182 ;
  assign n7184 = n1476 & n4287 ;
  assign n7185 = n888 ^ x10 ;
  assign n7186 = n7185 ^ n888 ;
  assign n7187 = n888 ^ n76 ;
  assign n7188 = n7187 ^ n888 ;
  assign n7189 = n7186 & n7188 ;
  assign n7190 = n7189 ^ n888 ;
  assign n7191 = x4 & n7190 ;
  assign n7192 = n7191 ^ n888 ;
  assign n7193 = n1682 & n7192 ;
  assign n7194 = ~n7184 & ~n7193 ;
  assign n7195 = ~n7183 & n7194 ;
  assign n7198 = n7195 ^ x4 ;
  assign n7199 = n7198 ^ n7195 ;
  assign n7196 = n7195 ^ n489 ;
  assign n7197 = n7196 ^ n7195 ;
  assign n7200 = n7199 ^ n7197 ;
  assign n7201 = n3021 & n5698 ;
  assign n7202 = n7201 ^ n7195 ;
  assign n7203 = n7202 ^ n7195 ;
  assign n7204 = n7203 ^ n7199 ;
  assign n7205 = ~n7199 & ~n7204 ;
  assign n7206 = n7205 ^ n7199 ;
  assign n7207 = ~n7200 & ~n7206 ;
  assign n7208 = n7207 ^ n7205 ;
  assign n7209 = n7208 ^ n7195 ;
  assign n7210 = n7209 ^ n7199 ;
  assign n7211 = ~x1 & n7210 ;
  assign n7212 = n7211 ^ n7195 ;
  assign n7213 = ~n7179 & n7212 ;
  assign n7214 = ~n7177 & n7213 ;
  assign n7215 = x6 & ~n7214 ;
  assign n7216 = ~x11 & ~n7024 ;
  assign n7218 = n4035 & n7217 ;
  assign n7219 = ~n2600 & n7218 ;
  assign n7220 = ~x0 & n2668 ;
  assign n7221 = n719 & n7220 ;
  assign n7222 = x12 & ~x15 ;
  assign n7223 = n24 & n7222 ;
  assign n7224 = n3517 & n7223 ;
  assign n7225 = ~n7221 & ~n7224 ;
  assign n7226 = ~n7219 & n7225 ;
  assign n7227 = x1 & ~n7226 ;
  assign n7228 = n7216 & ~n7227 ;
  assign n7229 = ~n7215 & n7228 ;
  assign n7230 = ~n7163 & ~n7223 ;
  assign n7231 = n7230 ^ n6452 ;
  assign n7232 = x10 & ~n7231 ;
  assign n7233 = n7232 ^ n6452 ;
  assign n7234 = x0 & n7233 ;
  assign n7235 = ~x12 & n780 ;
  assign n7236 = ~n7234 & ~n7235 ;
  assign n7237 = n6918 & ~n7236 ;
  assign n7238 = x1 & ~x6 ;
  assign n7239 = ~n1227 & n2631 ;
  assign n7240 = ~n1214 & ~n5698 ;
  assign n7241 = ~n1136 & ~n7240 ;
  assign n7242 = ~n1270 & n7241 ;
  assign n7243 = ~n7239 & ~n7242 ;
  assign n7244 = n7238 & ~n7243 ;
  assign n7245 = n178 & ~n7180 ;
  assign n7246 = x1 & ~n1227 ;
  assign n7247 = ~n7245 & ~n7246 ;
  assign n7248 = n1678 & ~n7247 ;
  assign n7249 = ~x0 & n2522 ;
  assign n7250 = ~x1 & ~n1499 ;
  assign n7251 = ~n7249 & ~n7250 ;
  assign n7252 = ~n7248 & n7251 ;
  assign n7253 = n2587 & ~n7252 ;
  assign n7254 = x11 & ~n7253 ;
  assign n7255 = ~n7244 & n7254 ;
  assign n7256 = n376 & n7163 ;
  assign n7257 = n7240 ^ x12 ;
  assign n7258 = n7257 ^ n7240 ;
  assign n7259 = n7240 ^ n302 ;
  assign n7260 = n7259 ^ n7240 ;
  assign n7261 = ~n7258 & n7260 ;
  assign n7262 = n7261 ^ n7240 ;
  assign n7263 = ~x1 & ~n7262 ;
  assign n7264 = n7263 ^ n7240 ;
  assign n7265 = n60 & ~n7264 ;
  assign n7266 = ~n828 & ~n2522 ;
  assign n7267 = ~n19 & ~n7266 ;
  assign n7268 = ~x4 & n311 ;
  assign n7269 = n4346 & ~n7268 ;
  assign n7270 = n1327 & ~n7269 ;
  assign n7271 = n19 & n3960 ;
  assign n7272 = n2182 & n7271 ;
  assign n7273 = ~n7270 & ~n7272 ;
  assign n7274 = ~n7267 & n7273 ;
  assign n7275 = n7274 ^ x0 ;
  assign n7276 = n7275 ^ n7274 ;
  assign n7277 = x1 & n1214 ;
  assign n7278 = n3960 & n7277 ;
  assign n7279 = n7278 ^ n7274 ;
  assign n7280 = ~n7276 & ~n7279 ;
  assign n7281 = n7280 ^ n7274 ;
  assign n7282 = ~n7265 & n7281 ;
  assign n7283 = ~n7256 & n7282 ;
  assign n7284 = n2839 & ~n7283 ;
  assign n7285 = n7255 & ~n7284 ;
  assign n7286 = ~n7237 & n7285 ;
  assign n7287 = ~n7229 & ~n7286 ;
  assign n7288 = ~n7081 & ~n7287 ;
  assign n7289 = ~n7156 & n7288 ;
  assign n7290 = n7289 ^ n7154 ;
  assign n7319 = n7318 ^ n7290 ;
  assign n7320 = n7290 ^ x9 ;
  assign n7321 = n7320 ^ n7290 ;
  assign n7322 = n7319 & ~n7321 ;
  assign n7323 = n7322 ^ n7290 ;
  assign n7324 = x3 & ~n7323 ;
  assign n7325 = n7324 ^ n7154 ;
  assign n7326 = n7325 ^ x5 ;
  assign n7327 = n7326 ^ n7325 ;
  assign n7328 = n7327 ^ n7011 ;
  assign n7329 = n845 & n870 ;
  assign n7330 = ~n1627 & ~n4339 ;
  assign n7331 = n7329 & ~n7330 ;
  assign n7332 = ~n3229 & n7331 ;
  assign n7333 = ~x1 & n3960 ;
  assign n7334 = n828 & n7333 ;
  assign n7335 = ~n4280 & ~n7334 ;
  assign n7336 = ~n370 & ~n1198 ;
  assign n7337 = ~x14 & n414 ;
  assign n7338 = n7337 ^ x13 ;
  assign n7339 = n7338 ^ n7337 ;
  assign n7340 = n7339 ^ n7336 ;
  assign n7341 = ~n4351 & ~n6597 ;
  assign n7342 = n7341 ^ x12 ;
  assign n7343 = ~x12 & n7342 ;
  assign n7344 = n7343 ^ n7337 ;
  assign n7345 = n7344 ^ x12 ;
  assign n7346 = ~n7340 & ~n7345 ;
  assign n7347 = n7346 ^ n7343 ;
  assign n7348 = n7347 ^ x12 ;
  assign n7349 = ~n7336 & ~n7348 ;
  assign n7350 = n7349 ^ n7336 ;
  assign n7351 = n7335 & ~n7350 ;
  assign n7352 = x11 & n370 ;
  assign n7353 = n1349 & n4497 ;
  assign n7354 = ~n7352 & ~n7353 ;
  assign n7355 = x10 & ~n7354 ;
  assign n7356 = ~n7351 & ~n7355 ;
  assign n7357 = ~n7332 & n7356 ;
  assign n7358 = n3530 & ~n7357 ;
  assign n7359 = x14 & n1423 ;
  assign n7360 = ~n307 & ~n7359 ;
  assign n7361 = n2271 & n2398 ;
  assign n7363 = n105 & ~n1671 ;
  assign n7362 = x15 ^ x1 ;
  assign n7364 = n7363 ^ n7362 ;
  assign n7365 = n7364 ^ n7361 ;
  assign n7366 = n1114 ^ x1 ;
  assign n7367 = n7363 & n7366 ;
  assign n7368 = n7367 ^ n1114 ;
  assign n7369 = n7365 & n7368 ;
  assign n7370 = n7369 ^ n7367 ;
  assign n7371 = n7370 ^ n1114 ;
  assign n7372 = n7371 ^ n7363 ;
  assign n7373 = ~n7361 & n7372 ;
  assign n7374 = ~n7360 & n7373 ;
  assign n7375 = ~n306 & ~n4339 ;
  assign n7376 = ~n1270 & ~n5067 ;
  assign n7377 = ~n7375 & n7376 ;
  assign n7378 = n524 & n1214 ;
  assign n7379 = ~n306 & ~n7333 ;
  assign n7380 = n7378 & ~n7379 ;
  assign n7381 = ~n7377 & ~n7380 ;
  assign n7382 = ~n7374 & n7381 ;
  assign n7383 = n2826 & ~n7382 ;
  assign n7384 = ~x10 & ~n817 ;
  assign n7385 = ~n5410 & ~n7384 ;
  assign n7386 = n517 & ~n1270 ;
  assign n7387 = n346 & ~n3960 ;
  assign n7388 = n1113 & n7387 ;
  assign n7389 = ~n2741 & ~n7388 ;
  assign n7390 = ~n7386 & n7389 ;
  assign n7391 = ~x12 & ~n7390 ;
  assign n7392 = ~n7385 & ~n7391 ;
  assign n7393 = ~x1 & n2608 ;
  assign n7394 = ~n104 & n7393 ;
  assign n7395 = ~n7392 & n7394 ;
  assign n7396 = ~n7383 & ~n7395 ;
  assign n7397 = ~n7358 & n7396 ;
  assign n7398 = n7397 ^ x3 ;
  assign n7399 = ~n7397 & ~n7398 ;
  assign n7400 = n7399 ^ n7325 ;
  assign n7401 = n7400 ^ n7397 ;
  assign n7402 = ~n7328 & ~n7401 ;
  assign n7403 = n7402 ^ n7399 ;
  assign n7404 = n7403 ^ n7397 ;
  assign n7405 = ~n7011 & ~n7404 ;
  assign n7406 = n7405 ^ n7011 ;
  assign n7407 = n7406 ^ x7 ;
  assign n7408 = n7407 ^ n7406 ;
  assign n7409 = n2587 & n5507 ;
  assign n7410 = n1246 & n7409 ;
  assign n7411 = x15 ^ x14 ;
  assign n7412 = ~x1 & ~x6 ;
  assign n7413 = n7412 ^ x15 ;
  assign n7414 = n7411 & ~n7413 ;
  assign n7415 = n7414 ^ x15 ;
  assign n7416 = n828 & n7415 ;
  assign n7417 = n2668 ^ n57 ;
  assign n7418 = n7417 ^ n57 ;
  assign n7419 = n7418 ^ n7416 ;
  assign n7420 = ~n2811 & ~n4829 ;
  assign n7421 = n7420 ^ n6905 ;
  assign n7422 = n7420 & ~n7421 ;
  assign n7423 = n7422 ^ n57 ;
  assign n7424 = n7423 ^ n7420 ;
  assign n7425 = n7419 & n7424 ;
  assign n7426 = n7425 ^ n7422 ;
  assign n7427 = n7426 ^ n7420 ;
  assign n7428 = ~n7416 & n7427 ;
  assign n7429 = n7428 ^ n7416 ;
  assign n7430 = n978 & n7429 ;
  assign n7431 = ~x12 & n2850 ;
  assign n7432 = ~n1246 & ~n1283 ;
  assign n7433 = ~n2509 & n7432 ;
  assign n7434 = ~n7431 & n7433 ;
  assign n7435 = ~x1 & ~n7434 ;
  assign n7436 = ~n248 & ~n1327 ;
  assign n7437 = ~x15 & ~n7436 ;
  assign n7438 = ~n6620 & ~n7337 ;
  assign n7439 = ~x0 & n1214 ;
  assign n7440 = ~n60 & ~n7439 ;
  assign n7441 = n7438 & ~n7440 ;
  assign n7442 = ~n7437 & n7441 ;
  assign n7443 = n240 & ~n1627 ;
  assign n7444 = ~n1283 & ~n7443 ;
  assign n7445 = ~n7333 & n7444 ;
  assign n7446 = ~x6 & ~n7445 ;
  assign n7447 = n7442 & ~n7446 ;
  assign n7448 = ~n7435 & n7447 ;
  assign n7449 = x14 & n7412 ;
  assign n7450 = ~n986 & n7449 ;
  assign n7451 = ~n7246 & ~n7450 ;
  assign n7452 = n2810 & ~n7451 ;
  assign n7453 = ~n414 & ~n642 ;
  assign n7454 = x6 & n4196 ;
  assign n7455 = ~n7453 & n7454 ;
  assign n7456 = n7271 ^ x6 ;
  assign n7457 = n7456 ^ n7271 ;
  assign n7458 = n7457 ^ n2605 ;
  assign n7459 = x13 ^ x1 ;
  assign n7460 = ~x1 & n7459 ;
  assign n7461 = n7460 ^ n7271 ;
  assign n7462 = n7461 ^ x1 ;
  assign n7463 = n7458 & n7462 ;
  assign n7464 = n7463 ^ n7460 ;
  assign n7465 = n7464 ^ x1 ;
  assign n7466 = n2605 & ~n7465 ;
  assign n7467 = n7466 ^ n2605 ;
  assign n7468 = ~n7455 & ~n7467 ;
  assign n7469 = ~n7452 & n7468 ;
  assign n7470 = ~n7448 & n7469 ;
  assign n7471 = ~n7430 & n7470 ;
  assign n7472 = n1679 & ~n7471 ;
  assign n7473 = ~n3098 & ~n7022 ;
  assign n7474 = ~n7132 & ~n7473 ;
  assign n7475 = n4155 & n4829 ;
  assign n7476 = n2562 & n7475 ;
  assign n7477 = ~n7474 & ~n7476 ;
  assign n7478 = x15 & ~n7477 ;
  assign n7479 = n6158 & n7096 ;
  assign n7480 = ~n453 & n2312 ;
  assign n7481 = ~n718 & n7139 ;
  assign n7482 = n5526 & ~n7481 ;
  assign n7483 = ~n2398 & ~n7482 ;
  assign n7484 = ~n7480 & n7483 ;
  assign n7485 = n2562 & ~n7484 ;
  assign n7486 = ~n7479 & ~n7485 ;
  assign n7487 = ~n7478 & n7486 ;
  assign n7488 = ~x3 & ~n7487 ;
  assign n7489 = ~n2290 & ~n4351 ;
  assign n7490 = ~n392 & n7489 ;
  assign n7491 = ~x0 & ~n6118 ;
  assign n7492 = ~n7490 & n7491 ;
  assign n7493 = n2815 ^ n748 ;
  assign n7494 = n7493 ^ n748 ;
  assign n7495 = ~n1555 & ~n2116 ;
  assign n7496 = ~n7271 & ~n7495 ;
  assign n7497 = n7496 ^ n748 ;
  assign n7498 = n7494 & ~n7497 ;
  assign n7499 = n7498 ^ n748 ;
  assign n7500 = n405 & ~n7499 ;
  assign n7501 = ~n7492 & n7500 ;
  assign n7502 = x9 & ~n6907 ;
  assign n7503 = ~n7501 & n7502 ;
  assign n7504 = ~n7488 & n7503 ;
  assign n7505 = ~n7472 & n7504 ;
  assign n7506 = n240 & ~n3080 ;
  assign n7507 = n4428 & n7506 ;
  assign n7508 = n57 & n2668 ;
  assign n7509 = n5625 & n7508 ;
  assign n7510 = ~n7507 & ~n7509 ;
  assign n7511 = ~n2600 & n4155 ;
  assign n7512 = n2948 & n6943 ;
  assign n7513 = ~n7511 & ~n7512 ;
  assign n7514 = n4333 & ~n7513 ;
  assign n7515 = n7510 & ~n7514 ;
  assign n7516 = n1270 & ~n7515 ;
  assign n7517 = n2562 & n4735 ;
  assign n7518 = ~x14 & ~n7082 ;
  assign n7519 = n7517 & ~n7518 ;
  assign n7520 = n4656 & n6943 ;
  assign n7521 = n759 & n4333 ;
  assign n7522 = n7520 & n7521 ;
  assign n7523 = ~x9 & ~n7522 ;
  assign n7524 = ~n7519 & n7523 ;
  assign n7538 = ~x15 & n673 ;
  assign n7539 = ~x12 & ~n7538 ;
  assign n7540 = x6 & ~n7539 ;
  assign n7541 = ~n7506 & ~n7540 ;
  assign n7542 = x1 & ~n7541 ;
  assign n7543 = n828 & n6905 ;
  assign n7544 = ~n1349 & n4685 ;
  assign n7545 = ~x6 & n7544 ;
  assign n7546 = ~n7543 & ~n7545 ;
  assign n7547 = x14 & ~n7546 ;
  assign n7548 = ~n7542 & ~n7547 ;
  assign n7549 = n489 & ~n7548 ;
  assign n7525 = n7308 ^ x1 ;
  assign n7526 = n7525 ^ n7308 ;
  assign n7527 = n7308 ^ n7139 ;
  assign n7528 = n7527 ^ n7308 ;
  assign n7529 = n7526 & ~n7528 ;
  assign n7530 = n7529 ^ n7308 ;
  assign n7531 = ~x6 & ~n7530 ;
  assign n7532 = n7531 ^ n7308 ;
  assign n7533 = n1104 & ~n7532 ;
  assign n7534 = n2562 & n7293 ;
  assign n7535 = n1743 & n2587 ;
  assign n7536 = ~n7534 & ~n7535 ;
  assign n7537 = ~n7533 & n7536 ;
  assign n7550 = n7549 ^ n7537 ;
  assign n7551 = n7550 ^ n7537 ;
  assign n7552 = ~n727 & n1656 ;
  assign n7553 = ~n122 & n7552 ;
  assign n7554 = ~n45 & ~n105 ;
  assign n7555 = n1905 & ~n2271 ;
  assign n7556 = n7554 & n7555 ;
  assign n7557 = ~x0 & n2312 ;
  assign n7558 = ~n7556 & ~n7557 ;
  assign n7559 = ~n7553 & n7558 ;
  assign n7560 = n7041 & ~n7559 ;
  assign n7561 = n7560 ^ n7537 ;
  assign n7562 = n7561 ^ n7537 ;
  assign n7563 = ~n7551 & ~n7562 ;
  assign n7564 = n7563 ^ n7537 ;
  assign n7565 = ~x3 & n7564 ;
  assign n7566 = n7565 ^ n7537 ;
  assign n7567 = n7524 & n7566 ;
  assign n7568 = ~n7516 & n7567 ;
  assign n7569 = ~n7505 & ~n7568 ;
  assign n7570 = ~n7410 & ~n7569 ;
  assign n7571 = n795 & ~n7570 ;
  assign n7572 = ~n1658 & ~n5650 ;
  assign n7573 = ~n4295 & ~n7572 ;
  assign n7574 = n26 & ~n7573 ;
  assign n7575 = ~x10 & ~n7163 ;
  assign n7576 = n843 & ~n7575 ;
  assign n7577 = n2693 & n4035 ;
  assign n7578 = n2612 & n7181 ;
  assign n7579 = ~n1601 & ~n7578 ;
  assign n7580 = ~n7577 & n7579 ;
  assign n7581 = n739 & ~n7580 ;
  assign n7582 = ~n7576 & ~n7581 ;
  assign n7583 = ~n7574 & n7582 ;
  assign n7584 = n517 & ~n7583 ;
  assign n7585 = ~x6 & n739 ;
  assign n7586 = n5699 & n7585 ;
  assign n7587 = ~n3229 & n7586 ;
  assign n7588 = ~n7584 & ~n7587 ;
  assign n7589 = n224 & ~n7588 ;
  assign n7590 = n739 & n2803 ;
  assign n7591 = n3835 & n7590 ;
  assign n7592 = n1353 & n1423 ;
  assign n7593 = n7591 & n7592 ;
  assign n7594 = x12 & n104 ;
  assign n7595 = ~n240 & ~n1353 ;
  assign n7596 = n7595 ^ x11 ;
  assign n7597 = n7596 ^ n7595 ;
  assign n7598 = n7595 ^ n1227 ;
  assign n7599 = n7598 ^ n7595 ;
  assign n7600 = n7597 & n7599 ;
  assign n7601 = n7600 ^ n7595 ;
  assign n7602 = ~x5 & ~n7601 ;
  assign n7603 = n7602 ^ n7595 ;
  assign n7604 = n7594 & ~n7603 ;
  assign n7605 = n4015 & n4155 ;
  assign n7606 = n7605 ^ x5 ;
  assign n7607 = n7606 ^ n7605 ;
  assign n7608 = ~x13 & n845 ;
  assign n7609 = n7222 & n7608 ;
  assign n7610 = ~n427 & n828 ;
  assign n7611 = x10 & x15 ;
  assign n7612 = ~n1010 & ~n7611 ;
  assign n7613 = n7610 & ~n7612 ;
  assign n7614 = ~n474 & ~n7613 ;
  assign n7615 = ~n7609 & n7614 ;
  assign n7616 = n7615 ^ n7605 ;
  assign n7617 = n7616 ^ n7605 ;
  assign n7618 = n7607 & ~n7617 ;
  assign n7619 = n7618 ^ n7605 ;
  assign n7620 = ~x9 & n7619 ;
  assign n7621 = n7620 ^ n7605 ;
  assign n7622 = ~n5947 & ~n7621 ;
  assign n7623 = x14 & ~n7622 ;
  assign n7624 = ~n7604 & ~n7623 ;
  assign n7625 = x0 & n3002 ;
  assign n7626 = ~n7624 & n7625 ;
  assign n7627 = ~n624 & n7577 ;
  assign n7628 = ~n1270 & ~n1905 ;
  assign n7629 = n3894 & ~n7628 ;
  assign n7630 = ~n890 & n7629 ;
  assign n7631 = ~x6 & x13 ;
  assign n7632 = x10 & n3960 ;
  assign n7633 = ~n7631 & ~n7632 ;
  assign n7634 = x5 & ~n473 ;
  assign n7635 = ~n7633 & n7634 ;
  assign n7636 = ~n7630 & ~n7635 ;
  assign n7637 = x12 & ~n7636 ;
  assign n7638 = ~n7627 & ~n7637 ;
  assign n7639 = x3 & n817 ;
  assign n7640 = n1880 & n7639 ;
  assign n7641 = ~n7638 & n7640 ;
  assign n7642 = ~n7626 & ~n7641 ;
  assign n7643 = ~n7593 & n7642 ;
  assign n7644 = ~n7589 & n7643 ;
  assign n7645 = x1 & ~n7644 ;
  assign n7646 = n75 & n366 ;
  assign n7647 = n195 & ~n2370 ;
  assign n7648 = ~n7646 & ~n7647 ;
  assign n7649 = x1 & ~n7648 ;
  assign n7650 = ~n1995 & ~n7649 ;
  assign n7651 = n346 & ~n7650 ;
  assign n7652 = n373 & n739 ;
  assign n7653 = n2389 & n7652 ;
  assign n7654 = ~n7651 & ~n7653 ;
  assign n7655 = n1214 & ~n7654 ;
  assign n7656 = n1948 & n2387 ;
  assign n7657 = n1114 & n7656 ;
  assign n7658 = ~n7655 & ~n7657 ;
  assign n7659 = n6991 & ~n7658 ;
  assign n7660 = n1283 & n3126 ;
  assign n7661 = n6997 & n7660 ;
  assign n7662 = ~n7659 & ~n7661 ;
  assign n7663 = ~n3012 & ~n7662 ;
  assign n7664 = x3 & n2755 ;
  assign n7665 = x11 & n306 ;
  assign n7666 = ~n7575 & n7665 ;
  assign n7667 = n122 & n7233 ;
  assign n7668 = ~n6163 & ~n7667 ;
  assign n7669 = n7668 ^ x1 ;
  assign n7670 = n7669 ^ n7668 ;
  assign n7671 = n7670 ^ n7666 ;
  assign n7672 = n3030 ^ n471 ;
  assign n7673 = n471 & n7672 ;
  assign n7674 = n7673 ^ n7668 ;
  assign n7675 = n7674 ^ n471 ;
  assign n7676 = n7671 & ~n7675 ;
  assign n7677 = n7676 ^ n7673 ;
  assign n7678 = n7677 ^ n471 ;
  assign n7679 = ~n7666 & n7678 ;
  assign n7680 = n7679 ^ n7666 ;
  assign n7681 = n7664 & n7680 ;
  assign n7682 = n1538 & n7681 ;
  assign n7683 = ~n7663 & ~n7682 ;
  assign n7684 = ~n7645 & n7683 ;
  assign n7685 = n5044 & n7045 ;
  assign n7686 = n2300 & n7685 ;
  assign n7687 = ~n1214 & ~n1226 ;
  assign n7688 = n89 & n5521 ;
  assign n7689 = n7687 & n7688 ;
  assign n7690 = ~n7686 & ~n7689 ;
  assign n7691 = ~x9 & ~n7690 ;
  assign n7692 = ~x13 & n7045 ;
  assign n7693 = ~n2036 & ~n7692 ;
  assign n7694 = n978 & n1920 ;
  assign n7695 = ~n7693 & n7694 ;
  assign n7696 = ~n7691 & ~n7695 ;
  assign n7697 = ~n1692 & ~n3728 ;
  assign n7698 = x12 & n414 ;
  assign n7699 = ~n4170 & n7698 ;
  assign n7700 = ~n7697 & n7699 ;
  assign n7701 = ~n319 & n7387 ;
  assign n7702 = ~n75 & ~n571 ;
  assign n7703 = n7701 & ~n7702 ;
  assign n7704 = ~n7700 & ~n7703 ;
  assign n7705 = x13 & ~n7704 ;
  assign n7706 = ~x15 & n1920 ;
  assign n7707 = ~n1630 & ~n7706 ;
  assign n7708 = n2282 & ~n7707 ;
  assign n7709 = n105 & n7708 ;
  assign n7710 = ~n7705 & ~n7709 ;
  assign n7711 = n7696 & n7710 ;
  assign n7712 = n2279 & ~n7711 ;
  assign n7713 = ~n427 & n624 ;
  assign n7714 = x12 & n7713 ;
  assign n7715 = ~n1010 & n7714 ;
  assign n7716 = ~n105 & ~n557 ;
  assign n7717 = n6037 & ~n7716 ;
  assign n7718 = x5 & ~x15 ;
  assign n7719 = ~n2119 & n7718 ;
  assign n7720 = ~n7717 & ~n7719 ;
  assign n7721 = ~n7715 & n7720 ;
  assign n7722 = n2282 & ~n7721 ;
  assign n7723 = n1435 & n7685 ;
  assign n7724 = n571 & n1353 ;
  assign n7725 = n1246 & n7724 ;
  assign n7726 = ~n7723 & ~n7725 ;
  assign n7727 = ~n7722 & n7726 ;
  assign n7728 = n3075 & ~n7727 ;
  assign n7729 = n1785 ^ n381 ;
  assign n7730 = n371 ^ x12 ;
  assign n7731 = n1353 ^ x12 ;
  assign n7732 = n7730 & n7731 ;
  assign n7733 = n7732 ^ x12 ;
  assign n7734 = n7733 ^ n1785 ;
  assign n7735 = ~n7729 & n7734 ;
  assign n7736 = n7735 ^ n7732 ;
  assign n7737 = n7736 ^ x12 ;
  assign n7738 = n7737 ^ n381 ;
  assign n7739 = n1785 & ~n7738 ;
  assign n7740 = n7739 ^ n1785 ;
  assign n7741 = ~n7728 & ~n7740 ;
  assign n7742 = ~n7712 & n7741 ;
  assign n7745 = n7742 ^ x5 ;
  assign n7746 = n7745 ^ n7742 ;
  assign n7743 = n7742 ^ n346 ;
  assign n7744 = n7743 ^ n7742 ;
  assign n7747 = n7746 ^ n7744 ;
  assign n7748 = ~x0 & n1656 ;
  assign n7749 = n1353 & n7748 ;
  assign n7750 = n1136 & ~n7749 ;
  assign n7751 = n4005 & ~n7750 ;
  assign n7752 = n7751 ^ n7742 ;
  assign n7753 = n7752 ^ n7742 ;
  assign n7754 = n7753 ^ n7746 ;
  assign n7755 = n7746 & n7754 ;
  assign n7756 = n7755 ^ n7746 ;
  assign n7757 = n7747 & n7756 ;
  assign n7758 = n7757 ^ n7755 ;
  assign n7759 = n7758 ^ n7742 ;
  assign n7760 = n7759 ^ n7746 ;
  assign n7761 = x6 & ~n7760 ;
  assign n7762 = n7761 ^ n7742 ;
  assign n7763 = n442 & ~n7762 ;
  assign n7764 = ~n1353 & n1678 ;
  assign n7765 = ~n787 & n4647 ;
  assign n7766 = ~n7764 & n7765 ;
  assign n7767 = n307 & n404 ;
  assign n7768 = ~x15 & n4206 ;
  assign n7769 = n4422 & n7768 ;
  assign n7770 = ~n7767 & ~n7769 ;
  assign n7771 = ~x3 & ~n7770 ;
  assign n7772 = n76 & ~n1169 ;
  assign n7773 = n224 & n7772 ;
  assign n7774 = ~n7771 & ~n7773 ;
  assign n7775 = n5410 & ~n7774 ;
  assign n7776 = ~n270 & ~n7639 ;
  assign n7777 = n4909 & ~n7776 ;
  assign n7778 = ~n306 & n7777 ;
  assign n7779 = n373 & n5332 ;
  assign n7780 = n1678 & n6095 ;
  assign n7781 = x0 & n395 ;
  assign n7782 = n6359 & n7781 ;
  assign n7783 = n727 & n1263 ;
  assign n7784 = ~n1743 & ~n7783 ;
  assign n7785 = ~n7782 & n7784 ;
  assign n7786 = ~n7780 & n7785 ;
  assign n7787 = n383 & ~n7786 ;
  assign n7788 = ~n7779 & ~n7787 ;
  assign n7789 = ~n7778 & n7788 ;
  assign n7790 = n7789 ^ x10 ;
  assign n7791 = n7790 ^ n7789 ;
  assign n7792 = n7791 ^ n7775 ;
  assign n7793 = n5516 & n7693 ;
  assign n7794 = n1169 & ~n7793 ;
  assign n7795 = ~n404 & ~n1282 ;
  assign n7796 = x1 & ~n7795 ;
  assign n7797 = ~n1364 & n7796 ;
  assign n7798 = ~n7794 & ~n7797 ;
  assign n7799 = n25 & ~n7798 ;
  assign n7800 = n870 & n6097 ;
  assign n7801 = ~n1565 & ~n5819 ;
  assign n7802 = x0 & ~n4881 ;
  assign n7803 = ~n7801 & n7802 ;
  assign n7804 = ~n7800 & ~n7803 ;
  assign n7805 = n1627 & ~n7804 ;
  assign n7806 = n28 & n2154 ;
  assign n7807 = n1227 & n4751 ;
  assign n7808 = n1382 & n3960 ;
  assign n7809 = x9 & n7808 ;
  assign n7810 = ~n7807 & ~n7809 ;
  assign n7811 = ~n7806 & n7810 ;
  assign n7812 = n373 & ~n7811 ;
  assign n7813 = n6295 & n7639 ;
  assign n7814 = n530 & n4421 ;
  assign n7815 = ~n7813 & ~n7814 ;
  assign n7816 = ~n6993 & n7815 ;
  assign n7817 = ~n7812 & n7816 ;
  assign n7818 = ~n7805 & n7817 ;
  assign n7819 = ~n7799 & n7818 ;
  assign n7820 = n7819 ^ x11 ;
  assign n7821 = ~n7819 & n7820 ;
  assign n7822 = n7821 ^ n7789 ;
  assign n7823 = n7822 ^ n7819 ;
  assign n7824 = n7792 & n7823 ;
  assign n7825 = n7824 ^ n7821 ;
  assign n7826 = n7825 ^ n7819 ;
  assign n7827 = ~n7775 & ~n7826 ;
  assign n7828 = n7827 ^ n7775 ;
  assign n7829 = ~n7766 & ~n7828 ;
  assign n7830 = n2870 & ~n7829 ;
  assign n7831 = ~n7763 & ~n7830 ;
  assign n7832 = n2781 & n5838 ;
  assign n7833 = ~n329 & n2755 ;
  assign n7834 = x15 & n888 ;
  assign n7835 = ~n452 & ~n7834 ;
  assign n7836 = ~n34 & n3030 ;
  assign n7837 = ~n7835 & n7836 ;
  assign n7838 = n7833 & n7837 ;
  assign n7839 = n1565 & n2188 ;
  assign n7840 = x0 & ~n3130 ;
  assign n7841 = n311 & n517 ;
  assign n7842 = ~n46 & n7841 ;
  assign n7843 = ~n7840 & n7842 ;
  assign n7844 = n7843 ^ x12 ;
  assign n7845 = n7844 ^ n7843 ;
  assign n7846 = n7845 ^ n2612 ;
  assign n7847 = x15 ^ x13 ;
  assign n7848 = n526 ^ x15 ;
  assign n7849 = n7848 ^ n526 ;
  assign n7850 = n1923 & n7849 ;
  assign n7851 = n7850 ^ n526 ;
  assign n7852 = ~n7847 & n7851 ;
  assign n7853 = n2568 & n7852 ;
  assign n7854 = ~n145 & ~n530 ;
  assign n7855 = ~n86 & ~n526 ;
  assign n7856 = ~n7854 & ~n7855 ;
  assign n7857 = ~n7853 & ~n7856 ;
  assign n7858 = x11 & ~n7857 ;
  assign n7859 = n1114 & ~n7697 ;
  assign n7860 = n7859 ^ n7858 ;
  assign n7861 = ~n7858 & n7860 ;
  assign n7862 = n7861 ^ n7843 ;
  assign n7863 = n7862 ^ n7858 ;
  assign n7864 = n7846 & n7863 ;
  assign n7865 = n7864 ^ n7861 ;
  assign n7866 = n7865 ^ n7858 ;
  assign n7867 = n2612 & ~n7866 ;
  assign n7868 = n7867 ^ n2612 ;
  assign n7869 = ~n7839 & ~n7868 ;
  assign n7870 = ~n7838 & n7869 ;
  assign n7871 = ~x4 & ~n7870 ;
  assign n7872 = ~n7832 & ~n7871 ;
  assign n7873 = n38 & ~n7872 ;
  assign n7874 = x14 ^ x12 ;
  assign n7875 = ~x13 & n2587 ;
  assign n7876 = ~n1679 & n2537 ;
  assign n7877 = ~n1657 & ~n7876 ;
  assign n7878 = ~n7875 & ~n7877 ;
  assign n7879 = n863 & n1785 ;
  assign n7882 = n7879 ^ n2575 ;
  assign n7883 = n7882 ^ n7879 ;
  assign n7880 = n7879 ^ n1903 ;
  assign n7881 = n7880 ^ n7879 ;
  assign n7884 = n7883 ^ n7881 ;
  assign n7885 = n7879 ^ x15 ;
  assign n7886 = n7885 ^ n7879 ;
  assign n7887 = n7886 ^ n7883 ;
  assign n7888 = ~n7883 & ~n7887 ;
  assign n7889 = n7888 ^ n7883 ;
  assign n7890 = ~n7884 & ~n7889 ;
  assign n7891 = n7890 ^ n7888 ;
  assign n7892 = n7891 ^ n7879 ;
  assign n7893 = n7892 ^ n7883 ;
  assign n7894 = x3 & ~n7893 ;
  assign n7895 = n7894 ^ n7879 ;
  assign n7896 = n7878 & n7895 ;
  assign n7897 = x15 & n168 ;
  assign n7898 = n2741 & n7897 ;
  assign n7899 = ~x5 & n6923 ;
  assign n7900 = n276 & n392 ;
  assign n7901 = n7899 & n7900 ;
  assign n7902 = ~n7898 & ~n7901 ;
  assign n7903 = n2279 & ~n7902 ;
  assign n7904 = ~n7896 & ~n7903 ;
  assign n7905 = n7904 ^ n7874 ;
  assign n7906 = n7905 ^ x14 ;
  assign n7907 = n7906 ^ n7905 ;
  assign n7908 = x9 & n383 ;
  assign n7909 = ~n1991 & n7908 ;
  assign n7910 = n7909 ^ n26 ;
  assign n7911 = n7909 ^ n3761 ;
  assign n7912 = n7911 ^ n3761 ;
  assign n7913 = n7912 ^ n7910 ;
  assign n7914 = n346 & n2811 ;
  assign n7915 = n7914 ^ x3 ;
  assign n7916 = n7914 & ~n7915 ;
  assign n7917 = n7916 ^ n3761 ;
  assign n7918 = n7917 ^ n7914 ;
  assign n7919 = ~n7913 & ~n7918 ;
  assign n7920 = n7919 ^ n7916 ;
  assign n7921 = n7920 ^ n7914 ;
  assign n7922 = n7910 & n7921 ;
  assign n7923 = n7922 ^ n7909 ;
  assign n7924 = n7632 & n7923 ;
  assign n7925 = n7608 & n7718 ;
  assign n7926 = ~n145 & ~n863 ;
  assign n7927 = ~n511 & n739 ;
  assign n7928 = ~n7926 & n7927 ;
  assign n7929 = n7928 ^ x11 ;
  assign n7930 = n7929 ^ n7928 ;
  assign n7931 = n7930 ^ n7925 ;
  assign n7932 = n411 ^ x4 ;
  assign n7933 = ~x4 & ~n7932 ;
  assign n7934 = n7933 ^ n7928 ;
  assign n7935 = n7934 ^ x4 ;
  assign n7936 = n7931 & ~n7935 ;
  assign n7937 = n7936 ^ n7933 ;
  assign n7938 = n7937 ^ x4 ;
  assign n7939 = ~n7925 & ~n7938 ;
  assign n7940 = n7939 ^ n7925 ;
  assign n7941 = n1559 & n7940 ;
  assign n7942 = ~x6 & n7941 ;
  assign n7943 = ~n7924 & ~n7942 ;
  assign n7944 = n7943 ^ n7905 ;
  assign n7945 = n7944 ^ n7874 ;
  assign n7946 = n7907 & ~n7945 ;
  assign n7947 = n7946 ^ n7943 ;
  assign n7948 = ~x4 & x13 ;
  assign n7949 = n4649 ^ x15 ;
  assign n7950 = n7949 ^ n4649 ;
  assign n7951 = n4649 ^ n2693 ;
  assign n7952 = n7951 ^ n4649 ;
  assign n7953 = n7950 & n7952 ;
  assign n7954 = n7953 ^ n4649 ;
  assign n7955 = ~x5 & ~n7954 ;
  assign n7956 = n7955 ^ n4649 ;
  assign n7957 = n7948 & ~n7956 ;
  assign n7958 = ~n644 & n843 ;
  assign n7959 = ~x10 & n7958 ;
  assign n7960 = ~n7957 & ~n7959 ;
  assign n7961 = n375 & ~n7960 ;
  assign n7962 = n7943 & ~n7961 ;
  assign n7963 = n7962 ^ n7874 ;
  assign n7964 = n7947 & ~n7963 ;
  assign n7965 = n7964 ^ n7962 ;
  assign n7966 = ~n7874 & n7965 ;
  assign n7967 = n7966 ^ n7946 ;
  assign n7968 = n7967 ^ x12 ;
  assign n7969 = n7968 ^ n7943 ;
  assign n7970 = n1954 & n7969 ;
  assign n7971 = ~n7873 & ~n7970 ;
  assign n7972 = n7831 & n7971 ;
  assign n7973 = n7684 & n7972 ;
  assign n7974 = ~n7571 & n7973 ;
  assign n7975 = n7974 ^ n7406 ;
  assign n7976 = ~n7408 & ~n7975 ;
  assign n7977 = n7976 ^ n7406 ;
  assign n7978 = ~n7006 & ~n7977 ;
  assign n7979 = ~n6972 & n7978 ;
  assign n7980 = ~n850 & ~n7979 ;
  assign n7981 = n2810 & n3192 ;
  assign n7982 = n105 & ~n319 ;
  assign n7983 = ~n1050 & ~n7982 ;
  assign n7984 = n1683 & ~n2848 ;
  assign n7985 = n1905 & n7984 ;
  assign n7986 = n7983 & n7985 ;
  assign n7987 = ~n7981 & ~n7986 ;
  assign n7993 = n673 & n4167 ;
  assign n7994 = n2180 & n7993 ;
  assign n7995 = n762 & ~n6709 ;
  assign n7996 = ~n7994 & ~n7995 ;
  assign n7988 = n4392 & n4656 ;
  assign n7989 = ~n3972 & ~n7988 ;
  assign n7990 = n60 & ~n7989 ;
  assign n7991 = n4033 & n4069 ;
  assign n7992 = ~n7990 & ~n7991 ;
  assign n7997 = n7996 ^ n7992 ;
  assign n7998 = n7997 ^ n7992 ;
  assign n7999 = n787 & n7201 ;
  assign n8000 = ~n1240 & ~n7999 ;
  assign n8001 = n2653 & ~n8000 ;
  assign n8002 = n8001 ^ n7992 ;
  assign n8003 = n8002 ^ n7992 ;
  assign n8004 = n7998 & ~n8003 ;
  assign n8005 = n8004 ^ n7992 ;
  assign n8006 = x10 & n8005 ;
  assign n8007 = n8006 ^ n7992 ;
  assign n8008 = n7987 & n8007 ;
  assign n8009 = n778 & ~n8008 ;
  assign n8010 = ~n768 & n6514 ;
  assign n8011 = n465 & ~n1226 ;
  assign n8012 = n8010 & n8011 ;
  assign n8013 = n928 & n3681 ;
  assign n8014 = ~n8012 & ~n8013 ;
  assign n8015 = ~n8009 & n8014 ;
  assign n8016 = n7393 & ~n8015 ;
  assign n8017 = n739 & n2806 ;
  assign n8018 = n795 & n1422 ;
  assign n8019 = ~n8017 & ~n8018 ;
  assign n8020 = n306 & ~n8019 ;
  assign n8021 = n66 & n2806 ;
  assign n8022 = n795 & n8021 ;
  assign n8023 = ~n8020 & ~n8022 ;
  assign n8024 = n4644 & ~n8023 ;
  assign n8025 = n778 & n4829 ;
  assign n8026 = n1002 & n8025 ;
  assign n8027 = n3425 & n8026 ;
  assign n8028 = ~n4422 & n4513 ;
  assign n8029 = n988 & n4829 ;
  assign n8030 = ~n8028 & ~n8029 ;
  assign n8031 = ~n8019 & ~n8030 ;
  assign n8032 = n2568 & ~n3566 ;
  assign n8033 = ~x6 & n786 ;
  assign n8034 = n43 & n8033 ;
  assign n8035 = ~n8032 & ~n8034 ;
  assign n8036 = n4561 & ~n8035 ;
  assign n8037 = ~n8031 & ~n8036 ;
  assign n8038 = ~n8027 & n8037 ;
  assign n8039 = x15 & ~n8038 ;
  assign n8040 = ~n8024 & ~n8039 ;
  assign n8041 = n4155 & ~n8040 ;
  assign n8042 = n3462 & n4513 ;
  assign n8043 = n743 & n3561 ;
  assign n8044 = ~x2 & n2224 ;
  assign n8045 = n6452 & n8044 ;
  assign n8046 = n4330 & n6286 ;
  assign n8047 = ~n8045 & ~n8046 ;
  assign n8048 = ~n8043 & n8047 ;
  assign n8049 = n122 & ~n8048 ;
  assign n8050 = ~n8042 & ~n8049 ;
  assign n8051 = ~x1 & n8050 ;
  assign n8052 = n1295 & n4898 ;
  assign n8053 = n145 & n4644 ;
  assign n8054 = ~n8052 & ~n8053 ;
  assign n8055 = n7748 & ~n8054 ;
  assign n8056 = ~n311 & ~n954 ;
  assign n8057 = ~n58 & n8056 ;
  assign n8058 = n1264 & ~n3013 ;
  assign n8059 = ~n727 & n4898 ;
  assign n8060 = ~n8058 & ~n8059 ;
  assign n8061 = n371 & ~n5888 ;
  assign n8062 = n7181 & ~n8061 ;
  assign n8063 = ~n8060 & n8062 ;
  assign n8064 = ~n8057 & n8063 ;
  assign n8065 = ~n8055 & ~n8064 ;
  assign n8066 = n406 & n784 ;
  assign n8067 = n7201 & n8066 ;
  assign n8068 = n8067 ^ x1 ;
  assign n8069 = n198 & n471 ;
  assign n8070 = n8069 ^ n306 ;
  assign n8071 = ~n8068 & n8070 ;
  assign n8072 = n8071 ^ n8069 ;
  assign n8073 = n306 & n8072 ;
  assign n8074 = n8073 ^ x1 ;
  assign n8075 = n8065 & n8074 ;
  assign n8076 = ~n8019 & ~n8075 ;
  assign n8077 = ~n8051 & n8076 ;
  assign n8078 = n712 & n1078 ;
  assign n8079 = n3088 ^ n2806 ;
  assign n8080 = n8079 ^ n2806 ;
  assign n8081 = n2806 ^ n1246 ;
  assign n8082 = n8081 ^ n2806 ;
  assign n8083 = n8080 & n8082 ;
  assign n8084 = n8083 ^ n2806 ;
  assign n8085 = ~x4 & n8084 ;
  assign n8086 = n8085 ^ n2806 ;
  assign n8087 = n8078 & n8086 ;
  assign n8088 = ~n8077 & ~n8087 ;
  assign n8089 = n2658 & n7378 ;
  assign n8090 = n3777 & n4813 ;
  assign n8091 = ~n8089 & ~n8090 ;
  assign n8092 = ~x15 & ~n700 ;
  assign n8093 = ~n4829 & ~n8092 ;
  assign n8094 = n4513 & n8093 ;
  assign n8095 = x8 & n1270 ;
  assign n8096 = n6574 & n8095 ;
  assign n8097 = ~n8094 & ~n8096 ;
  assign n8098 = ~n8091 & ~n8097 ;
  assign n8099 = n8088 & ~n8098 ;
  assign n8100 = ~n8041 & n8099 ;
  assign n8101 = ~n8016 & n8100 ;
  assign n8128 = ~n1240 & n3530 ;
  assign n8129 = n198 & n8128 ;
  assign n8130 = n199 & n1948 ;
  assign n8131 = ~n4330 & ~n8130 ;
  assign n8132 = n122 & ~n8131 ;
  assign n8103 = ~x2 & n2239 ;
  assign n8133 = n1327 & n8103 ;
  assign n8134 = n406 & n8133 ;
  assign n8135 = ~n8132 & ~n8134 ;
  assign n8136 = n2591 & ~n8135 ;
  assign n8137 = n1682 & ~n7595 ;
  assign n8138 = n392 & n4023 ;
  assign n8139 = ~n2350 & ~n8138 ;
  assign n8140 = n2282 & ~n7082 ;
  assign n8141 = n8139 & ~n8140 ;
  assign n8142 = ~n8137 & n8141 ;
  assign n8143 = n3428 & ~n8142 ;
  assign n8144 = ~n8136 & ~n8143 ;
  assign n8145 = ~n8129 & n8144 ;
  assign n8146 = n3490 & ~n8145 ;
  assign n8147 = n928 & n2608 ;
  assign n8148 = n3208 & n8147 ;
  assign n8149 = n106 & n2271 ;
  assign n8150 = n226 & n8149 ;
  assign n8151 = ~n8148 & ~n8150 ;
  assign n8152 = n411 & ~n8151 ;
  assign n8153 = n759 & n1948 ;
  assign n8154 = ~n5838 & ~n8153 ;
  assign n8155 = n843 & n4513 ;
  assign n8156 = ~n8154 & n8155 ;
  assign n8157 = ~n8152 & ~n8156 ;
  assign n8158 = ~n673 & n3561 ;
  assign n8159 = ~x8 & n6436 ;
  assign n8160 = ~n8158 & ~n8159 ;
  assign n8161 = n787 & ~n8160 ;
  assign n8162 = ~x2 & ~n718 ;
  assign n8163 = n978 & ~n8162 ;
  assign n8164 = n850 & n8163 ;
  assign n8165 = n58 & n1563 ;
  assign n8166 = n6359 & n8165 ;
  assign n8167 = ~n8164 & ~n8166 ;
  assign n8168 = ~n8161 & n8167 ;
  assign n8169 = n3207 & ~n8168 ;
  assign n8170 = n719 & n4513 ;
  assign n8171 = n2115 & n7585 ;
  assign n8172 = n8170 & n8171 ;
  assign n8173 = ~n8169 & ~n8172 ;
  assign n8174 = n8157 & n8173 ;
  assign n8175 = ~n8146 & n8174 ;
  assign n8176 = ~x7 & ~n8175 ;
  assign n8102 = n466 & n2356 ;
  assign n8104 = n2684 & n8103 ;
  assign n8105 = n8102 & n8104 ;
  assign n8106 = n371 & n862 ;
  assign n8107 = n1247 & n8106 ;
  assign n8108 = n3186 & n8107 ;
  assign n8109 = n145 & n778 ;
  assign n8110 = ~n4774 & ~n8109 ;
  assign n8111 = n2271 & ~n8110 ;
  assign n8112 = n199 & n4656 ;
  assign n8113 = ~n8111 & ~n8112 ;
  assign n8114 = x14 & n524 ;
  assign n8115 = n2684 & n8114 ;
  assign n8116 = ~n8113 & n8115 ;
  assign n8117 = n3365 & n6872 ;
  assign n8118 = ~n248 & ~n6597 ;
  assign n8119 = n1656 & n8118 ;
  assign n8120 = n2684 & n8119 ;
  assign n8121 = n198 & n8120 ;
  assign n8122 = ~n8117 & ~n8121 ;
  assign n8123 = x14 & ~n8122 ;
  assign n8124 = ~n8116 & ~n8123 ;
  assign n8125 = ~n8108 & n8124 ;
  assign n8126 = n26 & ~n8125 ;
  assign n8127 = ~n8105 & ~n8126 ;
  assign n8177 = n8176 ^ n8127 ;
  assign n8178 = n8177 ^ n8127 ;
  assign n8179 = n1524 & n3702 ;
  assign n8180 = n874 & n8179 ;
  assign n8181 = ~x11 & n7103 ;
  assign n8182 = ~n1214 & ~n4035 ;
  assign n8183 = ~x2 & n8182 ;
  assign n8184 = n8181 & ~n8183 ;
  assign n8185 = n850 & n8184 ;
  assign n8186 = n5117 & ~n5121 ;
  assign n8187 = n3428 & ~n8186 ;
  assign n8188 = x0 & n8187 ;
  assign n8189 = ~n8185 & ~n8188 ;
  assign n8190 = ~n8180 & n8189 ;
  assign n8191 = n2653 & ~n8190 ;
  assign n8192 = ~x5 & n8102 ;
  assign n8193 = n8147 & n8192 ;
  assign n8194 = ~n8191 & ~n8193 ;
  assign n8195 = n8194 ^ n8127 ;
  assign n8196 = n8195 ^ n8127 ;
  assign n8197 = ~n8178 & n8196 ;
  assign n8198 = n8197 ^ n8127 ;
  assign n8199 = x1 & n8198 ;
  assign n8200 = n8199 ^ n8127 ;
  assign n8201 = n8101 & n8200 ;
  assign n8202 = ~n4672 & ~n8201 ;
  assign n8203 = ~n2263 & ~n4262 ;
  assign n8204 = x13 & n17 ;
  assign n8205 = x9 & n8204 ;
  assign n8206 = ~n8203 & n8205 ;
  assign n8207 = ~n3418 & ~n5130 ;
  assign n8208 = n8207 ^ n7594 ;
  assign n8209 = n8208 ^ n7594 ;
  assign n8210 = n7594 ^ x9 ;
  assign n8211 = n8210 ^ n7594 ;
  assign n8212 = ~n8209 & n8211 ;
  assign n8213 = n8212 ^ n7594 ;
  assign n8214 = x7 & n8213 ;
  assign n8215 = n8214 ^ n7594 ;
  assign n8216 = n261 & n8215 ;
  assign n8217 = x14 & n2637 ;
  assign n8218 = n1954 & ~n4273 ;
  assign n8219 = ~x10 & ~n7240 ;
  assign n8220 = ~n5463 & ~n8219 ;
  assign n8221 = n109 & ~n8220 ;
  assign n8222 = n511 & n5384 ;
  assign n8223 = ~n1423 & n4350 ;
  assign n8224 = n7363 & n8223 ;
  assign n8225 = ~n8222 & ~n8224 ;
  assign n8226 = ~x0 & ~n8225 ;
  assign n8227 = ~n8221 & ~n8226 ;
  assign n8228 = ~n8218 & n8227 ;
  assign n8229 = n8217 & ~n8228 ;
  assign n8230 = ~n8216 & ~n8229 ;
  assign n8231 = ~n8206 & n8230 ;
  assign n8232 = n1905 & n4542 ;
  assign n8233 = ~n240 & ~n260 ;
  assign n8234 = ~n8232 & n8233 ;
  assign n8235 = ~x12 & ~n8234 ;
  assign n8236 = n6160 & ~n8235 ;
  assign n8237 = ~n524 & n8236 ;
  assign n8238 = n2863 & ~n8237 ;
  assign n8239 = x1 & n8238 ;
  assign n8240 = n8231 & ~n8239 ;
  assign n8241 = n168 & ~n8240 ;
  assign n8242 = n60 & ~n7716 ;
  assign n8243 = ~n5215 & ~n8242 ;
  assign n8244 = n4014 & ~n8243 ;
  assign n8245 = ~n392 & ~n1010 ;
  assign n8246 = x0 & n8245 ;
  assign n8247 = ~n605 & ~n8246 ;
  assign n8248 = ~n759 & n8247 ;
  assign n8249 = n4253 & ~n8248 ;
  assign n8250 = ~n8244 & ~n8249 ;
  assign n8251 = n846 & ~n8250 ;
  assign n8252 = ~n60 & ~n1353 ;
  assign n8253 = n6956 & ~n8252 ;
  assign n8254 = x11 & n5976 ;
  assign n8255 = ~n4203 & ~n8254 ;
  assign n8256 = n5619 & ~n8255 ;
  assign n8257 = n1180 & ~n5516 ;
  assign n8258 = ~n8256 & ~n8257 ;
  assign n8259 = ~n8253 & n8258 ;
  assign n8260 = n5908 & ~n8259 ;
  assign n8261 = ~n8251 & ~n8260 ;
  assign n8262 = n1920 & ~n8261 ;
  assign n8263 = ~n1050 & ~n4014 ;
  assign n8264 = n224 & ~n8263 ;
  assign n8265 = ~n45 & ~n462 ;
  assign n8266 = ~n109 & n5908 ;
  assign n8267 = ~n8265 & n8266 ;
  assign n8268 = ~n8264 & ~n8267 ;
  assign n8269 = n5947 & ~n8268 ;
  assign n8270 = ~n8262 & ~n8269 ;
  assign n8271 = ~n8241 & n8270 ;
  assign n8276 = n4253 & n6973 ;
  assign n8277 = n846 & n8276 ;
  assign n8272 = n306 & ~n2468 ;
  assign n8273 = n105 & n6326 ;
  assign n8274 = ~n8272 & ~n8273 ;
  assign n8275 = n5431 & ~n8274 ;
  assign n8278 = n8277 ^ n8275 ;
  assign n8279 = ~x5 & n8278 ;
  assign n8280 = n8279 ^ n8277 ;
  assign n8281 = n8271 & ~n8280 ;
  assign n8282 = ~n3566 & ~n8281 ;
  assign n8283 = x14 & n1214 ;
  assign n8284 = n2471 & n8283 ;
  assign n8285 = n6392 & n8284 ;
  assign n8286 = n4253 & n8285 ;
  assign n8328 = n3862 & n6562 ;
  assign n8329 = n928 & n4253 ;
  assign n8330 = n2814 & n8329 ;
  assign n8331 = ~x7 & n20 ;
  assign n8332 = n248 & n8331 ;
  assign n8333 = n226 & n4206 ;
  assign n8334 = ~n8332 & ~n8333 ;
  assign n8335 = n1349 & ~n8334 ;
  assign n8336 = n8335 ^ x3 ;
  assign n8337 = n8336 ^ n8335 ;
  assign n8338 = n8337 ^ n8330 ;
  assign n8339 = n3264 & n5291 ;
  assign n8340 = ~n1169 & n8339 ;
  assign n8341 = ~x2 & n66 ;
  assign n8342 = n641 & n8341 ;
  assign n8343 = n20 & n1028 ;
  assign n8344 = ~n8342 & ~n8343 ;
  assign n8345 = ~n8340 & n8344 ;
  assign n8346 = n8345 ^ x12 ;
  assign n8347 = ~n8345 & n8346 ;
  assign n8348 = n8347 ^ n8335 ;
  assign n8349 = n8348 ^ n8345 ;
  assign n8350 = n8338 & ~n8349 ;
  assign n8351 = n8350 ^ n8347 ;
  assign n8352 = n8351 ^ n8345 ;
  assign n8353 = ~n8330 & ~n8352 ;
  assign n8354 = n8353 ^ n8330 ;
  assign n8355 = x14 & n8354 ;
  assign n8356 = ~n8328 & ~n8355 ;
  assign n8357 = n411 & ~n8356 ;
  assign n8359 = n1665 & n1693 ;
  assign n8360 = ~n5735 & ~n8359 ;
  assign n8358 = n2290 & n6104 ;
  assign n8361 = n8360 ^ n8358 ;
  assign n8362 = n8361 ^ n8360 ;
  assign n8363 = n8360 ^ n58 ;
  assign n8364 = n8363 ^ n8360 ;
  assign n8365 = n8362 & ~n8364 ;
  assign n8366 = n8365 ^ n8360 ;
  assign n8367 = ~n928 & ~n8366 ;
  assign n8368 = n8367 ^ n8360 ;
  assign n8369 = n779 & ~n8368 ;
  assign n8370 = n492 & n7178 ;
  assign n8371 = ~x9 & n168 ;
  assign n8372 = n3555 & n8371 ;
  assign n8373 = ~n8370 & ~n8372 ;
  assign n8374 = n20 & ~n8373 ;
  assign n8375 = n375 & n1656 ;
  assign n8376 = n104 & n5469 ;
  assign n8377 = ~n8375 & ~n8376 ;
  assign n8378 = n740 & ~n8377 ;
  assign n8379 = n196 & n1030 ;
  assign n8380 = ~n785 & ~n8379 ;
  assign n8381 = n76 & ~n8380 ;
  assign n8382 = n1682 & n8381 ;
  assign n8383 = ~n8378 & ~n8382 ;
  assign n8384 = ~n8374 & n8383 ;
  assign n8385 = x11 & ~n8384 ;
  assign n8386 = ~n8369 & ~n8385 ;
  assign n8387 = n1042 & ~n8386 ;
  assign n8388 = ~x2 & n517 ;
  assign n8389 = n1954 & n8388 ;
  assign n8390 = ~n7139 & n8389 ;
  assign n8391 = ~n741 & n4684 ;
  assign n8392 = ~n8390 & ~n8391 ;
  assign n8393 = n5908 & ~n8392 ;
  assign n8394 = x10 & n8393 ;
  assign n8395 = n217 & n1030 ;
  assign n8396 = n1095 & n8395 ;
  assign n8397 = n713 & n847 ;
  assign n8398 = n65 & ~n354 ;
  assign n8399 = ~n8397 & ~n8398 ;
  assign n8400 = ~n8396 & n8399 ;
  assign n8401 = n8400 ^ n529 ;
  assign n8402 = n8401 ^ n8400 ;
  assign n8403 = ~n24 & ~n346 ;
  assign n8404 = ~n517 & ~n8403 ;
  assign n8405 = n1095 & ~n8404 ;
  assign n8406 = n176 & n1435 ;
  assign n8407 = n633 & n8406 ;
  assign n8408 = ~n8405 & ~n8407 ;
  assign n8409 = n8408 ^ n8400 ;
  assign n8410 = n8409 ^ n8400 ;
  assign n8411 = n8402 & ~n8410 ;
  assign n8412 = n8411 ^ n8400 ;
  assign n8413 = ~x0 & ~n8412 ;
  assign n8414 = n8413 ^ n8400 ;
  assign n8415 = n1034 & ~n8414 ;
  assign n8416 = n71 & n517 ;
  assign n8417 = n712 & n978 ;
  assign n8418 = n55 & n8417 ;
  assign n8419 = ~n8416 & ~n8418 ;
  assign n8420 = n6146 & ~n8419 ;
  assign n8421 = ~n8415 & ~n8420 ;
  assign n8422 = ~n8394 & n8421 ;
  assign n8423 = ~n8387 & n8422 ;
  assign n8424 = ~n8357 & n8423 ;
  assign n8287 = n196 & n4180 ;
  assign n8288 = ~n750 & n4014 ;
  assign n8289 = n8288 ^ n76 ;
  assign n8290 = n8289 ^ n8288 ;
  assign n8291 = n8288 ^ n1806 ;
  assign n8292 = n8291 ^ n8288 ;
  assign n8293 = n8290 & n8292 ;
  assign n8294 = n8293 ^ n8288 ;
  assign n8295 = ~x12 & n8294 ;
  assign n8296 = n8295 ^ n8288 ;
  assign n8297 = n1165 & n8296 ;
  assign n8298 = ~n8287 & ~n8297 ;
  assign n8299 = n277 & ~n8298 ;
  assign n8300 = ~x7 & n524 ;
  assign n8301 = ~n4851 & ~n8300 ;
  assign n8302 = x0 & ~n8301 ;
  assign n8303 = ~n1170 & ~n8302 ;
  assign n8304 = ~x1 & n712 ;
  assign n8305 = ~n8303 & n8304 ;
  assign n8306 = n2301 & n8305 ;
  assign n8307 = ~n8299 & ~n8306 ;
  assign n8308 = n65 & n845 ;
  assign n8309 = n262 & n524 ;
  assign n8310 = ~n8308 & ~n8309 ;
  assign n8311 = x1 & ~n8310 ;
  assign n8312 = n8311 ^ n65 ;
  assign n8313 = n8312 ^ n8311 ;
  assign n8314 = n8311 ^ n6129 ;
  assign n8315 = n8314 ^ n8311 ;
  assign n8316 = n8313 & n8315 ;
  assign n8317 = n8316 ^ n8311 ;
  assign n8318 = ~x0 & n8317 ;
  assign n8319 = n8318 ^ n8311 ;
  assign n8320 = ~n2678 & n8319 ;
  assign n8321 = ~x3 & n524 ;
  assign n8322 = ~n77 & ~n1781 ;
  assign n8323 = n8321 & ~n8322 ;
  assign n8324 = n1042 & n8323 ;
  assign n8325 = ~n8320 & ~n8324 ;
  assign n8326 = n1263 & ~n8325 ;
  assign n8327 = n8307 & ~n8326 ;
  assign n8425 = n8424 ^ n8327 ;
  assign n8426 = ~x8 & n8425 ;
  assign n8427 = n8426 ^ n8424 ;
  assign n8428 = ~n8286 & n8427 ;
  assign n8429 = n2701 & ~n8428 ;
  assign n8430 = ~n8282 & ~n8429 ;
  assign n8431 = ~n8202 & n8430 ;
  assign n8432 = n146 & n4019 ;
  assign n8433 = n2711 & n8432 ;
  assign n8434 = ~n1738 & ~n2270 ;
  assign n8435 = n28 & ~n8434 ;
  assign n8436 = ~n106 & ~n556 ;
  assign n8437 = n1806 & ~n8436 ;
  assign n8438 = ~n8435 & ~n8437 ;
  assign n8439 = n1656 & ~n8438 ;
  assign n8440 = n442 & n5463 ;
  assign n8441 = n2394 & n8440 ;
  assign n8442 = ~x13 & ~n3908 ;
  assign n8443 = n349 & n456 ;
  assign n8444 = n8442 & n8443 ;
  assign n8445 = ~n8441 & ~n8444 ;
  assign n8446 = n1841 & n4313 ;
  assign n8447 = n1665 & n8446 ;
  assign n8448 = n8445 & ~n8447 ;
  assign n8449 = ~n8439 & n8448 ;
  assign n8450 = ~n8433 & n8449 ;
  assign n8451 = n20 & ~n8450 ;
  assign n8452 = ~n1630 & ~n7897 ;
  assign n8453 = ~n110 & n562 ;
  assign n8454 = n7217 & n8453 ;
  assign n8455 = n55 & n292 ;
  assign n8456 = n2799 & n8455 ;
  assign n8457 = ~n8454 & ~n8456 ;
  assign n8458 = n740 & ~n8457 ;
  assign n8459 = ~n8452 & n8458 ;
  assign n8460 = n8459 ^ n8451 ;
  assign n8461 = n124 & n1656 ;
  assign n8462 = n1117 & n7611 ;
  assign n8463 = ~n8461 & ~n8462 ;
  assign n8464 = ~x2 & x4 ;
  assign n8465 = n5729 & n8464 ;
  assign n8466 = ~n8463 & n8465 ;
  assign n8467 = n168 & n2754 ;
  assign n8468 = n124 & n2873 ;
  assign n8469 = x13 & n8468 ;
  assign n8470 = ~n8467 & ~n8469 ;
  assign n8471 = n332 & n1618 ;
  assign n8472 = ~n8470 & n8471 ;
  assign n8473 = ~n8466 & ~n8472 ;
  assign n8474 = n8473 ^ x0 ;
  assign n8475 = n8474 ^ n8473 ;
  assign n8476 = ~n467 & n1327 ;
  assign n8477 = ~n214 & ~n4333 ;
  assign n8478 = n8476 & ~n8477 ;
  assign n8479 = ~x8 & n1656 ;
  assign n8480 = n55 & n8479 ;
  assign n8481 = ~n8478 & ~n8480 ;
  assign n8482 = n1624 & ~n8481 ;
  assign n8483 = n8482 ^ n8473 ;
  assign n8484 = n8475 & ~n8483 ;
  assign n8485 = n8484 ^ n8473 ;
  assign n8486 = n8485 ^ n8451 ;
  assign n8487 = n8460 & ~n8486 ;
  assign n8488 = n8487 ^ n8484 ;
  assign n8489 = n8488 ^ n8473 ;
  assign n8490 = n8489 ^ n8459 ;
  assign n8491 = ~n8451 & ~n8490 ;
  assign n8492 = n8491 ^ n8451 ;
  assign n8493 = n623 & n8492 ;
  assign n8494 = n2030 ^ n795 ;
  assign n8495 = n8494 ^ n2030 ;
  assign n8496 = n2030 ^ n1601 ;
  assign n8497 = n8496 ^ n2030 ;
  assign n8498 = n8495 & n8497 ;
  assign n8499 = n8498 ^ n2030 ;
  assign n8500 = ~x3 & n8499 ;
  assign n8501 = n8500 ^ n2030 ;
  assign n8502 = n778 & n8501 ;
  assign n8503 = ~x4 & n65 ;
  assign n8504 = n5029 & n8503 ;
  assign n8505 = x5 & n8504 ;
  assign n8506 = ~n8502 & ~n8505 ;
  assign n8507 = n7665 & ~n8506 ;
  assign n8508 = x2 & n1667 ;
  assign n8509 = n1265 & n8508 ;
  assign n8510 = n1608 & n8509 ;
  assign n8511 = n463 & ~n3803 ;
  assign n8512 = n1563 & n1678 ;
  assign n8513 = n8442 & n8512 ;
  assign n8514 = ~n8511 & ~n8513 ;
  assign n8515 = x2 & n168 ;
  assign n8516 = ~n8514 & n8515 ;
  assign n8517 = ~n467 & n1682 ;
  assign n8518 = n105 & n1626 ;
  assign n8519 = n8517 & n8518 ;
  assign n8520 = ~n8516 & ~n8519 ;
  assign n8521 = x1 & ~n8520 ;
  assign n8522 = ~n8510 & ~n8521 ;
  assign n8523 = ~n8507 & n8522 ;
  assign n8524 = n2370 & ~n5714 ;
  assign n8525 = n7948 & ~n8524 ;
  assign n8526 = n1683 & n8525 ;
  assign n8527 = ~n1327 & ~n6037 ;
  assign n8528 = ~n2183 & ~n8527 ;
  assign n8529 = ~x0 & ~n56 ;
  assign n8530 = n8528 & n8529 ;
  assign n8531 = n795 & n5129 ;
  assign n8532 = ~n1631 & ~n8531 ;
  assign n8533 = n1874 & ~n8532 ;
  assign n8534 = ~n8530 & ~n8533 ;
  assign n8535 = ~n8526 & n8534 ;
  assign n8536 = n1003 & ~n8535 ;
  assign n8537 = n463 & n1327 ;
  assign n8538 = n43 & n8537 ;
  assign n8539 = n164 & ~n5998 ;
  assign n8540 = ~n344 & ~n8539 ;
  assign n8541 = n8538 & n8540 ;
  assign n8542 = n168 & n1382 ;
  assign n8543 = ~n3803 & n8109 ;
  assign n8544 = n8542 & n8543 ;
  assign n8545 = ~n8541 & ~n8544 ;
  assign n8546 = ~n8536 & n8545 ;
  assign n8547 = n260 & ~n8546 ;
  assign n8548 = n8523 & ~n8547 ;
  assign n8549 = ~n8493 & n8548 ;
  assign n8550 = n1025 & ~n8549 ;
  assign n8551 = ~n56 & n195 ;
  assign n8552 = n373 & ~n3798 ;
  assign n8553 = ~n1034 & n8552 ;
  assign n8554 = ~n8551 & ~n8553 ;
  assign n8555 = n779 & ~n8554 ;
  assign n8556 = ~x6 & n8555 ;
  assign n8557 = n3798 & n7409 ;
  assign n8558 = x1 & n2633 ;
  assign n8559 = ~x4 & n8558 ;
  assign n8560 = ~n8021 & ~n8559 ;
  assign n8561 = n1679 & ~n8560 ;
  assign n8562 = ~x7 & n312 ;
  assign n8563 = ~x3 & n3666 ;
  assign n8564 = ~n8562 & ~n8563 ;
  assign n8565 = n4027 & ~n8564 ;
  assign n8566 = ~n8561 & ~n8565 ;
  assign n8567 = x14 & ~n8566 ;
  assign n8568 = ~n8557 & ~n8567 ;
  assign n8569 = ~n8556 & n8568 ;
  assign n8570 = n1363 & ~n8569 ;
  assign n8571 = ~n2569 & ~n4338 ;
  assign n8572 = ~x6 & ~n8571 ;
  assign n8573 = ~n8562 & ~n8572 ;
  assign n8574 = n307 & ~n8573 ;
  assign n8576 = n3578 ^ x3 ;
  assign n8575 = n3578 ^ x7 ;
  assign n8577 = n8576 ^ n8575 ;
  assign n8578 = n8577 ^ n8576 ;
  assign n8579 = n8578 ^ n3578 ;
  assign n8580 = n8576 ^ n3578 ;
  assign n8581 = n8578 & ~n8580 ;
  assign n8582 = n8581 ^ n8579 ;
  assign n8583 = n249 & n8582 ;
  assign n8584 = n8583 ^ n8581 ;
  assign n8585 = n8579 & n8584 ;
  assign n8586 = n8585 ^ n8581 ;
  assign n8587 = n6905 & n8586 ;
  assign n8588 = ~n8574 & ~n8587 ;
  assign n8589 = x11 & n784 ;
  assign n8590 = ~n8588 & n8589 ;
  assign n8591 = ~x10 & n226 ;
  assign n8593 = ~x4 & n2806 ;
  assign n8594 = n4007 & n8593 ;
  assign n8595 = n1422 & n2226 ;
  assign n8596 = n2584 & n6905 ;
  assign n8597 = ~n3803 & n8596 ;
  assign n8598 = ~n8595 & ~n8597 ;
  assign n8599 = ~n8594 & n8598 ;
  assign n8592 = n306 & ~n2702 ;
  assign n8600 = n8599 ^ n8592 ;
  assign n8601 = n8600 ^ n8599 ;
  assign n8602 = n8599 ^ x7 ;
  assign n8603 = n8602 ^ n8599 ;
  assign n8604 = n8601 & ~n8603 ;
  assign n8605 = n8604 ^ n8599 ;
  assign n8606 = ~x3 & ~n8605 ;
  assign n8607 = n8606 ^ n8599 ;
  assign n8608 = n8591 & ~n8607 ;
  assign n8609 = x7 & ~n225 ;
  assign n8610 = x6 & n845 ;
  assign n8611 = ~n21 & ~n5189 ;
  assign n8612 = n8610 & n8611 ;
  assign n8613 = n306 & n8612 ;
  assign n8614 = ~n8609 & n8613 ;
  assign n8615 = ~x2 & n8614 ;
  assign n8616 = ~n8608 & ~n8615 ;
  assign n8617 = ~n8590 & n8616 ;
  assign n8618 = ~x2 & x6 ;
  assign n8619 = ~n3427 & ~n8618 ;
  assign n8620 = n1494 & n2583 ;
  assign n8621 = n21 & n3091 ;
  assign n8622 = ~n8620 & ~n8621 ;
  assign n8623 = ~n8619 & ~n8622 ;
  assign n8624 = n366 & n7022 ;
  assign n8625 = n3568 & n8624 ;
  assign n8626 = ~n8623 & ~n8625 ;
  assign n8627 = n306 & ~n8626 ;
  assign n8628 = n225 & n1422 ;
  assign n8629 = n65 & n8628 ;
  assign n8630 = n301 & n8593 ;
  assign n8631 = ~x2 & n2575 ;
  assign n8632 = n314 ^ x7 ;
  assign n8633 = n8632 ^ n314 ;
  assign n8634 = n6448 ^ n314 ;
  assign n8635 = n8633 & n8634 ;
  assign n8636 = n8635 ^ n314 ;
  assign n8637 = n8631 & n8636 ;
  assign n8638 = ~n8630 & ~n8637 ;
  assign n8639 = ~n8629 & n8638 ;
  assign n8640 = n261 & ~n8639 ;
  assign n8641 = n1581 & n2583 ;
  assign n8642 = n178 & n3091 ;
  assign n8643 = ~n8641 & ~n8642 ;
  assign n8644 = n65 & ~n8643 ;
  assign n8645 = ~n42 & ~n8464 ;
  assign n8646 = ~n700 & ~n4253 ;
  assign n8647 = ~x3 & ~n2583 ;
  assign n8648 = n8646 & n8647 ;
  assign n8649 = ~n8645 & n8648 ;
  assign n8650 = ~n8644 & ~n8649 ;
  assign n8651 = n2599 & ~n8650 ;
  assign n8652 = x4 & n3427 ;
  assign n8653 = ~n442 & n2458 ;
  assign n8654 = ~n314 & ~n700 ;
  assign n8655 = n8653 & n8654 ;
  assign n8656 = n8652 & n8655 ;
  assign n8657 = ~n8651 & ~n8656 ;
  assign n8658 = ~n8640 & n8657 ;
  assign n8659 = ~n8627 & n8658 ;
  assign n8660 = n845 & ~n8659 ;
  assign n8661 = n1514 & n2881 ;
  assign n8662 = n318 & n2684 ;
  assign n8663 = ~n8661 & ~n8662 ;
  assign n8664 = n1555 & n7217 ;
  assign n8665 = n261 & n8664 ;
  assign n8666 = ~n109 & ~n2477 ;
  assign n8667 = n1476 & n4422 ;
  assign n8668 = n8666 & n8667 ;
  assign n8669 = ~n8665 & ~n8668 ;
  assign n8670 = ~n8663 & ~n8669 ;
  assign n8671 = n1495 & n8114 ;
  assign n8672 = n1042 & n2562 ;
  assign n8673 = n8671 & n8672 ;
  assign n8674 = ~n8670 & ~n8673 ;
  assign n8675 = ~n8660 & n8674 ;
  assign n8676 = n8675 ^ x15 ;
  assign n8677 = n8676 ^ n8675 ;
  assign n8678 = n8021 & n8309 ;
  assign n8679 = n348 & n2633 ;
  assign n8680 = n845 & n3427 ;
  assign n8681 = n8679 & n8680 ;
  assign n8682 = ~n8678 & ~n8681 ;
  assign n8683 = ~n7129 & ~n8682 ;
  assign n8684 = ~x4 & n3098 ;
  assign n8685 = n66 & n862 ;
  assign n8686 = ~n1042 & ~n4014 ;
  assign n8687 = n20 & ~n8686 ;
  assign n8688 = ~n8685 & ~n8687 ;
  assign n8689 = n8321 & ~n8688 ;
  assign n8690 = n8591 & n8679 ;
  assign n8691 = n67 & n8300 ;
  assign n8692 = ~n8690 & ~n8691 ;
  assign n8693 = ~n8689 & n8692 ;
  assign n8694 = n8684 & ~n8693 ;
  assign n8695 = ~n8683 & ~n8694 ;
  assign n8696 = n8695 ^ n8675 ;
  assign n8697 = n8677 & n8696 ;
  assign n8698 = n8697 ^ n8675 ;
  assign n8699 = n8617 & n8698 ;
  assign n8700 = ~n8570 & n8699 ;
  assign n8701 = ~x5 & ~n8700 ;
  assign n8702 = ~n8300 & ~n8610 ;
  assign n8703 = ~n2881 & ~n8702 ;
  assign n8704 = n929 & n1270 ;
  assign n8705 = ~x2 & n311 ;
  assign n8706 = ~x0 & n8705 ;
  assign n8707 = ~n8704 & ~n8706 ;
  assign n8708 = n366 & ~n8707 ;
  assign n8709 = n652 & ~n8645 ;
  assign n8710 = ~n8708 & ~n8709 ;
  assign n8711 = n159 & ~n8710 ;
  assign n8712 = n3019 & n7646 ;
  assign n8713 = n8645 ^ n352 ;
  assign n8714 = x0 & ~n8713 ;
  assign n8715 = n8714 ^ n352 ;
  assign n8716 = n345 & n8715 ;
  assign n8717 = ~n70 & ~n7129 ;
  assign n8718 = n3010 & n8551 ;
  assign n8719 = ~n8717 & ~n8718 ;
  assign n8720 = n4015 & ~n8719 ;
  assign n8721 = ~n8716 & ~n8720 ;
  assign n8722 = ~n8712 & n8721 ;
  assign n8723 = ~n8711 & n8722 ;
  assign n8724 = n8703 & ~n8723 ;
  assign n8725 = ~x2 & n225 ;
  assign n8726 = n261 & n2806 ;
  assign n8727 = n8725 & n8726 ;
  assign n8728 = n249 & n2562 ;
  assign n8729 = n233 & n8728 ;
  assign n8730 = ~n8727 & ~n8729 ;
  assign n8731 = n8321 & ~n8730 ;
  assign n8732 = ~x6 & n159 ;
  assign n8733 = n1545 & n8732 ;
  assign n8734 = n1050 & n1905 ;
  assign n8735 = n8733 & n8734 ;
  assign n8736 = ~x7 & ~n70 ;
  assign n8737 = n3128 ^ x14 ;
  assign n8738 = n6632 ^ x14 ;
  assign n8739 = n8738 ^ x6 ;
  assign n8740 = n8739 ^ n6632 ;
  assign n8741 = n8740 ^ n8737 ;
  assign n8742 = n524 ^ x6 ;
  assign n8743 = n524 & n8742 ;
  assign n8744 = n8743 ^ n6632 ;
  assign n8745 = n8744 ^ n524 ;
  assign n8746 = n8741 & n8745 ;
  assign n8747 = n8746 ^ n8743 ;
  assign n8748 = n8747 ^ n524 ;
  assign n8749 = ~n8737 & n8748 ;
  assign n8750 = n8736 & n8749 ;
  assign n8751 = ~n8735 & ~n8750 ;
  assign n8752 = ~n8731 & n8751 ;
  assign n8753 = ~n2702 & n3960 ;
  assign n8754 = n306 & n8591 ;
  assign n8755 = n8753 & n8754 ;
  assign n8756 = ~n66 & ~n352 ;
  assign n8757 = ~n2612 & ~n8756 ;
  assign n8758 = ~n306 & ~n8757 ;
  assign n8759 = n2282 & ~n2839 ;
  assign n8760 = ~n249 & ~n8759 ;
  assign n8761 = ~n6992 & ~n8760 ;
  assign n8762 = ~n66 & ~n332 ;
  assign n8763 = ~n2839 & n8762 ;
  assign n8764 = ~n2477 & ~n8763 ;
  assign n8765 = n8761 & n8764 ;
  assign n8766 = n8758 & n8765 ;
  assign n8767 = ~n8755 & ~n8766 ;
  assign n8768 = n4344 & ~n8767 ;
  assign n8769 = x6 & ~n1092 ;
  assign n8770 = ~n302 & n8769 ;
  assign n8772 = ~x0 & n8464 ;
  assign n8771 = n6905 ^ n55 ;
  assign n8773 = n8772 ^ n8771 ;
  assign n8774 = n8773 ^ n6905 ;
  assign n8779 = n8774 ^ n8771 ;
  assign n8780 = n8779 ^ n6905 ;
  assign n8781 = n8780 ^ n6905 ;
  assign n8782 = ~x4 & n6490 ;
  assign n8783 = n8782 ^ n8771 ;
  assign n8784 = n8783 ^ n8771 ;
  assign n8785 = n8784 ^ n6905 ;
  assign n8786 = n8781 & n8785 ;
  assign n8775 = n8771 ^ n2973 ;
  assign n8776 = n8775 ^ n8774 ;
  assign n8777 = n8776 ^ n6905 ;
  assign n8778 = n8774 & n8777 ;
  assign n8787 = n8786 ^ n8778 ;
  assign n8788 = n8787 ^ n8774 ;
  assign n8789 = n8778 ^ n6905 ;
  assign n8790 = n8789 ^ n8780 ;
  assign n8791 = ~n6905 & n8790 ;
  assign n8792 = n8791 ^ n8778 ;
  assign n8793 = n8788 & n8792 ;
  assign n8794 = n8793 ^ n8786 ;
  assign n8795 = n8794 ^ n8791 ;
  assign n8796 = n8795 ^ n8774 ;
  assign n8797 = n8796 ^ n6905 ;
  assign n8798 = n8797 ^ n8780 ;
  assign n8799 = n8798 ^ n55 ;
  assign n8800 = ~n8770 & ~n8799 ;
  assign n8801 = n8114 & ~n8800 ;
  assign n8802 = x6 & ~x15 ;
  assign n8803 = n74 & n8802 ;
  assign n8804 = n6448 & n8803 ;
  assign n8805 = n348 & ~n1270 ;
  assign n8806 = ~n7473 & n8805 ;
  assign n8807 = x2 & n8806 ;
  assign n8808 = x2 & ~x15 ;
  assign n8809 = ~x6 & ~x14 ;
  assign n8810 = n8808 & n8809 ;
  assign n8811 = n442 & n8810 ;
  assign n8812 = ~n8807 & ~n8811 ;
  assign n8813 = ~n8804 & n8812 ;
  assign n8814 = n195 & ~n8813 ;
  assign n8815 = n442 & ~n8809 ;
  assign n8816 = ~n6991 & n8815 ;
  assign n8817 = ~n8806 & ~n8816 ;
  assign n8818 = x4 & ~n8817 ;
  assign n8819 = ~n741 & n8818 ;
  assign n8820 = ~x3 & n249 ;
  assign n8821 = n8803 & n8820 ;
  assign n8822 = ~x4 & n318 ;
  assign n8823 = n8802 & n8822 ;
  assign n8824 = n4422 & n8823 ;
  assign n8825 = ~n8821 & ~n8824 ;
  assign n8826 = n8825 ^ x0 ;
  assign n8827 = n8826 ^ n8825 ;
  assign n8828 = x1 & ~n6097 ;
  assign n8829 = ~x15 & n314 ;
  assign n8830 = n8652 & ~n8829 ;
  assign n8831 = ~n8828 & n8830 ;
  assign n8832 = n8831 ^ n8825 ;
  assign n8833 = n8827 & ~n8832 ;
  assign n8834 = n8833 ^ n8825 ;
  assign n8835 = ~n8819 & n8834 ;
  assign n8836 = ~n8814 & n8835 ;
  assign n8837 = n845 & ~n8836 ;
  assign n8838 = n1270 & n2608 ;
  assign n8839 = n524 & n8838 ;
  assign n8840 = n4954 & n8839 ;
  assign n8841 = ~n8837 & ~n8840 ;
  assign n8842 = ~n8801 & n8841 ;
  assign n8843 = n2848 & ~n8842 ;
  assign n8844 = ~n8768 & ~n8843 ;
  assign n8845 = n8752 & n8844 ;
  assign n8846 = ~n8724 & n8845 ;
  assign n8847 = ~n8701 & n8846 ;
  assign n8848 = ~n2754 & ~n2824 ;
  assign n8849 = ~n265 & ~n8848 ;
  assign n8850 = ~n8847 & n8849 ;
  assign n8851 = ~n8550 & ~n8850 ;
  assign n8852 = n8431 & n8851 ;
  assign n8853 = ~x7 & n1515 ;
  assign n8877 = n26 & n1708 ;
  assign n8854 = n225 & n4942 ;
  assign n8855 = n196 & n8854 ;
  assign n8856 = n730 & n2528 ;
  assign n8857 = n978 & n3908 ;
  assign n8858 = ~n2607 & n8857 ;
  assign n8859 = ~n8856 & ~n8858 ;
  assign n8860 = n168 & ~n8859 ;
  assign n8861 = ~n8855 & ~n8860 ;
  assign n8862 = n1095 & ~n8861 ;
  assign n8863 = ~x0 & n352 ;
  assign n8864 = n4280 & n8863 ;
  assign n8865 = ~n489 & n6163 ;
  assign n8866 = ~n6973 & ~n8865 ;
  assign n8867 = ~n8645 & ~n8866 ;
  assign n8868 = ~n8864 & ~n8867 ;
  assign n8869 = n168 & ~n8868 ;
  assign n8870 = n561 & n4942 ;
  assign n8871 = n6436 & n8870 ;
  assign n8872 = ~x4 & n8871 ;
  assign n8873 = ~n8869 & ~n8872 ;
  assign n8874 = ~n8862 & n8873 ;
  assign n8878 = n8877 ^ n8874 ;
  assign n8879 = n8878 ^ n8874 ;
  assign n8875 = n8874 ^ n8114 ;
  assign n8876 = n8875 ^ n8874 ;
  assign n8880 = n8879 ^ n8876 ;
  assign n8881 = n8874 ^ x0 ;
  assign n8882 = n8881 ^ n8874 ;
  assign n8883 = n8882 ^ n8879 ;
  assign n8884 = n8879 & ~n8883 ;
  assign n8885 = n8884 ^ n8879 ;
  assign n8886 = n8880 & n8885 ;
  assign n8887 = n8886 ^ n8884 ;
  assign n8888 = n8887 ^ n8874 ;
  assign n8889 = n8888 ^ n8879 ;
  assign n8890 = ~x1 & ~n8889 ;
  assign n8891 = n8890 ^ n8874 ;
  assign n8892 = n8853 & ~n8891 ;
  assign n8893 = n348 & n2848 ;
  assign n8894 = n4605 & n8893 ;
  assign n8895 = n345 & n858 ;
  assign n8896 = n4087 & n8895 ;
  assign n8897 = ~n8894 & ~n8896 ;
  assign n8898 = ~n3803 & n6823 ;
  assign n8899 = n106 & n740 ;
  assign n8900 = n798 & n8464 ;
  assign n8901 = ~n8899 & ~n8900 ;
  assign n8902 = ~n1658 & ~n8901 ;
  assign n8903 = ~n8898 & ~n8902 ;
  assign n8904 = ~n8897 & ~n8903 ;
  assign n8905 = n367 & n7431 ;
  assign n8906 = n2326 & n2536 ;
  assign n8907 = ~n8905 & ~n8906 ;
  assign n8908 = n277 & n845 ;
  assign n8909 = n1909 & n8908 ;
  assign n8910 = n6563 & n8909 ;
  assign n8911 = n4582 & n7337 ;
  assign n8912 = n1648 & n8911 ;
  assign n8913 = ~n8910 & ~n8912 ;
  assign n8914 = ~n8907 & ~n8913 ;
  assign n8915 = ~x4 & n20 ;
  assign n8916 = ~n43 & ~n8772 ;
  assign n8917 = ~n8915 & n8916 ;
  assign n8918 = n730 & n8893 ;
  assign n8919 = n1515 & ~n1658 ;
  assign n8920 = n8918 & n8919 ;
  assign n8921 = ~n8917 & n8920 ;
  assign n8922 = ~n8914 & ~n8921 ;
  assign n8923 = ~n8904 & n8922 ;
  assign n8924 = ~n8892 & n8923 ;
  assign n8925 = n2975 & n4770 ;
  assign n8926 = n2613 & n5225 ;
  assign n8927 = x8 & n8926 ;
  assign n8928 = ~n8925 & ~n8927 ;
  assign n8929 = n1382 & n6562 ;
  assign n8930 = x12 & n67 ;
  assign n8931 = n1214 ^ n828 ;
  assign n8932 = n8931 ^ n828 ;
  assign n8933 = n828 ^ n442 ;
  assign n8934 = n8933 ^ n828 ;
  assign n8935 = n8932 & ~n8934 ;
  assign n8936 = n8935 ^ n828 ;
  assign n8937 = ~n348 & n8936 ;
  assign n8938 = n8937 ^ n828 ;
  assign n8939 = n58 & n8938 ;
  assign n8940 = ~n8930 & ~n8939 ;
  assign n8941 = ~n8929 & n8940 ;
  assign n8942 = n3960 & ~n8941 ;
  assign n8943 = ~n4627 & ~n6492 ;
  assign n8944 = ~n2036 & ~n3030 ;
  assign n8945 = ~n8943 & ~n8944 ;
  assign n8946 = n364 & n1960 ;
  assign n8947 = x2 & n2271 ;
  assign n8948 = ~n28 & n8947 ;
  assign n8949 = n56 & n8948 ;
  assign n8950 = ~n8946 & ~n8949 ;
  assign n8951 = ~n8945 & n8950 ;
  assign n8952 = ~n1327 & ~n2036 ;
  assign n8953 = n328 & n1377 ;
  assign n8954 = ~x1 & ~n3019 ;
  assign n8955 = n6448 & n8954 ;
  assign n8956 = n929 & n8955 ;
  assign n8957 = ~n8953 & ~n8956 ;
  assign n8958 = n8952 & ~n8957 ;
  assign n8959 = ~x15 & n8958 ;
  assign n8960 = n8951 & ~n8959 ;
  assign n8961 = ~n8942 & n8960 ;
  assign n8962 = ~n8928 & ~n8961 ;
  assign n8963 = n263 & n1422 ;
  assign n8964 = n2027 & n8963 ;
  assign n8965 = n3777 & n5025 ;
  assign n8966 = ~n8964 & ~n8965 ;
  assign n8967 = n318 & n471 ;
  assign n8968 = ~n2904 & ~n8967 ;
  assign n8969 = n8968 ^ x2 ;
  assign n8970 = n8969 ^ n8968 ;
  assign n8971 = n8968 ^ n5277 ;
  assign n8972 = n8971 ^ n8968 ;
  assign n8973 = n8970 & n8972 ;
  assign n8974 = n8973 ^ n8968 ;
  assign n8975 = ~x0 & ~n8974 ;
  assign n8976 = n8975 ^ n8968 ;
  assign n8977 = n4829 & ~n8976 ;
  assign n8978 = n691 & ~n8968 ;
  assign n8979 = n1124 & n6562 ;
  assign n8980 = n55 & n784 ;
  assign n8981 = n787 & n8980 ;
  assign n8982 = ~n8979 & ~n8981 ;
  assign n8983 = n8982 ^ x14 ;
  assign n8984 = n8983 ^ n8982 ;
  assign n8985 = n8984 ^ n8978 ;
  assign n8986 = n8308 ^ n262 ;
  assign n8987 = n8986 ^ x0 ;
  assign n8994 = n8987 ^ n8986 ;
  assign n8988 = n8987 ^ n4942 ;
  assign n8989 = n8988 ^ n8986 ;
  assign n8990 = n8987 ^ n8308 ;
  assign n8991 = n8990 ^ n4942 ;
  assign n8992 = n8991 ^ n8989 ;
  assign n8993 = n8989 & ~n8992 ;
  assign n8995 = n8994 ^ n8993 ;
  assign n8996 = n8995 ^ n8989 ;
  assign n8997 = n8986 ^ n2477 ;
  assign n8998 = n8993 ^ n8989 ;
  assign n8999 = ~n8997 & n8998 ;
  assign n9000 = n8999 ^ n8986 ;
  assign n9001 = ~n8996 & n9000 ;
  assign n9002 = n9001 ^ n8986 ;
  assign n9003 = n9002 ^ n262 ;
  assign n9004 = n9003 ^ n8986 ;
  assign n9005 = n9004 ^ x1 ;
  assign n9006 = x1 & n9005 ;
  assign n9007 = n9006 ^ n8982 ;
  assign n9008 = n9007 ^ x1 ;
  assign n9009 = n8985 & ~n9008 ;
  assign n9010 = n9009 ^ n9006 ;
  assign n9011 = n9010 ^ x1 ;
  assign n9012 = ~n8978 & n9011 ;
  assign n9013 = n9012 ^ n8978 ;
  assign n9014 = ~n8977 & ~n9013 ;
  assign n9015 = x15 & ~n9014 ;
  assign n9016 = ~n1680 & ~n8980 ;
  assign n9017 = ~x0 & ~n9016 ;
  assign n9018 = ~x10 & n69 ;
  assign n9019 = ~n9017 & ~n9018 ;
  assign n9020 = n623 & ~n9019 ;
  assign n9021 = ~n9015 & ~n9020 ;
  assign n9022 = ~n8966 & ~n9021 ;
  assign n9023 = ~n8962 & ~n9022 ;
  assign n9024 = n66 & n1214 ;
  assign n9025 = n264 & n9024 ;
  assign n9026 = n266 & n5143 ;
  assign n9027 = ~n9025 & ~n9026 ;
  assign n9028 = n2612 & n2848 ;
  assign n9029 = ~n3907 & ~n9028 ;
  assign n9030 = ~n414 & ~n623 ;
  assign n9031 = ~n9029 & ~n9030 ;
  assign n9032 = ~x4 & n9031 ;
  assign n9033 = n1876 & n4470 ;
  assign n9034 = ~n3106 & ~n3894 ;
  assign n9035 = n9033 & n9034 ;
  assign n9036 = ~n2591 & ~n3960 ;
  assign n9037 = n9035 & n9036 ;
  assign n9038 = n2612 & n4730 ;
  assign n9039 = n3467 & n9038 ;
  assign n9040 = ~n9037 & ~n9039 ;
  assign n9041 = ~n9032 & n9040 ;
  assign n9042 = ~n9027 & ~n9041 ;
  assign n9043 = n2154 & n4769 ;
  assign n9044 = n18 & n5968 ;
  assign n9045 = ~n5231 & n9044 ;
  assign n9046 = ~n9043 & ~n9045 ;
  assign n9047 = ~n3803 & ~n9046 ;
  assign n9048 = n7594 & n8900 ;
  assign n9049 = n18 & n1977 ;
  assign n9050 = n8899 & n9049 ;
  assign n9051 = ~n9048 & ~n9050 ;
  assign n9052 = x9 ^ x8 ;
  assign n9053 = n9052 ^ n1228 ;
  assign n9054 = n718 ^ n76 ;
  assign n9055 = x2 & ~n9054 ;
  assign n9056 = n9055 ^ n76 ;
  assign n9057 = ~n9053 & n9056 ;
  assign n9058 = n9057 ^ n9055 ;
  assign n9059 = n9058 ^ n76 ;
  assign n9060 = n9059 ^ x2 ;
  assign n9061 = n9052 & n9060 ;
  assign n9062 = n2528 & n9061 ;
  assign n9063 = x12 & n9062 ;
  assign n9064 = n9051 & ~n9063 ;
  assign n9065 = ~n9047 & n9064 ;
  assign n9066 = n345 & ~n9065 ;
  assign n9067 = n104 & n8283 ;
  assign n9068 = n1427 & n8341 ;
  assign n9069 = n739 & n1954 ;
  assign n9070 = n262 & n9069 ;
  assign n9071 = ~n9068 & ~n9070 ;
  assign n9072 = n26 & n4954 ;
  assign n9073 = n9071 & ~n9072 ;
  assign n9074 = n9067 & ~n9073 ;
  assign n9075 = x8 & n9074 ;
  assign n9076 = ~n9066 & ~n9075 ;
  assign n9077 = n1050 & ~n9076 ;
  assign n9078 = ~n9042 & ~n9077 ;
  assign n9079 = n9023 & n9078 ;
  assign n9080 = n8924 & n9079 ;
  assign n9081 = n69 & n302 ;
  assign n9082 = n4632 & n9081 ;
  assign n9083 = x15 & n795 ;
  assign n9084 = n8341 & n9083 ;
  assign n9085 = n739 & n4350 ;
  assign n9086 = ~n1996 & ~n9085 ;
  assign n9087 = ~n741 & ~n9086 ;
  assign n9088 = ~n9084 & ~n9087 ;
  assign n9089 = x3 & ~n9088 ;
  assign n9090 = n4350 & n7646 ;
  assign n9091 = ~x2 & n9090 ;
  assign n9092 = ~n9089 & ~n9091 ;
  assign n9093 = n265 & ~n9092 ;
  assign n9094 = n33 & n2034 ;
  assign n9095 = n274 & n9094 ;
  assign n9096 = ~n9093 & ~n9095 ;
  assign n9097 = x14 & ~n9096 ;
  assign n9098 = n69 & n2033 ;
  assign n9099 = n1626 & n2031 ;
  assign n9100 = ~n9098 & ~n9099 ;
  assign n9101 = ~n9097 & n9100 ;
  assign n9102 = ~n3960 & ~n9101 ;
  assign n9103 = ~n9082 & ~n9102 ;
  assign n9104 = n8703 & ~n9103 ;
  assign n9105 = ~n267 & n1606 ;
  assign n9106 = n2033 & n3686 ;
  assign n9107 = ~n9105 & ~n9106 ;
  assign n9108 = n524 & ~n9107 ;
  assign n9109 = n366 & n740 ;
  assign n9110 = n246 & n9109 ;
  assign n9111 = n1198 & n9110 ;
  assign n9112 = ~n9108 & ~n9111 ;
  assign n9113 = n1422 & ~n9112 ;
  assign n9114 = x8 & n2806 ;
  assign n9115 = ~x3 & n7217 ;
  assign n9116 = n9114 & n9115 ;
  assign n9117 = n2300 & n3257 ;
  assign n9118 = n9116 & n9117 ;
  assign n9119 = ~n9113 & ~n9118 ;
  assign n9120 = n700 & ~n9119 ;
  assign n9121 = n328 & n1954 ;
  assign n9122 = n1014 & n8017 ;
  assign n9123 = n5164 & n8018 ;
  assign n9124 = ~n9122 & ~n9123 ;
  assign n9125 = n9121 & ~n9124 ;
  assign n9126 = ~n263 & ~n652 ;
  assign n9127 = n4146 & n8017 ;
  assign n9128 = n4145 & n8018 ;
  assign n9129 = ~n9127 & ~n9128 ;
  assign n9130 = ~n265 & ~n2991 ;
  assign n9131 = ~n9129 & ~n9130 ;
  assign n9132 = ~n9126 & n9131 ;
  assign n9133 = ~n9125 & ~n9132 ;
  assign n9134 = n679 & ~n9133 ;
  assign n9135 = ~n2035 & n2816 ;
  assign n9136 = n65 & n4222 ;
  assign n9137 = n4350 & n9136 ;
  assign n9138 = n9135 & n9137 ;
  assign n9139 = ~n9134 & ~n9138 ;
  assign n9140 = n265 & n2806 ;
  assign n9141 = n8309 & n9140 ;
  assign n9142 = n8308 & n8963 ;
  assign n9143 = ~n9141 & ~n9142 ;
  assign n9144 = ~n3960 & ~n9143 ;
  assign n9145 = ~n1511 & n9144 ;
  assign n9146 = ~x8 & n2806 ;
  assign n9147 = n691 & n1989 ;
  assign n9148 = n1427 & n9147 ;
  assign n9149 = n9146 & n9148 ;
  assign n9150 = ~n9145 & ~n9149 ;
  assign n9151 = n9139 & n9150 ;
  assign n9152 = ~n9120 & n9151 ;
  assign n9153 = ~n9104 & n9152 ;
  assign n9154 = n4832 & ~n9153 ;
  assign n9155 = n9080 & ~n9154 ;
  assign n9156 = ~n3172 & ~n3177 ;
  assign n9157 = n175 & n2608 ;
  assign n9158 = ~x4 & ~n2815 ;
  assign n9159 = ~n2910 & n9158 ;
  assign n9160 = ~n274 & n9159 ;
  assign n9161 = ~n9157 & ~n9160 ;
  assign n9162 = n3091 & ~n9161 ;
  assign n9163 = n8371 & n9162 ;
  assign n9164 = n26 & n2881 ;
  assign n9165 = n5530 & n9164 ;
  assign n9166 = n2637 & n9157 ;
  assign n9167 = n798 & n6923 ;
  assign n9168 = n2637 ^ n2480 ;
  assign n9169 = x4 & n9168 ;
  assign n9170 = n9169 ^ n2480 ;
  assign n9171 = n9167 & n9170 ;
  assign n9172 = ~n9166 & ~n9171 ;
  assign n9173 = n1464 & ~n9172 ;
  assign n9174 = ~n9165 & ~n9173 ;
  assign n9175 = x14 & ~n9174 ;
  assign n9176 = ~n9163 & ~n9175 ;
  assign n9177 = n9176 ^ x2 ;
  assign n9178 = n9177 ^ n2480 ;
  assign n9179 = n9178 ^ n9176 ;
  assign n9208 = n9179 ^ n9177 ;
  assign n9209 = n9208 ^ n9176 ;
  assign n9210 = n9209 ^ n9176 ;
  assign n9211 = n26 & n3960 ;
  assign n9212 = n224 ^ x6 ;
  assign n9213 = n224 ^ x8 ;
  assign n9214 = n9213 ^ x8 ;
  assign n9215 = n1906 ^ x8 ;
  assign n9216 = ~n9214 & ~n9215 ;
  assign n9217 = n9216 ^ x8 ;
  assign n9218 = n9212 & n9217 ;
  assign n9219 = n9218 ^ x6 ;
  assign n9220 = n9211 & n9219 ;
  assign n9221 = ~n2239 & ~n3288 ;
  assign n9222 = ~x6 & ~x8 ;
  assign n9223 = ~x0 & n168 ;
  assign n9224 = n9223 ^ n1464 ;
  assign n9225 = ~n9222 & n9224 ;
  assign n9226 = n9225 ^ n1464 ;
  assign n9227 = ~n274 & n9226 ;
  assign n9228 = ~n9221 & n9227 ;
  assign n9229 = x2 & ~n9228 ;
  assign n9230 = ~n9220 & n9229 ;
  assign n9231 = n9230 ^ n9177 ;
  assign n9232 = n9231 ^ n9177 ;
  assign n9233 = n9232 ^ n9176 ;
  assign n9234 = ~n9210 & n9233 ;
  assign n9180 = ~x8 & n7473 ;
  assign n9181 = ~n1270 & n1494 ;
  assign n9182 = n89 & n9181 ;
  assign n9183 = ~n9180 & n9182 ;
  assign n9186 = n2679 & n3960 ;
  assign n9187 = x5 & ~n7045 ;
  assign n9188 = x0 & ~n2711 ;
  assign n9189 = ~n9187 & n9188 ;
  assign n9190 = ~n9186 & ~n9189 ;
  assign n9191 = n3287 & ~n9190 ;
  assign n9184 = n1909 & n7899 ;
  assign n9185 = n68 & n9184 ;
  assign n9192 = n9191 ^ n9185 ;
  assign n9193 = n9192 ^ n9191 ;
  assign n9194 = x8 & n2599 ;
  assign n9195 = ~n5239 & ~n9187 ;
  assign n9196 = n9194 & n9195 ;
  assign n9197 = n9196 ^ n9191 ;
  assign n9198 = n9197 ^ n9191 ;
  assign n9199 = ~n9193 & ~n9198 ;
  assign n9200 = n9199 ^ n9191 ;
  assign n9201 = x4 & ~n9200 ;
  assign n9202 = n9201 ^ n9191 ;
  assign n9203 = ~n9183 & ~n9202 ;
  assign n9204 = n9203 ^ n9177 ;
  assign n9205 = n9204 ^ n9179 ;
  assign n9206 = n9205 ^ n9176 ;
  assign n9207 = n9179 & ~n9206 ;
  assign n9235 = n9234 ^ n9207 ;
  assign n9236 = n9235 ^ n9179 ;
  assign n9237 = n9207 ^ n9176 ;
  assign n9238 = n9237 ^ n9209 ;
  assign n9239 = ~n9176 & ~n9238 ;
  assign n9240 = n9239 ^ n9207 ;
  assign n9241 = n9236 & n9240 ;
  assign n9242 = n9241 ^ n9234 ;
  assign n9243 = n9242 ^ n9239 ;
  assign n9244 = n9243 ^ n9179 ;
  assign n9245 = n9244 ^ n9176 ;
  assign n9246 = n9245 ^ n9209 ;
  assign n9247 = n9246 ^ x2 ;
  assign n9248 = x1 & n9247 ;
  assign n9249 = n3967 & n7045 ;
  assign n9250 = n1514 & n1538 ;
  assign n9251 = n9249 & n9250 ;
  assign n9252 = x4 & n2480 ;
  assign n9253 = ~n8217 & ~n9252 ;
  assign n9254 = n20 & ~n9253 ;
  assign n9255 = n60 & n352 ;
  assign n9256 = ~n40 & n2568 ;
  assign n9257 = ~n9255 & ~n9256 ;
  assign n9258 = n2637 & ~n9257 ;
  assign n9259 = ~n8725 & n8916 ;
  assign n9260 = ~n60 & n2480 ;
  assign n9261 = ~n9259 & n9260 ;
  assign n9262 = ~n9258 & ~n9261 ;
  assign n9263 = ~x15 & ~n9262 ;
  assign n9264 = n58 & ~n3288 ;
  assign n9265 = n9170 & n9264 ;
  assign n9266 = ~n9263 & ~n9265 ;
  assign n9267 = ~n9254 & n9266 ;
  assign n9268 = n1464 & ~n9267 ;
  assign n9269 = n1499 & n6824 ;
  assign n9270 = n714 & n9269 ;
  assign n9271 = ~n9268 & ~n9270 ;
  assign n9272 = ~n9251 & n9271 ;
  assign n9273 = ~n3494 & ~n9272 ;
  assign n9274 = x7 & ~x15 ;
  assign n9275 = ~n4166 & ~n9274 ;
  assign n9276 = n4955 & ~n9275 ;
  assign n9277 = x7 & n786 ;
  assign n9278 = ~n9276 & ~n9277 ;
  assign n9279 = n3835 & ~n9278 ;
  assign n9280 = n1048 & n3960 ;
  assign n9281 = ~x6 & n9280 ;
  assign n9282 = n2581 & n2686 ;
  assign n9283 = x14 & n9282 ;
  assign n9284 = ~n9281 & ~n9283 ;
  assign n9285 = ~n9279 & n9284 ;
  assign n9286 = x0 & ~n9285 ;
  assign n9287 = ~x15 & n60 ;
  assign n9288 = n9282 & n9287 ;
  assign n9289 = ~n9286 & ~n9288 ;
  assign n9290 = n352 & ~n9289 ;
  assign n9291 = n928 & n2701 ;
  assign n9292 = n7045 & n9291 ;
  assign n9293 = n8853 & n9292 ;
  assign n9294 = x8 & ~n3729 ;
  assign n9295 = ~x6 & ~n9274 ;
  assign n9296 = n9294 & ~n9295 ;
  assign n9297 = n9255 & n9296 ;
  assign n9298 = ~n9293 & ~n9297 ;
  assign n9299 = ~n9290 & n9298 ;
  assign n9300 = n2711 & ~n9299 ;
  assign n9301 = n9109 & n9184 ;
  assign n9302 = ~n300 & ~n1623 ;
  assign n9303 = ~x0 & ~n9302 ;
  assign n9304 = n574 & ~n9303 ;
  assign n9305 = n3960 & ~n9304 ;
  assign n9306 = ~n652 & ~n6097 ;
  assign n9307 = ~n312 & ~n366 ;
  assign n9308 = n572 & n9307 ;
  assign n9309 = ~n9306 & n9308 ;
  assign n9310 = ~n9305 & ~n9309 ;
  assign n9311 = n42 & n196 ;
  assign n9312 = n9311 ^ n9287 ;
  assign n9313 = n9311 ^ n9250 ;
  assign n9314 = n9313 ^ n9250 ;
  assign n9315 = n9250 ^ n2282 ;
  assign n9316 = n9314 & ~n9315 ;
  assign n9317 = n9316 ^ n9250 ;
  assign n9318 = n9312 & ~n9317 ;
  assign n9319 = n9318 ^ n9287 ;
  assign n9320 = n9310 & ~n9319 ;
  assign n9321 = n3287 & ~n9320 ;
  assign n9322 = ~n9301 & ~n9321 ;
  assign n9323 = ~n3729 & ~n9322 ;
  assign n9324 = n25 & n249 ;
  assign n9325 = n213 & n9324 ;
  assign n9326 = ~n44 & ~n7129 ;
  assign n9327 = n68 & n9326 ;
  assign n9328 = n9327 ^ x5 ;
  assign n9329 = n9328 ^ n9327 ;
  assign n9330 = n9329 ^ x15 ;
  assign n9331 = n7129 ^ n249 ;
  assign n9332 = x2 & ~n9331 ;
  assign n9333 = n9332 ^ n249 ;
  assign n9334 = n25 & n9333 ;
  assign n9335 = ~n250 & ~n3010 ;
  assign n9336 = n224 & ~n9335 ;
  assign n9337 = n9336 ^ n9334 ;
  assign n9338 = ~n9334 & n9337 ;
  assign n9339 = n9338 ^ n9327 ;
  assign n9340 = n9339 ^ n9334 ;
  assign n9341 = n9330 & n9340 ;
  assign n9342 = n9341 ^ n9338 ;
  assign n9343 = n9342 ^ n9334 ;
  assign n9344 = ~x15 & ~n9343 ;
  assign n9345 = n9344 ^ x15 ;
  assign n9346 = ~n9325 & n9345 ;
  assign n9347 = n3165 & n3835 ;
  assign n9348 = ~n9282 & ~n9347 ;
  assign n9349 = ~n9346 & ~n9348 ;
  assign n9350 = ~n9323 & ~n9349 ;
  assign n9351 = ~n9300 & n9350 ;
  assign n9352 = ~n9273 & n9351 ;
  assign n9353 = n9248 & n9352 ;
  assign n9354 = n3960 & n9294 ;
  assign n9355 = ~n175 & n858 ;
  assign n9356 = ~n456 & n5785 ;
  assign n9357 = ~n9355 & ~n9356 ;
  assign n9358 = x14 & ~n9357 ;
  assign n9359 = ~n9354 & ~n9358 ;
  assign n9360 = n168 & ~n9359 ;
  assign n9361 = x7 & n8095 ;
  assign n9362 = ~n9280 & ~n9361 ;
  assign n9363 = ~n9294 & n9362 ;
  assign n9364 = n2679 & ~n9363 ;
  assign n9365 = ~n9360 & ~n9364 ;
  assign n9366 = x6 & ~n9365 ;
  assign n9367 = ~x5 & ~n633 ;
  assign n9368 = ~n1217 & n9367 ;
  assign n9369 = ~x3 & ~n9368 ;
  assign n9370 = ~n561 & n6923 ;
  assign n9371 = ~n3091 & n9370 ;
  assign n9372 = n2508 & ~n5908 ;
  assign n9373 = ~n68 & ~n1515 ;
  assign n9374 = ~n9372 & ~n9373 ;
  assign n9375 = ~n314 & ~n373 ;
  assign n9376 = ~n2480 & n9375 ;
  assign n9377 = n9374 & n9376 ;
  assign n9378 = n9371 & n9377 ;
  assign n9379 = ~n9369 & n9378 ;
  assign n9380 = ~n9366 & ~n9379 ;
  assign n9381 = ~n8645 & ~n9380 ;
  assign n9382 = n3967 ^ n2711 ;
  assign n9383 = n884 & n1565 ;
  assign n9384 = n9383 ^ n3967 ;
  assign n9385 = n9384 ^ n9383 ;
  assign n9386 = n9385 ^ n9382 ;
  assign n9387 = n319 ^ n314 ;
  assign n9388 = n314 & n9387 ;
  assign n9389 = n9388 ^ n9383 ;
  assign n9390 = n9389 ^ n314 ;
  assign n9391 = n9386 & ~n9390 ;
  assign n9392 = n9391 ^ n9388 ;
  assign n9393 = n9392 ^ n314 ;
  assign n9394 = n9382 & n9393 ;
  assign n9395 = n9394 ^ n2711 ;
  assign n9396 = n352 & n9395 ;
  assign n9397 = x2 & n3728 ;
  assign n9398 = n8620 & n9397 ;
  assign n9399 = ~n9250 & ~n9311 ;
  assign n9400 = ~x14 & n3967 ;
  assign n9401 = ~n9383 & ~n9400 ;
  assign n9402 = ~n9399 & ~n9401 ;
  assign n9403 = x5 & n8634 ;
  assign n9404 = n9403 ^ n314 ;
  assign n9405 = n8915 & n9404 ;
  assign n9406 = n2480 & n9405 ;
  assign n9407 = ~n9402 & ~n9406 ;
  assign n9408 = ~n9398 & n9407 ;
  assign n9409 = ~x15 & ~n9408 ;
  assign n9410 = ~n9396 & ~n9409 ;
  assign n9411 = ~n3494 & ~n9410 ;
  assign n9412 = n1909 & n8652 ;
  assign n9413 = n111 & n8684 ;
  assign n9414 = ~n9412 & ~n9413 ;
  assign n9415 = n2747 & ~n9414 ;
  assign n9416 = n6862 & n7029 ;
  assign n9417 = n778 & n9416 ;
  assign n9418 = ~n9415 & ~n9417 ;
  assign n9419 = n6824 & ~n9418 ;
  assign n9420 = ~x7 & n2562 ;
  assign n9421 = n277 & n556 ;
  assign n9422 = n9420 & n9421 ;
  assign n9423 = x0 & n7045 ;
  assign n9424 = x4 ^ x2 ;
  assign n9425 = n282 ^ x4 ;
  assign n9426 = n9425 ^ n282 ;
  assign n9427 = n1515 ^ n282 ;
  assign n9428 = ~n9426 & n9427 ;
  assign n9429 = n9428 ^ n282 ;
  assign n9430 = ~n9424 & n9429 ;
  assign n9431 = n9423 & n9430 ;
  assign n9432 = n2684 & n9431 ;
  assign n9433 = ~n9422 & ~n9432 ;
  assign n9434 = ~n9419 & n9433 ;
  assign n9435 = n2711 & ~n9434 ;
  assign n9436 = n1422 & n2033 ;
  assign n9437 = n65 & n9436 ;
  assign n9438 = n264 & n8017 ;
  assign n9439 = ~n9437 & ~n9438 ;
  assign n9440 = x15 & ~n4170 ;
  assign n9441 = ~n9439 & n9440 ;
  assign n9442 = x14 ^ x9 ;
  assign n9443 = n9114 ^ x14 ;
  assign n9444 = n9443 ^ n9114 ;
  assign n9445 = n6824 & n9222 ;
  assign n9446 = n9445 ^ n9114 ;
  assign n9447 = ~n9444 & n9446 ;
  assign n9448 = n9447 ^ n9114 ;
  assign n9449 = ~n9442 & n9448 ;
  assign n9450 = ~n9399 & n9449 ;
  assign n9451 = x0 & n9450 ;
  assign n9452 = ~n9441 & ~n9451 ;
  assign n9453 = n9348 ^ n2282 ;
  assign n9454 = n1994 ^ x3 ;
  assign n9455 = n9454 ^ n1994 ;
  assign n9456 = n1994 ^ n1606 ;
  assign n9457 = n9456 ^ n1994 ;
  assign n9458 = ~n9455 & n9457 ;
  assign n9459 = n9458 ^ n1994 ;
  assign n9460 = ~x2 & n9459 ;
  assign n9461 = n9460 ^ n1994 ;
  assign n9462 = n3960 & n9461 ;
  assign n9463 = n9462 ^ n9453 ;
  assign n9464 = n9463 ^ n9348 ;
  assign n9465 = n9464 ^ n9463 ;
  assign n9466 = n1538 & n2684 ;
  assign n9467 = n1513 & n9466 ;
  assign n9468 = n1516 & n9164 ;
  assign n9469 = ~n9467 & ~n9468 ;
  assign n9470 = n9469 ^ n9463 ;
  assign n9471 = n9470 ^ n9453 ;
  assign n9472 = ~n9465 & n9471 ;
  assign n9473 = n9472 ^ n9469 ;
  assign n9474 = n712 & n9307 ;
  assign n9475 = ~n9250 & ~n9474 ;
  assign n9476 = n9469 & n9475 ;
  assign n9477 = n9476 ^ n9453 ;
  assign n9478 = n9473 & n9477 ;
  assign n9479 = n9478 ^ n9476 ;
  assign n9480 = n9453 & n9479 ;
  assign n9481 = n9480 ^ n9472 ;
  assign n9482 = n9481 ^ n2282 ;
  assign n9483 = n9482 ^ n9469 ;
  assign n9484 = n9452 & ~n9483 ;
  assign n9485 = n34 & n263 ;
  assign n9486 = ~n2033 & ~n9485 ;
  assign n9487 = x3 & n363 ;
  assign n9488 = n3427 & n9487 ;
  assign n9489 = ~n9486 & n9488 ;
  assign n9490 = n844 & n6562 ;
  assign n9491 = n9294 & n9490 ;
  assign n9492 = x4 & ~n3494 ;
  assign n9493 = n25 & n363 ;
  assign n9494 = n526 & n9493 ;
  assign n9495 = n9492 & n9494 ;
  assign n9496 = ~n9491 & ~n9495 ;
  assign n9497 = ~n9489 & n9496 ;
  assign n9498 = n9484 & n9497 ;
  assign n9499 = ~n9435 & n9498 ;
  assign n9500 = ~n9411 & n9499 ;
  assign n9501 = ~x4 & n7022 ;
  assign n9502 = n80 & n9501 ;
  assign n9503 = n720 & n9502 ;
  assign n9504 = n3287 & n8725 ;
  assign n9505 = n4955 & n8652 ;
  assign n9506 = ~n9504 & ~n9505 ;
  assign n9507 = n2679 & ~n9506 ;
  assign n9508 = n556 & n3894 ;
  assign n9509 = n106 & n3106 ;
  assign n9510 = ~n9508 & ~n9509 ;
  assign n9511 = n1514 & n2282 ;
  assign n9512 = ~n9510 & n9511 ;
  assign n9513 = ~n9507 & ~n9512 ;
  assign n9514 = ~n9503 & n9513 ;
  assign n9515 = ~n3729 & ~n9514 ;
  assign n9516 = ~n9348 & ~n9399 ;
  assign n9517 = n9469 & ~n9516 ;
  assign n9518 = ~n4170 & ~n9517 ;
  assign n9519 = ~n9515 & ~n9518 ;
  assign n9520 = ~x15 & ~n9519 ;
  assign n9521 = ~x1 & ~n9520 ;
  assign n9522 = n9500 & n9521 ;
  assign n9523 = ~n9381 & n9522 ;
  assign n9524 = ~n9353 & ~n9523 ;
  assign n9525 = ~n8963 & ~n9140 ;
  assign n9526 = n66 & n313 ;
  assign n9527 = ~x4 & ~n7045 ;
  assign n9528 = n66 & ~n9527 ;
  assign n9529 = ~n6924 & ~n9528 ;
  assign n9530 = ~x3 & ~n9529 ;
  assign n9531 = n66 & n1494 ;
  assign n9532 = ~n8551 & ~n9531 ;
  assign n9533 = n1270 & ~n9532 ;
  assign n9534 = n1494 & n1954 ;
  assign n9535 = n3960 & n9534 ;
  assign n9536 = ~n9533 & ~n9535 ;
  assign n9537 = ~n9530 & n9536 ;
  assign n9538 = ~n9526 & n9537 ;
  assign n9539 = n213 & ~n9538 ;
  assign n9540 = n5507 & n7052 ;
  assign n9541 = n9527 ^ x15 ;
  assign n9542 = n9541 ^ n9527 ;
  assign n9543 = n9527 ^ n7129 ;
  assign n9544 = n9543 ^ n9527 ;
  assign n9545 = n9542 & ~n9544 ;
  assign n9546 = n9545 ^ n9527 ;
  assign n9547 = x1 & ~n9546 ;
  assign n9548 = n9547 ^ n9527 ;
  assign n9549 = n68 & ~n9548 ;
  assign n9550 = n1581 & n8829 ;
  assign n9551 = x0 & n9550 ;
  assign n9552 = ~n9549 & ~n9551 ;
  assign n9553 = ~n9540 & n9552 ;
  assign n9554 = n180 & ~n9553 ;
  assign n9555 = x15 ^ x2 ;
  assign n9556 = n513 ^ n376 ;
  assign n9557 = n376 ^ x15 ;
  assign n9558 = n9557 ^ n376 ;
  assign n9559 = n9556 & ~n9558 ;
  assign n9560 = n9559 ^ n376 ;
  assign n9561 = n9555 & n9560 ;
  assign n9562 = n2568 & n9561 ;
  assign n9563 = x15 & n60 ;
  assign n9564 = n376 & n9563 ;
  assign n9565 = ~n9255 & ~n9564 ;
  assign n9566 = n5976 & n8863 ;
  assign n9567 = n9565 & ~n9566 ;
  assign n9568 = ~n9562 & n9567 ;
  assign n9569 = n196 & ~n9568 ;
  assign n9570 = ~n9554 & ~n9569 ;
  assign n9571 = ~n9539 & n9570 ;
  assign n9572 = ~n9525 & ~n9571 ;
  assign n9573 = x0 & ~n2508 ;
  assign n9574 = ~n858 & n9573 ;
  assign n9575 = ~n9249 & ~n9574 ;
  assign n9576 = n3186 & ~n9575 ;
  assign n9577 = ~n1270 & ~n2480 ;
  assign n9578 = ~n2637 & ~n9577 ;
  assign n9579 = n9194 & n9578 ;
  assign n9580 = ~n7029 & ~n7045 ;
  assign n9581 = ~n2815 & n6893 ;
  assign n9582 = ~n9580 & n9581 ;
  assign n9583 = ~n9579 & ~n9582 ;
  assign n9584 = ~n9576 & n9583 ;
  assign n9585 = ~x1 & ~n9584 ;
  assign n9586 = n434 & n4014 ;
  assign n9587 = ~n786 & n9586 ;
  assign n9588 = ~n9180 & n9587 ;
  assign n9589 = x15 & n9588 ;
  assign n9590 = ~n3287 & n9589 ;
  assign n9591 = ~n9585 & ~n9590 ;
  assign n9592 = n1626 & ~n9591 ;
  assign n9593 = ~n9572 & ~n9592 ;
  assign n9594 = ~n9524 & n9593 ;
  assign n9595 = ~n9156 & ~n9594 ;
  assign n9596 = n9155 & ~n9595 ;
  assign n9597 = n8852 & n9596 ;
  assign n9598 = ~n9164 & ~n9466 ;
  assign n9599 = ~n1014 & ~n5164 ;
  assign n9600 = ~n2326 & ~n5238 ;
  assign n9601 = n32 & n2282 ;
  assign n9602 = ~n863 & n9601 ;
  assign n9603 = n9600 & n9602 ;
  assign n9604 = x13 & n690 ;
  assign n9605 = n1113 & n5976 ;
  assign n9606 = ~n28 & n9563 ;
  assign n9607 = ~n9605 & ~n9606 ;
  assign n9608 = ~n9604 & n9607 ;
  assign n9609 = n65 & ~n9608 ;
  assign n9610 = n828 & ~n4346 ;
  assign n9611 = ~x12 & ~n80 ;
  assign n9612 = ~n3003 & ~n9611 ;
  assign n9613 = ~n9610 & n9612 ;
  assign n9614 = ~n9609 & ~n9613 ;
  assign n9615 = ~n9603 & n9614 ;
  assign n9616 = ~n3019 & ~n8162 ;
  assign n9617 = n66 & n9616 ;
  assign n9618 = ~n3164 & ~n9617 ;
  assign n9619 = x15 & ~n9618 ;
  assign n9620 = n1954 & n8808 ;
  assign n9621 = ~n4421 & ~n9121 ;
  assign n9622 = ~n9620 & n9621 ;
  assign n9623 = ~n310 & ~n6484 ;
  assign n9624 = x13 & ~n9623 ;
  assign n9625 = n20 & ~n5239 ;
  assign n9626 = ~n19 & ~n700 ;
  assign n9627 = ~n38 & ~n741 ;
  assign n9628 = ~n9626 & n9627 ;
  assign n9629 = ~n9625 & ~n9628 ;
  assign n9630 = ~n9624 & n9629 ;
  assign n9631 = x12 & n9630 ;
  assign n9632 = n9622 & n9631 ;
  assign n9633 = ~n9619 & n9632 ;
  assign n9634 = ~n9615 & ~n9633 ;
  assign n9635 = x1 & n6490 ;
  assign n9636 = ~n9634 & ~n9635 ;
  assign n9637 = ~n9599 & ~n9636 ;
  assign n9638 = ~n673 & ~n1270 ;
  assign n9639 = n1514 & n9638 ;
  assign n9640 = ~n177 & ~n9639 ;
  assign n9641 = n4684 & ~n9640 ;
  assign n9642 = ~n163 & ~n8829 ;
  assign n9643 = n9642 ^ x2 ;
  assign n9644 = n9643 ^ n9642 ;
  assign n9645 = n9644 ^ x11 ;
  assign n9646 = ~n328 & ~n863 ;
  assign n9647 = n9646 ^ n314 ;
  assign n9648 = ~n314 & n9647 ;
  assign n9649 = n9648 ^ n9642 ;
  assign n9650 = n9649 ^ n314 ;
  assign n9651 = n9645 & n9650 ;
  assign n9652 = n9651 ^ n9648 ;
  assign n9653 = n9652 ^ n314 ;
  assign n9654 = ~x11 & ~n9653 ;
  assign n9655 = n396 & n9654 ;
  assign n9656 = ~x14 & ~n8808 ;
  assign n9657 = n2402 & ~n9656 ;
  assign n9658 = ~n9655 & ~n9657 ;
  assign n9659 = ~n9641 & n9658 ;
  assign n9660 = n639 & ~n1270 ;
  assign n9661 = ~n7841 & ~n9660 ;
  assign n9662 = n55 & ~n9661 ;
  assign n9663 = n702 & n1290 ;
  assign n9664 = ~n9662 & ~n9663 ;
  assign n9665 = x13 & ~n9664 ;
  assign n9666 = n9659 & ~n9665 ;
  assign n9667 = n1682 & ~n9666 ;
  assign n9668 = ~x15 & n718 ;
  assign n9669 = n8341 & n9668 ;
  assign n9670 = n306 & n5968 ;
  assign n9671 = ~n1645 & ~n9670 ;
  assign n9672 = ~n9669 & n9671 ;
  assign n9673 = ~x3 & ~n9672 ;
  assign n9674 = n6484 & n9604 ;
  assign n9675 = ~n9673 & ~n9674 ;
  assign n9676 = n346 & ~n9675 ;
  assign n9677 = ~n163 & ~n442 ;
  assign n9678 = ~n3992 & n9677 ;
  assign n9679 = n66 & ~n5998 ;
  assign n9680 = ~n110 & n9679 ;
  assign n9681 = ~n9678 & ~n9680 ;
  assign n9682 = n639 & ~n9681 ;
  assign n9683 = ~n702 & ~n4992 ;
  assign n9684 = n518 & ~n9683 ;
  assign n9685 = ~n126 & ~n4350 ;
  assign n9686 = n346 & n6562 ;
  assign n9687 = n9685 & n9686 ;
  assign n9688 = ~n9684 & ~n9687 ;
  assign n9689 = ~n9682 & n9688 ;
  assign n9690 = n1282 & ~n9689 ;
  assign n9691 = ~n9676 & ~n9690 ;
  assign n9692 = n327 & n8829 ;
  assign n9693 = n1090 & n3960 ;
  assign n9694 = ~n6491 & ~n8805 ;
  assign n9695 = ~n9693 & ~n9694 ;
  assign n9696 = ~n9692 & n9695 ;
  assign n9697 = n2738 & ~n9696 ;
  assign n9698 = n9697 ^ x12 ;
  assign n9699 = n9698 ^ n9697 ;
  assign n9700 = n56 & ~n673 ;
  assign n9701 = ~n110 & ~n126 ;
  assign n9702 = ~n9700 & n9701 ;
  assign n9703 = n757 & n762 ;
  assign n9704 = ~n9702 & n9703 ;
  assign n9705 = ~n6097 & n9642 ;
  assign n9706 = n978 & ~n9705 ;
  assign n9707 = n396 & n9706 ;
  assign n9708 = ~x2 & n9707 ;
  assign n9709 = ~n1227 & n1966 ;
  assign n9710 = x15 & n110 ;
  assign n9711 = ~x14 & n68 ;
  assign n9712 = ~n9710 & ~n9711 ;
  assign n9713 = n7386 & ~n9712 ;
  assign n9714 = ~n9709 & ~n9713 ;
  assign n9715 = n74 & ~n9714 ;
  assign n9716 = ~n9708 & ~n9715 ;
  assign n9717 = ~n9704 & n9716 ;
  assign n9718 = n9717 ^ n9697 ;
  assign n9719 = n9699 & ~n9718 ;
  assign n9720 = n9719 ^ n9697 ;
  assign n9721 = n9691 & ~n9720 ;
  assign n9722 = ~n9667 & n9721 ;
  assign n9723 = ~n467 & ~n9722 ;
  assign n9724 = ~n9637 & ~n9723 ;
  assign n9725 = n3019 ^ n2607 ;
  assign n9726 = n9725 ^ x8 ;
  assign n9733 = n9726 ^ n9725 ;
  assign n9727 = n9726 ^ n198 ;
  assign n9728 = n9727 ^ n9725 ;
  assign n9729 = n9726 ^ n3019 ;
  assign n9730 = n9729 ^ n198 ;
  assign n9731 = n9730 ^ n9728 ;
  assign n9732 = n9728 & n9731 ;
  assign n9734 = n9733 ^ n9732 ;
  assign n9735 = n9734 ^ n9728 ;
  assign n9736 = n9725 ^ n1270 ;
  assign n9737 = n9732 ^ n9728 ;
  assign n9738 = n9736 & n9737 ;
  assign n9739 = n9738 ^ n9725 ;
  assign n9740 = ~n9735 & ~n9739 ;
  assign n9741 = n9740 ^ n9725 ;
  assign n9742 = n9741 ^ n2607 ;
  assign n9743 = n9742 ^ n9725 ;
  assign n9744 = n55 & ~n9743 ;
  assign n9745 = n65 & ~n4955 ;
  assign n9746 = ~n465 & ~n568 ;
  assign n9747 = n9745 & n9746 ;
  assign n9748 = ~x8 & n3960 ;
  assign n9749 = n946 & n9748 ;
  assign n9750 = ~n1003 & ~n9749 ;
  assign n9751 = n442 & ~n9750 ;
  assign n9752 = ~n9747 & ~n9751 ;
  assign n9753 = ~n9744 & n9752 ;
  assign n9754 = n5619 & ~n9753 ;
  assign n9755 = n453 & n4952 ;
  assign n9756 = n1146 & n9755 ;
  assign n9757 = ~n9754 & ~n9756 ;
  assign n9758 = ~n463 & ~n9749 ;
  assign n9759 = x13 & n8829 ;
  assign n9760 = ~n65 & ~n9759 ;
  assign n9761 = ~n9758 & ~n9760 ;
  assign n9762 = x8 ^ x3 ;
  assign n9763 = n946 ^ n784 ;
  assign n9764 = n784 ^ x8 ;
  assign n9765 = n9764 ^ n784 ;
  assign n9766 = n9763 & ~n9765 ;
  assign n9767 = n9766 ^ n784 ;
  assign n9768 = ~n9762 & n9767 ;
  assign n9769 = ~n673 & n9768 ;
  assign n9770 = ~n9761 & ~n9769 ;
  assign n9771 = n1742 & ~n9770 ;
  assign n9772 = n364 & n4952 ;
  assign n9773 = x1 & n7834 ;
  assign n9774 = n9772 & n9773 ;
  assign n9775 = n110 & n1003 ;
  assign n9776 = n2224 & ~n9656 ;
  assign n9777 = ~x3 & n9776 ;
  assign n9778 = ~n9775 & ~n9777 ;
  assign n9779 = n1382 & ~n9778 ;
  assign n9780 = ~n9774 & ~n9779 ;
  assign n9781 = ~n9771 & n9780 ;
  assign n9782 = n9781 ^ x0 ;
  assign n9783 = n9782 ^ n9781 ;
  assign n9784 = n9783 ^ n9757 ;
  assign n9785 = n141 & n1214 ;
  assign n9786 = ~n6097 & n9785 ;
  assign n9787 = n442 & ~n4098 ;
  assign n9788 = ~n76 & ~n4333 ;
  assign n9789 = ~n2338 & ~n9788 ;
  assign n9790 = ~x15 & n9789 ;
  assign n9791 = ~n9787 & ~n9790 ;
  assign n9792 = n1095 & ~n9791 ;
  assign n9793 = x3 & ~n5976 ;
  assign n9794 = ~n1349 & ~n1382 ;
  assign n9795 = n176 & ~n9794 ;
  assign n9796 = ~n9793 & n9795 ;
  assign n9797 = ~n9792 & ~n9796 ;
  assign n9798 = ~n9786 & n9797 ;
  assign n9799 = n9798 ^ n463 ;
  assign n9800 = n463 & ~n9799 ;
  assign n9801 = n9800 ^ n9781 ;
  assign n9802 = n9801 ^ n463 ;
  assign n9803 = ~n9784 & ~n9802 ;
  assign n9804 = n9803 ^ n9800 ;
  assign n9805 = n9804 ^ n463 ;
  assign n9806 = n9757 & n9805 ;
  assign n9807 = n9806 ^ n9757 ;
  assign n9808 = ~n555 & ~n9807 ;
  assign n9809 = n4350 & n5462 ;
  assign n9810 = n442 & ~n5698 ;
  assign n9811 = ~n4832 & n9810 ;
  assign n9812 = ~n9809 & ~n9811 ;
  assign n9813 = ~x8 & ~n9812 ;
  assign n9814 = ~n8440 & ~n9813 ;
  assign n9815 = ~x9 & n623 ;
  assign n9816 = ~n9814 & n9815 ;
  assign n9817 = ~x9 & n1667 ;
  assign n9818 = n965 & n4098 ;
  assign n9819 = n9817 & n9818 ;
  assign n9820 = ~n18 & n230 ;
  assign n9821 = n2356 & n9820 ;
  assign n9822 = ~n786 & ~n4955 ;
  assign n9823 = ~n1270 & n5656 ;
  assign n9824 = n9822 & n9823 ;
  assign n9825 = ~n9821 & ~n9824 ;
  assign n9826 = x3 & ~n9825 ;
  assign n9827 = ~n9819 & ~n9826 ;
  assign n9828 = x1 & ~n9827 ;
  assign n9829 = ~n9816 & ~n9828 ;
  assign n9830 = ~x8 & n1667 ;
  assign n9831 = ~x15 & n3555 ;
  assign n9832 = ~n633 & ~n9831 ;
  assign n9833 = n9830 & ~n9832 ;
  assign n9834 = x9 & n3960 ;
  assign n9835 = n2358 & n9834 ;
  assign n9836 = ~n2508 & ~n6020 ;
  assign n9837 = ~n9835 & ~n9836 ;
  assign n9838 = n464 & ~n9837 ;
  assign n9839 = ~n9833 & ~n9838 ;
  assign n9840 = n462 & ~n9839 ;
  assign n9841 = n1202 & n4196 ;
  assign n9842 = n7854 & n9841 ;
  assign n9843 = n3228 & n7926 ;
  assign n9844 = ~n870 & n900 ;
  assign n9845 = n9843 & n9844 ;
  assign n9846 = ~n9842 & ~n9845 ;
  assign n9847 = n1563 & ~n9846 ;
  assign n9848 = ~x9 & n76 ;
  assign n9849 = ~n1263 & ~n9848 ;
  assign n9850 = n405 & ~n9849 ;
  assign n9851 = n1272 & n9850 ;
  assign n9852 = n557 & n1742 ;
  assign n9853 = n162 & n9852 ;
  assign n9854 = n633 & n9853 ;
  assign n9855 = ~n9851 & ~n9854 ;
  assign n9856 = ~n9847 & n9855 ;
  assign n9857 = n18 & n76 ;
  assign n9858 = n2358 & n9857 ;
  assign n9859 = n2023 & n2083 ;
  assign n9860 = n328 & n530 ;
  assign n9861 = n453 & n9860 ;
  assign n9862 = ~n9859 & ~n9861 ;
  assign n9863 = ~n9858 & n9862 ;
  assign n9864 = n230 & ~n9863 ;
  assign n9865 = n265 & n986 ;
  assign n9866 = n863 & n1364 ;
  assign n9867 = ~n4794 & ~n9866 ;
  assign n9868 = ~n9865 & n9867 ;
  assign n9869 = n690 & n4851 ;
  assign n9870 = ~n9868 & n9869 ;
  assign n9871 = ~n9864 & ~n9870 ;
  assign n9872 = n9856 & n9871 ;
  assign n9873 = ~n9840 & n9872 ;
  assign n9874 = n9829 & n9873 ;
  assign n9875 = n929 & ~n9874 ;
  assign n9876 = ~n9808 & ~n9875 ;
  assign n9877 = n438 & ~n1658 ;
  assign n9878 = n4954 & n7692 ;
  assign n9879 = n9877 & n9878 ;
  assign n9880 = n414 & n1869 ;
  assign n9881 = n5193 & n6936 ;
  assign n9882 = ~n9880 & ~n9881 ;
  assign n9883 = n1664 & ~n9882 ;
  assign n9884 = n151 & n9883 ;
  assign n9885 = n333 & n986 ;
  assign n9886 = n1980 & n9885 ;
  assign n9887 = n9886 ^ x8 ;
  assign n9888 = n9887 ^ n9886 ;
  assign n9889 = n9888 ^ n9884 ;
  assign n9890 = n5327 & n5698 ;
  assign n9891 = n442 & n986 ;
  assign n9892 = n9891 ^ n104 ;
  assign n9893 = n2477 ^ x11 ;
  assign n9894 = n2477 ^ x9 ;
  assign n9895 = n9894 ^ n2477 ;
  assign n9896 = ~n9893 & ~n9895 ;
  assign n9897 = n9896 ^ n2477 ;
  assign n9898 = n9897 ^ n9891 ;
  assign n9899 = ~n9892 & ~n9898 ;
  assign n9900 = n9899 ^ n9896 ;
  assign n9901 = n9900 ^ n2477 ;
  assign n9902 = n9901 ^ n104 ;
  assign n9903 = n9891 & n9902 ;
  assign n9904 = n9903 ^ n9891 ;
  assign n9905 = ~n9890 & ~n9904 ;
  assign n9906 = n9905 ^ n58 ;
  assign n9907 = ~n9905 & ~n9906 ;
  assign n9908 = n9907 ^ n9886 ;
  assign n9909 = n9908 ^ n9905 ;
  assign n9910 = n9889 & ~n9909 ;
  assign n9911 = n9910 ^ n9907 ;
  assign n9912 = n9911 ^ n9905 ;
  assign n9913 = ~n9884 & ~n9912 ;
  assign n9914 = n9913 ^ n9884 ;
  assign n9915 = ~n3229 & n9914 ;
  assign n9916 = ~n9879 & ~n9915 ;
  assign n9917 = n9916 ^ n9876 ;
  assign n9918 = n66 & n5888 ;
  assign n9919 = ~n24 & ~n1092 ;
  assign n9920 = ~n9918 & ~n9919 ;
  assign n9921 = ~n333 & n9920 ;
  assign n9922 = x12 & ~n9921 ;
  assign n9923 = n58 & n1665 ;
  assign n9924 = ~n1227 & n9923 ;
  assign n9925 = ~x2 & n38 ;
  assign n9926 = ~n1990 & ~n9925 ;
  assign n9927 = ~n7230 & ~n9926 ;
  assign n9928 = n9683 & ~n9927 ;
  assign n9929 = ~n9924 & n9928 ;
  assign n9930 = ~n9922 & n9929 ;
  assign n9931 = n517 & ~n9930 ;
  assign n9932 = n2738 & ~n4656 ;
  assign n9933 = n3146 & n4098 ;
  assign n9934 = ~n2356 & ~n9933 ;
  assign n9935 = ~n9932 & n9934 ;
  assign n9936 = n928 & ~n9935 ;
  assign n9937 = ~n56 & n9936 ;
  assign n9938 = n6436 & ~n9600 ;
  assign n9939 = n1667 ^ x2 ;
  assign n9940 = x12 ^ x0 ;
  assign n9941 = n9940 ^ x12 ;
  assign n9942 = n2326 ^ x12 ;
  assign n9943 = n9941 & n9942 ;
  assign n9944 = n9943 ^ x12 ;
  assign n9945 = n9944 ^ n1667 ;
  assign n9946 = ~n9939 & ~n9945 ;
  assign n9947 = n9946 ^ n9943 ;
  assign n9948 = n9947 ^ x12 ;
  assign n9949 = n9948 ^ x2 ;
  assign n9950 = ~n1667 & n9949 ;
  assign n9951 = n9950 ^ n1667 ;
  assign n9952 = ~n9938 & n9951 ;
  assign n9953 = ~n20 & n462 ;
  assign n9954 = ~n9952 & n9953 ;
  assign n9955 = n301 & n2290 ;
  assign n9956 = n66 & n9955 ;
  assign n9957 = ~n318 & ~n4887 ;
  assign n9958 = n261 & ~n9957 ;
  assign n9959 = ~n9956 & ~n9958 ;
  assign n9960 = n9958 ^ n7539 ;
  assign n9961 = n9959 ^ n70 ;
  assign n9962 = n9960 & n9961 ;
  assign n9963 = n9962 ^ n70 ;
  assign n9964 = n9959 & n9963 ;
  assign n9965 = ~n9954 & n9964 ;
  assign n9966 = ~x9 & ~n9965 ;
  assign n9967 = n439 & n1645 ;
  assign n9968 = n639 & n5163 ;
  assign n9969 = ~n9967 & ~n9968 ;
  assign n9970 = ~n9966 & n9969 ;
  assign n9971 = ~n9937 & n9970 ;
  assign n9972 = n434 & n4098 ;
  assign n9973 = n45 & n3960 ;
  assign n9974 = ~n9972 & ~n9973 ;
  assign n9975 = n1627 & ~n9974 ;
  assign n9976 = n318 & n9975 ;
  assign n9977 = n328 & n9918 ;
  assign n9978 = ~n757 & n3960 ;
  assign n9979 = n3697 & n9978 ;
  assign n9980 = ~n176 & ~n5888 ;
  assign n9981 = n9979 & n9980 ;
  assign n9982 = ~n9977 & ~n9981 ;
  assign n9983 = ~x12 & ~n9982 ;
  assign n9984 = n276 & n2272 ;
  assign n9985 = ~n9983 & ~n9984 ;
  assign n9986 = ~n9976 & n9985 ;
  assign n9987 = x11 & ~n9986 ;
  assign n9988 = n9971 & ~n9987 ;
  assign n9989 = ~n9931 & n9988 ;
  assign n9990 = x10 & ~n9989 ;
  assign n9991 = n276 & n928 ;
  assign n9992 = n863 & n9991 ;
  assign n9993 = ~n1030 & ~n2747 ;
  assign n9994 = n177 & ~n9993 ;
  assign n9995 = n888 & ~n5998 ;
  assign n9996 = n1059 & n9995 ;
  assign n9997 = ~n9994 & ~n9996 ;
  assign n9998 = ~n9992 & n9997 ;
  assign n9999 = n2116 & ~n9998 ;
  assign n10000 = x12 & n9991 ;
  assign n10001 = ~n7716 & n10000 ;
  assign n10002 = ~n277 & n5020 ;
  assign n10003 = n2290 & n10002 ;
  assign n10004 = ~n10001 & ~n10003 ;
  assign n10005 = ~n9999 & n10004 ;
  assign n10006 = n690 & ~n10005 ;
  assign n10007 = n109 & n5372 ;
  assign n10008 = n642 & n4333 ;
  assign n10009 = ~n10007 & ~n10008 ;
  assign n10010 = n6998 & ~n10009 ;
  assign n10011 = n659 & n2154 ;
  assign n10012 = ~n10010 & ~n10011 ;
  assign n10013 = n3330 & ~n10012 ;
  assign n10014 = ~x10 & ~n1642 ;
  assign n10015 = x2 & ~n10014 ;
  assign n10016 = ~n55 & ~n176 ;
  assign n10017 = ~n18 & ~n375 ;
  assign n10018 = ~n10016 & n10017 ;
  assign n10019 = ~n530 & n762 ;
  assign n10020 = x13 & ~n8808 ;
  assign n10021 = n10019 & ~n10020 ;
  assign n10022 = n10018 & n10021 ;
  assign n10023 = ~n10015 & n10022 ;
  assign n10024 = n845 & n1377 ;
  assign n10025 = n163 & n10024 ;
  assign n10026 = ~n10023 & ~n10025 ;
  assign n10027 = n1282 & ~n10026 ;
  assign n10028 = ~n10013 & ~n10027 ;
  assign n10029 = ~n10006 & n10028 ;
  assign n10030 = ~n9990 & n10029 ;
  assign n10031 = n10030 ^ x8 ;
  assign n10032 = n10031 ^ n10030 ;
  assign n10033 = ~n70 & ~n7926 ;
  assign n10034 = ~n142 & ~n1478 ;
  assign n10035 = n224 & n10034 ;
  assign n10036 = ~n10033 & ~n10035 ;
  assign n10037 = ~n1090 & n10036 ;
  assign n10038 = n346 & ~n10037 ;
  assign n10039 = ~x15 & ~n332 ;
  assign n10040 = n68 ^ n65 ;
  assign n10041 = ~n4339 & n10040 ;
  assign n10042 = n10041 ^ n65 ;
  assign n10043 = n698 & n10042 ;
  assign n10044 = ~n10039 & n10043 ;
  assign n10045 = ~n10038 & ~n10044 ;
  assign n10046 = n1905 & ~n10045 ;
  assign n10047 = n4954 & n6597 ;
  assign n10048 = n870 & n10047 ;
  assign n10049 = x14 & n10048 ;
  assign n10050 = ~n10046 & ~n10049 ;
  assign n10051 = ~n679 & n1990 ;
  assign n10052 = x3 & ~n142 ;
  assign n10053 = ~n274 & ~n740 ;
  assign n10054 = n10052 & n10053 ;
  assign n10055 = ~n10051 & ~n10054 ;
  assign n10056 = x9 & ~n10055 ;
  assign n10057 = ~n4954 & ~n10056 ;
  assign n10058 = n240 & ~n10057 ;
  assign n10059 = n32 & n284 ;
  assign n10060 = n274 & n10059 ;
  assign n10061 = n105 & n10060 ;
  assign n10062 = ~n10058 & ~n10061 ;
  assign n10063 = n779 & ~n10062 ;
  assign n10064 = n6492 & n7329 ;
  assign n10065 = ~n348 & ~n1270 ;
  assign n10066 = ~n442 & ~n10065 ;
  assign n10067 = n2118 & n10066 ;
  assign n10068 = ~n4735 & ~n10067 ;
  assign n10069 = n1059 & ~n10068 ;
  assign n10070 = ~n10064 & ~n10069 ;
  assign n10071 = n1031 & ~n1092 ;
  assign n10072 = n25 & n1648 ;
  assign n10073 = ~n10071 & ~n10072 ;
  assign n10074 = n10073 ^ n18 ;
  assign n10075 = n10074 ^ n10073 ;
  assign n10076 = n10073 ^ n9683 ;
  assign n10077 = n10076 ^ n10073 ;
  assign n10078 = n10075 & ~n10077 ;
  assign n10079 = n10078 ^ n10073 ;
  assign n10080 = x11 & ~n10079 ;
  assign n10081 = n10080 ^ n10073 ;
  assign n10082 = n7180 & ~n10081 ;
  assign n10083 = n10070 & ~n10082 ;
  assign n10084 = ~n10063 & n10083 ;
  assign n10085 = n10050 & n10084 ;
  assign n10086 = x12 & ~n10085 ;
  assign n10087 = n700 & n1328 ;
  assign n10088 = ~x11 & n9604 ;
  assign n10089 = ~n10087 & ~n10088 ;
  assign n10090 = n354 & ~n10089 ;
  assign n10091 = n3040 ^ x9 ;
  assign n10092 = n10091 ^ n3040 ;
  assign n10093 = n10092 ^ n1283 ;
  assign n10094 = n1283 ^ n24 ;
  assign n10095 = x10 & ~n10094 ;
  assign n10096 = n10095 ^ n3040 ;
  assign n10097 = n10093 & ~n10096 ;
  assign n10098 = n10097 ^ n10095 ;
  assign n10099 = ~n1283 & n10098 ;
  assign n10100 = n10099 ^ n10095 ;
  assign n10101 = n10100 ^ n10097 ;
  assign n10102 = ~x1 & n10101 ;
  assign n10103 = ~n10090 & ~n10102 ;
  assign n10104 = n6490 & ~n10103 ;
  assign n10105 = n4179 & n6075 ;
  assign n10106 = n393 & n453 ;
  assign n10107 = n568 & ~n1038 ;
  assign n10108 = ~n10106 & ~n10107 ;
  assign n10109 = n6998 & ~n10108 ;
  assign n10110 = n197 & n9857 ;
  assign n10111 = ~n1283 & n1967 ;
  assign n10112 = n346 & ~n10111 ;
  assign n10113 = ~x15 & n828 ;
  assign n10114 = n2389 & n10113 ;
  assign n10115 = ~n10112 & ~n10114 ;
  assign n10116 = n1905 & ~n10115 ;
  assign n10117 = ~n10110 & ~n10116 ;
  assign n10118 = ~n10109 & n10117 ;
  assign n10119 = n318 & ~n10118 ;
  assign n10120 = ~n10105 & ~n10119 ;
  assign n10121 = x0 & ~n10120 ;
  assign n10122 = n67 & n779 ;
  assign n10123 = n5615 & n10122 ;
  assign n10124 = ~n10121 & ~n10123 ;
  assign n10125 = ~n10104 & n10124 ;
  assign n10126 = ~n10086 & n10125 ;
  assign n10127 = n10126 ^ n10030 ;
  assign n10128 = ~n10032 & n10127 ;
  assign n10129 = n10128 ^ n10030 ;
  assign n10130 = n10129 ^ n9876 ;
  assign n10131 = n9917 & n10130 ;
  assign n10132 = n10131 ^ n10128 ;
  assign n10133 = n10132 ^ n10030 ;
  assign n10134 = n10133 ^ n9916 ;
  assign n10135 = n9876 & n10134 ;
  assign n10136 = n10135 ^ n9876 ;
  assign n10137 = n9724 & n10136 ;
  assign n10138 = ~n9598 & ~n10137 ;
  assign n10139 = ~n260 & ~n3307 ;
  assign n10140 = n65 & ~n10139 ;
  assign n10141 = n7585 & n10140 ;
  assign n10142 = ~x2 & n366 ;
  assign n10143 = n3106 & n10142 ;
  assign n10144 = n1555 & n10143 ;
  assign n10145 = ~n10141 & ~n10144 ;
  assign n10146 = n489 & ~n10145 ;
  assign n10147 = n2568 & n10142 ;
  assign n10148 = n2861 & n10147 ;
  assign n10149 = ~n10146 & ~n10148 ;
  assign n10150 = x15 & ~n10149 ;
  assign n10151 = n65 & n8854 ;
  assign n10152 = n3894 & n10151 ;
  assign n10153 = ~n10150 & ~n10152 ;
  assign n10154 = ~n8686 & ~n10153 ;
  assign n10155 = n65 & n1124 ;
  assign n10156 = ~n8311 & ~n10155 ;
  assign n10157 = n60 & ~n10156 ;
  assign n10158 = ~n9015 & ~n10157 ;
  assign n10159 = ~n8019 & ~n10158 ;
  assign n10160 = n301 & n427 ;
  assign n10161 = n10160 ^ n2973 ;
  assign n10162 = n10161 ^ n7103 ;
  assign n10163 = n10162 ^ n10160 ;
  assign n10164 = n10163 ^ n10162 ;
  assign n10165 = ~n3960 & ~n8310 ;
  assign n10166 = n10165 ^ n10162 ;
  assign n10167 = n10166 ^ n10161 ;
  assign n10168 = n10164 & ~n10167 ;
  assign n10169 = n10168 ^ n10165 ;
  assign n10170 = ~x10 & ~n10165 ;
  assign n10171 = n10170 ^ n10161 ;
  assign n10172 = ~n10169 & ~n10171 ;
  assign n10173 = n10172 ^ n10170 ;
  assign n10174 = ~n10161 & n10173 ;
  assign n10175 = n10174 ^ n10168 ;
  assign n10176 = n10175 ^ n2973 ;
  assign n10177 = n10176 ^ n10165 ;
  assign n10178 = n164 & ~n10177 ;
  assign n10179 = n2280 & ~n3012 ;
  assign n10180 = ~x10 & n1912 ;
  assign n10181 = ~n10179 & ~n10180 ;
  assign n10182 = x3 & n2995 ;
  assign n10183 = ~n10181 & n10182 ;
  assign n10184 = x10 ^ x0 ;
  assign n10185 = n10184 ^ x14 ;
  assign n10186 = n2608 ^ x10 ;
  assign n10187 = n10186 ^ n2608 ;
  assign n10188 = n10187 ^ n10185 ;
  assign n10189 = n2535 ^ x14 ;
  assign n10190 = n2535 & n10189 ;
  assign n10191 = n10190 ^ n2608 ;
  assign n10192 = n10191 ^ n2535 ;
  assign n10193 = n10188 & n10192 ;
  assign n10194 = n10193 ^ n10190 ;
  assign n10195 = n10194 ^ n2535 ;
  assign n10196 = n10185 & n10195 ;
  assign n10197 = n217 & n10196 ;
  assign n10198 = n1164 & n3072 ;
  assign n10199 = ~n10197 & ~n10198 ;
  assign n10200 = n232 & ~n10199 ;
  assign n10201 = n26 & n2612 ;
  assign n10202 = n260 & n10201 ;
  assign n10203 = n6484 & n10202 ;
  assign n10204 = ~n3207 & ~n10201 ;
  assign n10205 = n10204 ^ x10 ;
  assign n10206 = n10205 ^ n10204 ;
  assign n10207 = n10204 ^ n3425 ;
  assign n10208 = n10207 ^ n10204 ;
  assign n10209 = ~n10206 & n10208 ;
  assign n10210 = n10209 ^ n10204 ;
  assign n10211 = ~x3 & ~n10210 ;
  assign n10212 = n10211 ^ n10204 ;
  assign n10213 = n3307 & ~n10212 ;
  assign n10214 = n740 & n10213 ;
  assign n10215 = ~n10203 & ~n10214 ;
  assign n10216 = ~n10200 & n10215 ;
  assign n10217 = ~n10183 & n10216 ;
  assign n10218 = n4339 & ~n10217 ;
  assign n10219 = ~n260 & ~n6097 ;
  assign n10220 = n784 & ~n10219 ;
  assign n10221 = ~n328 & ~n1555 ;
  assign n10222 = n946 & ~n3960 ;
  assign n10223 = ~n10221 & n10222 ;
  assign n10224 = ~n10220 & ~n10223 ;
  assign n10225 = ~n2803 & n3530 ;
  assign n10226 = ~n10224 & n10225 ;
  assign n10227 = n311 & n2904 ;
  assign n10228 = n2973 & n10227 ;
  assign n10229 = n383 & ~n3960 ;
  assign n10230 = x14 & n414 ;
  assign n10231 = ~n10229 & ~n10230 ;
  assign n10232 = n2974 & ~n10231 ;
  assign n10233 = ~n10228 & ~n10232 ;
  assign n10234 = ~n10226 & n10233 ;
  assign n10235 = n79 & ~n10234 ;
  assign n10236 = n8732 & n10151 ;
  assign n10237 = ~n10235 & ~n10236 ;
  assign n10238 = ~n10218 & n10237 ;
  assign n10239 = ~n10178 & n10238 ;
  assign n10240 = n10239 ^ x7 ;
  assign n10241 = n10240 ^ n10239 ;
  assign n10242 = n10241 ^ n10159 ;
  assign n10243 = n5214 & n8147 ;
  assign n10244 = n524 & n2973 ;
  assign n10245 = ~n10243 & ~n10244 ;
  assign n10246 = n164 & ~n10245 ;
  assign n10247 = n762 & n2535 ;
  assign n10248 = n779 & n10247 ;
  assign n10249 = n427 & ~n3012 ;
  assign n10250 = n3530 & n10249 ;
  assign n10251 = n7611 & ~n10139 ;
  assign n10252 = n2973 & n10251 ;
  assign n10253 = ~n10250 & ~n10252 ;
  assign n10254 = ~n10248 & n10253 ;
  assign n10255 = n5851 & ~n10254 ;
  assign n10256 = n232 & ~n3960 ;
  assign n10257 = n3010 & n4015 ;
  assign n10258 = ~n10256 & ~n10257 ;
  assign n10259 = ~n8705 & n10258 ;
  assign n10260 = n7103 & ~n10259 ;
  assign n10261 = n40 & n3894 ;
  assign n10262 = n2282 & n10261 ;
  assign n10263 = n7611 & n10262 ;
  assign n10264 = ~n10260 & ~n10263 ;
  assign n10265 = n109 & ~n10264 ;
  assign n10266 = ~x3 & ~n10265 ;
  assign n10267 = ~n10255 & n10266 ;
  assign n10268 = ~n10246 & n10267 ;
  assign n10269 = ~x10 & n403 ;
  assign n10270 = ~n516 & ~n10269 ;
  assign n10271 = x11 & ~n10270 ;
  assign n10272 = n739 & n978 ;
  assign n10273 = n8093 ^ n5976 ;
  assign n10274 = n8093 ^ x10 ;
  assign n10275 = n10274 ^ n8093 ;
  assign n10276 = n10275 ^ n10272 ;
  assign n10277 = n10273 & n10276 ;
  assign n10278 = n10277 ^ n5976 ;
  assign n10279 = n10272 & n10278 ;
  assign n10280 = ~n10271 & ~n10279 ;
  assign n10281 = n3427 & ~n10280 ;
  assign n10282 = n3564 & n3867 ;
  assign n10283 = n5976 & n10282 ;
  assign n10284 = x3 & ~n10283 ;
  assign n10285 = ~n10281 & n10284 ;
  assign n10286 = n10285 ^ n10268 ;
  assign n10287 = ~n10268 & n10286 ;
  assign n10288 = n10287 ^ n10239 ;
  assign n10289 = n10288 ^ n10268 ;
  assign n10290 = ~n10242 & n10289 ;
  assign n10291 = n10290 ^ n10287 ;
  assign n10292 = n10291 ^ n10268 ;
  assign n10293 = ~n10159 & ~n10292 ;
  assign n10294 = n10293 ^ n10159 ;
  assign n10295 = ~n10154 & ~n10294 ;
  assign n10296 = ~n828 & ~n1275 ;
  assign n10297 = ~n10295 & ~n10296 ;
  assign n10298 = ~n1276 & n10297 ;
  assign n10299 = n58 & n363 ;
  assign n10300 = n2213 & n10299 ;
  assign n10301 = n2877 & n10300 ;
  assign n10302 = n4019 & n10301 ;
  assign n10303 = n739 & n8703 ;
  assign n10304 = n3403 & n4471 ;
  assign n10305 = ~n10303 & ~n10304 ;
  assign n10306 = n849 & ~n10305 ;
  assign n10307 = n311 & n10306 ;
  assign n10308 = n2394 & n2807 ;
  assign n10309 = n928 & n1010 ;
  assign n10310 = n10308 & n10309 ;
  assign n10311 = ~n6276 & ~n9033 ;
  assign n10312 = ~x9 & ~n8464 ;
  assign n10313 = n2599 & n10312 ;
  assign n10314 = ~n10311 & n10313 ;
  assign n10315 = n290 & n2995 ;
  assign n10316 = n4471 & n10315 ;
  assign n10317 = ~n10314 & ~n10316 ;
  assign n10318 = n365 & ~n10317 ;
  assign n10319 = ~n10310 & ~n10318 ;
  assign n10320 = n700 & ~n10319 ;
  assign n10334 = n1422 & ~n3960 ;
  assign n10335 = n4769 & n10334 ;
  assign n10336 = n44 & n9146 ;
  assign n10337 = ~n10335 & ~n10336 ;
  assign n10338 = n795 & ~n10337 ;
  assign n10339 = ~n1031 & n10338 ;
  assign n10340 = n739 & n1030 ;
  assign n10341 = n5996 & n10340 ;
  assign n10342 = n9114 & n10341 ;
  assign n10343 = ~n10339 & ~n10342 ;
  assign n10321 = n1422 & n5256 ;
  assign n10322 = n10321 ^ n633 ;
  assign n10323 = n10322 ^ n10321 ;
  assign n10324 = n10321 ^ n2806 ;
  assign n10325 = n10324 ^ n10321 ;
  assign n10326 = n10323 & n10325 ;
  assign n10327 = n10326 ^ n10321 ;
  assign n10328 = ~x8 & n10327 ;
  assign n10329 = n10328 ^ n10321 ;
  assign n10330 = n739 & n10329 ;
  assign n10331 = x2 & n10330 ;
  assign n10332 = n3019 & n9436 ;
  assign n10333 = ~n10331 & ~n10332 ;
  assign n10344 = n10343 ^ n10333 ;
  assign n10345 = n10344 ^ n10343 ;
  assign n10346 = n10343 ^ x10 ;
  assign n10347 = n10346 ^ n10343 ;
  assign n10348 = ~n10345 & n10347 ;
  assign n10349 = n10348 ^ n10343 ;
  assign n10350 = x11 & ~n10349 ;
  assign n10351 = n10350 ^ n10343 ;
  assign n10352 = n261 & ~n10351 ;
  assign n10353 = ~n10320 & ~n10352 ;
  assign n10354 = ~n10307 & n10353 ;
  assign n10355 = n10354 ^ x12 ;
  assign n10356 = n10355 ^ n10354 ;
  assign n10357 = n10356 ^ n10302 ;
  assign n10358 = n2634 & n3361 ;
  assign n10359 = n7337 & n10358 ;
  assign n10360 = n6924 & n10359 ;
  assign n10361 = n7044 & n8703 ;
  assign n10362 = n2806 & n5526 ;
  assign n10363 = n60 & n10362 ;
  assign n10364 = ~n10361 & ~n10363 ;
  assign n10365 = n2033 & ~n10364 ;
  assign n10366 = n4222 & n8963 ;
  assign n10367 = n2075 & n10366 ;
  assign n10368 = ~n10365 & ~n10367 ;
  assign n10369 = ~n10360 & n10368 ;
  assign n10370 = n10369 ^ x2 ;
  assign n10371 = ~n10369 & n10370 ;
  assign n10372 = n10371 ^ n10354 ;
  assign n10373 = n10372 ^ n10369 ;
  assign n10374 = ~n10357 & n10373 ;
  assign n10375 = n10374 ^ n10371 ;
  assign n10376 = n10375 ^ n10369 ;
  assign n10377 = ~n10302 & ~n10376 ;
  assign n10378 = n10377 ^ n10302 ;
  assign n10379 = ~n4881 & n10378 ;
  assign n10380 = ~n10298 & ~n10379 ;
  assign n10381 = ~n10138 & n10380 ;
  assign n10382 = ~n2461 & ~n2471 ;
  assign n10383 = n1464 & n7631 ;
  assign n10384 = ~x15 & n10383 ;
  assign n10385 = ~n6373 & ~n10384 ;
  assign n10386 = n66 & ~n10385 ;
  assign n10387 = n344 & n2562 ;
  assign n10388 = n1665 & n10387 ;
  assign n10389 = n163 & n7899 ;
  assign n10390 = n168 & ~n986 ;
  assign n10391 = ~n3761 & n10390 ;
  assign n10392 = ~n10389 & ~n10391 ;
  assign n10393 = ~x12 & ~n10392 ;
  assign n10394 = ~n10383 & ~n10393 ;
  assign n10395 = n306 & ~n10394 ;
  assign n10396 = ~n10388 & ~n10395 ;
  assign n10397 = ~n10386 & n10396 ;
  assign n10398 = n3091 & ~n10397 ;
  assign n10399 = ~n1227 & ~n7181 ;
  assign n10400 = ~x1 & n10399 ;
  assign n10401 = ~n7808 & ~n10400 ;
  assign n10402 = n4338 & ~n10401 ;
  assign n10403 = n2778 & n10402 ;
  assign n10404 = n145 & n1782 ;
  assign n10405 = n38 & n7718 ;
  assign n10406 = ~n10404 & ~n10405 ;
  assign n10407 = n3021 & n9420 ;
  assign n10408 = ~n10406 & n10407 ;
  assign n10409 = ~n10403 & ~n10408 ;
  assign n10410 = ~n10398 & n10409 ;
  assign n10411 = ~x7 & n10399 ;
  assign n10412 = ~x14 & n9274 ;
  assign n10413 = x12 & n10412 ;
  assign n10414 = ~n10411 & ~n10413 ;
  assign n10415 = n34 & ~n10414 ;
  assign n10416 = n2873 & ~n10412 ;
  assign n10417 = n1113 & n10416 ;
  assign n10418 = ~n10415 & ~n10417 ;
  assign n10419 = n10418 ^ x3 ;
  assign n10420 = n10419 ^ n10418 ;
  assign n10421 = n828 & n3960 ;
  assign n10422 = ~n1214 & ~n10421 ;
  assign n10423 = n10422 ^ x12 ;
  assign n10424 = ~x7 & ~n10423 ;
  assign n10425 = n10424 ^ x12 ;
  assign n10426 = n89 & n10425 ;
  assign n10427 = n10426 ^ n10418 ;
  assign n10428 = n10420 & ~n10427 ;
  assign n10429 = n10428 ^ n10418 ;
  assign n10430 = n7041 & ~n10429 ;
  assign n10431 = n10410 & ~n10430 ;
  assign n10432 = n25 & n85 ;
  assign n10433 = n1113 & ~n2370 ;
  assign n10434 = ~n10432 & ~n10433 ;
  assign n10435 = n10434 ^ n168 ;
  assign n10436 = n10435 ^ n10434 ;
  assign n10437 = x0 & ~n673 ;
  assign n10438 = ~n3960 & ~n10437 ;
  assign n10439 = n10438 ^ n10434 ;
  assign n10440 = n10439 ^ n10434 ;
  assign n10441 = n10436 & ~n10440 ;
  assign n10442 = n10441 ^ n10434 ;
  assign n10443 = x12 & ~n10442 ;
  assign n10444 = n10443 ^ n10434 ;
  assign n10445 = n10444 ^ x7 ;
  assign n10446 = n10445 ^ n10444 ;
  assign n10447 = n10446 ^ n6905 ;
  assign n10448 = n1282 & n10390 ;
  assign n10449 = ~n163 & ~n6037 ;
  assign n10450 = ~n196 & ~n2036 ;
  assign n10451 = x0 & n10450 ;
  assign n10452 = ~n10449 & n10451 ;
  assign n10453 = ~n10448 & ~n10452 ;
  assign n10454 = ~n4026 & ~n7692 ;
  assign n10455 = ~n2036 & n2679 ;
  assign n10456 = ~n10454 & n10455 ;
  assign n10457 = n10456 ^ n10453 ;
  assign n10458 = n10453 & ~n10457 ;
  assign n10459 = n10458 ^ n10444 ;
  assign n10460 = n10459 ^ n10453 ;
  assign n10461 = n10447 & n10460 ;
  assign n10462 = n10461 ^ n10458 ;
  assign n10463 = n10462 ^ n10453 ;
  assign n10464 = n6905 & n10463 ;
  assign n10465 = n10464 ^ n6905 ;
  assign n10466 = n10431 & ~n10465 ;
  assign n10467 = ~n8645 & ~n10466 ;
  assign n10468 = ~n7539 & n8017 ;
  assign n10469 = n8684 & n10113 ;
  assign n10470 = n2653 & n10469 ;
  assign n10471 = ~n10468 & ~n10470 ;
  assign n10472 = n1645 & ~n10471 ;
  assign n10473 = ~n10467 & ~n10472 ;
  assign n10474 = n690 & n3408 ;
  assign n10475 = x5 ^ x1 ;
  assign n10476 = n17 & ~n1227 ;
  assign n10477 = n344 & n10476 ;
  assign n10478 = n828 & n10412 ;
  assign n10479 = ~n6150 & ~n10478 ;
  assign n10480 = n344 & ~n10479 ;
  assign n10481 = ~n10477 & ~n10480 ;
  assign n10482 = n10481 ^ n10475 ;
  assign n10483 = ~x7 & n3960 ;
  assign n10484 = n1282 & n9274 ;
  assign n10485 = ~n10483 & ~n10484 ;
  assign n10486 = ~x13 & ~n10485 ;
  assign n10487 = ~n2512 & ~n10486 ;
  assign n10488 = ~n1227 & ~n10487 ;
  assign n10489 = n10488 ^ x1 ;
  assign n10490 = n10489 ^ n10488 ;
  assign n10491 = n3021 & ~n5698 ;
  assign n10492 = ~n9275 & n10491 ;
  assign n10493 = ~n2036 & ~n5698 ;
  assign n10494 = x14 & n10493 ;
  assign n10495 = ~x7 & n10494 ;
  assign n10496 = ~n10492 & ~n10495 ;
  assign n10497 = n10496 ^ n10488 ;
  assign n10498 = ~n10490 & ~n10497 ;
  assign n10499 = n10498 ^ n10488 ;
  assign n10500 = n10499 ^ n10475 ;
  assign n10501 = n10482 & n10500 ;
  assign n10502 = n10501 ^ n10498 ;
  assign n10503 = n10502 ^ n10488 ;
  assign n10504 = n10503 ^ n10481 ;
  assign n10505 = n10475 & n10504 ;
  assign n10506 = n10505 ^ n10475 ;
  assign n10507 = n10506 ^ n10481 ;
  assign n10508 = x2 & ~n10507 ;
  assign n10509 = ~n10474 & ~n10508 ;
  assign n10510 = n2815 & ~n10509 ;
  assign n10511 = ~n679 & ~n3960 ;
  assign n10512 = ~n332 & ~n10511 ;
  assign n10513 = ~n32 & n2678 ;
  assign n10514 = ~n10512 & n10513 ;
  assign n10515 = n718 & ~n9274 ;
  assign n10516 = ~n1042 & n10515 ;
  assign n10517 = n2558 & ~n4829 ;
  assign n10518 = ~n9656 & n10517 ;
  assign n10519 = ~n10516 & ~n10518 ;
  assign n10520 = ~n74 & ~n10519 ;
  assign n10521 = ~n10514 & ~n10520 ;
  assign n10522 = n1641 & ~n10521 ;
  assign n10523 = x7 ^ x1 ;
  assign n10524 = n10523 ^ n10476 ;
  assign n10525 = n1327 ^ x1 ;
  assign n10526 = n10525 ^ n1327 ;
  assign n10527 = n6294 ^ n1327 ;
  assign n10528 = n10526 & n10527 ;
  assign n10529 = n10528 ^ n1327 ;
  assign n10530 = n10529 ^ n10523 ;
  assign n10531 = ~n10524 & ~n10530 ;
  assign n10532 = n10531 ^ n10528 ;
  assign n10533 = n10532 ^ n1327 ;
  assign n10534 = n10533 ^ n10476 ;
  assign n10535 = n10523 & n10534 ;
  assign n10536 = n10535 ^ n10523 ;
  assign n10537 = n10536 ^ n10476 ;
  assign n10538 = n213 & n10537 ;
  assign n10539 = ~n176 & ~n3019 ;
  assign n10540 = ~n3960 & n10539 ;
  assign n10541 = n1042 & ~n10540 ;
  assign n10542 = ~n205 & ~n10541 ;
  assign n10543 = n6037 & ~n10542 ;
  assign n10544 = ~x1 & ~n4166 ;
  assign n10545 = x12 & ~n10544 ;
  assign n10546 = ~n3263 & n10545 ;
  assign n10547 = ~n6248 & ~n10546 ;
  assign n10548 = n497 & ~n10547 ;
  assign n10549 = ~n10543 & ~n10548 ;
  assign n10550 = ~n10538 & n10549 ;
  assign n10551 = ~n10522 & n10550 ;
  assign n10552 = n2562 & ~n10551 ;
  assign n10553 = n233 & n10494 ;
  assign n10554 = x2 & ~n160 ;
  assign n10555 = n8527 & n10554 ;
  assign n10556 = ~n10553 & ~n10555 ;
  assign n10557 = n2712 & ~n10556 ;
  assign n10558 = n6628 & n7041 ;
  assign n10559 = n1683 & n10558 ;
  assign n10560 = ~n10557 & ~n10559 ;
  assign n10561 = n1678 & n7180 ;
  assign n10562 = ~n76 & n8944 ;
  assign n10563 = ~x0 & n10562 ;
  assign n10564 = ~x5 & ~n2796 ;
  assign n10565 = ~n10563 & n10564 ;
  assign n10566 = ~n10561 & ~n10565 ;
  assign n10567 = n141 & ~n10566 ;
  assign n10568 = ~n58 & ~n2282 ;
  assign n10569 = n8707 & n10568 ;
  assign n10570 = n1349 & n1991 ;
  assign n10571 = ~n10569 & n10570 ;
  assign n10572 = ~n89 & ~n929 ;
  assign n10573 = ~x0 & n176 ;
  assign n10574 = ~x5 & n10573 ;
  assign n10575 = n7539 & ~n10574 ;
  assign n10576 = ~n10572 & ~n10575 ;
  assign n10577 = ~x1 & n10576 ;
  assign n10578 = ~n10571 & ~n10577 ;
  assign n10579 = ~n10567 & n10578 ;
  assign n10580 = n2806 & ~n10579 ;
  assign n10581 = n10560 & ~n10580 ;
  assign n10582 = ~n10552 & n10581 ;
  assign n10583 = ~n10510 & n10582 ;
  assign n10584 = n366 & ~n10583 ;
  assign n10585 = n7041 & n7163 ;
  assign n10586 = n4344 & n10585 ;
  assign n10587 = n33 & n3091 ;
  assign n10588 = n6037 & n10587 ;
  assign n10589 = n2583 & n4656 ;
  assign n10590 = n10589 ^ n10496 ;
  assign n10591 = n10590 ^ n10496 ;
  assign n10592 = n10496 ^ x13 ;
  assign n10593 = n10592 ^ n10496 ;
  assign n10594 = n10591 & ~n10593 ;
  assign n10595 = n10594 ^ n10496 ;
  assign n10596 = x6 & ~n10595 ;
  assign n10597 = n10596 ^ n10496 ;
  assign n10598 = n2343 & ~n10597 ;
  assign n10599 = ~n1227 & n2881 ;
  assign n10600 = n1382 & n10599 ;
  assign n10601 = n1422 & n7808 ;
  assign n10602 = ~n2356 & ~n7277 ;
  assign n10603 = n2806 & ~n10602 ;
  assign n10604 = ~n10601 & ~n10603 ;
  assign n10605 = ~n10600 & n10604 ;
  assign n10606 = n196 & ~n10605 ;
  assign n10607 = ~n10598 & ~n10606 ;
  assign n10608 = n10607 ^ x2 ;
  assign n10609 = n10608 ^ n10607 ;
  assign n10610 = n10609 ^ n10588 ;
  assign n10611 = x12 & n10483 ;
  assign n10612 = ~n3199 & ~n10611 ;
  assign n10613 = n1660 & ~n10612 ;
  assign n10614 = n2343 & ~n10414 ;
  assign n10615 = ~n10613 & ~n10614 ;
  assign n10616 = n10615 ^ x6 ;
  assign n10617 = x6 & ~n10616 ;
  assign n10618 = n10617 ^ n10607 ;
  assign n10619 = n10618 ^ x6 ;
  assign n10620 = n10610 & ~n10619 ;
  assign n10621 = n10620 ^ n10617 ;
  assign n10622 = n10621 ^ x6 ;
  assign n10623 = ~n10588 & n10622 ;
  assign n10624 = n10623 ^ n10588 ;
  assign n10625 = ~n10586 & ~n10624 ;
  assign n10626 = ~n3803 & ~n10625 ;
  assign n10627 = x15 ^ x7 ;
  assign n10628 = n5851 ^ x15 ;
  assign n10629 = n10628 ^ n5851 ;
  assign n10630 = n8304 ^ n5851 ;
  assign n10631 = ~n10629 & n10630 ;
  assign n10632 = n10631 ^ n5851 ;
  assign n10633 = n10627 & n10632 ;
  assign n10634 = n195 & n10633 ;
  assign n10635 = n233 & n4166 ;
  assign n10636 = n141 & n9274 ;
  assign n10637 = ~x5 & n10636 ;
  assign n10638 = ~n10635 & ~n10637 ;
  assign n10639 = n1476 & ~n10638 ;
  assign n10640 = ~n10634 & ~n10639 ;
  assign n10641 = ~x3 & ~n10640 ;
  assign n10642 = n302 & n3264 ;
  assign n10643 = n8103 & n9274 ;
  assign n10644 = ~n10642 & ~n10643 ;
  assign n10645 = n2343 & ~n10644 ;
  assign n10646 = ~n10641 & ~n10645 ;
  assign n10647 = n1214 & ~n10646 ;
  assign n10648 = ~x13 & n3286 ;
  assign n10649 = n306 & n1626 ;
  assign n10650 = n712 & n9531 ;
  assign n10651 = ~n10649 & ~n10650 ;
  assign n10652 = n10648 & ~n10651 ;
  assign n10653 = x15 & n10652 ;
  assign n10654 = ~n10647 & ~n10653 ;
  assign n10655 = ~n7473 & ~n10654 ;
  assign n10656 = ~n10626 & ~n10655 ;
  assign n10661 = ~x7 & ~n7539 ;
  assign n10662 = ~n10478 & ~n10661 ;
  assign n10663 = n3427 & ~n10662 ;
  assign n10657 = n919 & ~n7139 ;
  assign n10658 = n3019 & n3175 ;
  assign n10659 = ~n10657 & ~n10658 ;
  assign n10660 = x6 & ~n10659 ;
  assign n10664 = n10663 ^ n10660 ;
  assign n10665 = n10663 ^ x0 ;
  assign n10666 = n10665 ^ n10663 ;
  assign n10667 = n10666 ^ n1996 ;
  assign n10668 = n10664 & ~n10667 ;
  assign n10669 = n10668 ^ n10660 ;
  assign n10670 = n1996 & n10669 ;
  assign n10671 = n10656 & ~n10670 ;
  assign n10672 = ~n10584 & n10671 ;
  assign n10673 = n10473 & n10672 ;
  assign n10772 = n306 & n7631 ;
  assign n10773 = n213 & n10772 ;
  assign n10774 = n2850 & n8685 ;
  assign n10775 = ~n741 & n843 ;
  assign n10776 = x1 & n10483 ;
  assign n10777 = n10775 & n10776 ;
  assign n10778 = ~n10774 & ~n10777 ;
  assign n10779 = ~n10773 & n10778 ;
  assign n10780 = n2182 & ~n10779 ;
  assign n10781 = x1 & ~n10422 ;
  assign n10782 = ~n1382 & ~n10562 ;
  assign n10783 = ~n10781 & ~n10782 ;
  assign n10786 = n10783 ^ n828 ;
  assign n10787 = n10786 ^ n10783 ;
  assign n10784 = n10783 ^ n690 ;
  assign n10785 = n10784 ^ n10783 ;
  assign n10788 = n10787 ^ n10785 ;
  assign n10789 = n10783 ^ x15 ;
  assign n10790 = n10789 ^ n10783 ;
  assign n10791 = n10790 ^ n10787 ;
  assign n10792 = n10787 & ~n10791 ;
  assign n10793 = n10792 ^ n10787 ;
  assign n10794 = n10788 & n10793 ;
  assign n10795 = n10794 ^ n10792 ;
  assign n10796 = n10795 ^ n10783 ;
  assign n10797 = n10796 ^ n10787 ;
  assign n10798 = ~x6 & ~n10797 ;
  assign n10799 = n10798 ^ n10783 ;
  assign n10800 = n884 & ~n10799 ;
  assign n10801 = n673 & ~n6905 ;
  assign n10802 = n2633 & ~n7238 ;
  assign n10803 = x12 & n10802 ;
  assign n10804 = ~n10801 & n10803 ;
  assign n10805 = ~n10800 & ~n10804 ;
  assign n10806 = ~x5 & ~n10805 ;
  assign n10807 = ~n2568 & ~n7041 ;
  assign n10737 = ~x5 & n6824 ;
  assign n10808 = ~n60 & ~n7412 ;
  assign n10809 = n8952 & ~n10808 ;
  assign n10810 = n1382 & n2568 ;
  assign n10811 = ~n3761 & n10810 ;
  assign n10812 = ~n10809 & ~n10811 ;
  assign n10813 = n10737 & ~n10812 ;
  assign n10814 = ~n10807 & n10813 ;
  assign n10815 = n8726 & n10421 ;
  assign n10816 = ~n10814 & ~n10815 ;
  assign n10817 = ~n10806 & n10816 ;
  assign n10818 = n8464 & ~n10817 ;
  assign n10819 = ~n10780 & ~n10818 ;
  assign n10674 = n76 & n884 ;
  assign n10675 = n1382 & n10674 ;
  assign n10676 = n306 & n8204 ;
  assign n10677 = ~n3286 & ~n10113 ;
  assign n10678 = n261 & ~n10677 ;
  assign n10679 = ~n1241 & ~n6824 ;
  assign n10680 = n727 & ~n10679 ;
  assign n10681 = n10544 & n10680 ;
  assign n10682 = n8558 & n10493 ;
  assign n10683 = ~n10681 & ~n10682 ;
  assign n10684 = ~n10678 & n10683 ;
  assign n10685 = n85 & ~n10684 ;
  assign n10686 = ~n10676 & ~n10685 ;
  assign n10687 = ~n10675 & n10686 ;
  assign n10688 = ~x2 & ~n10687 ;
  assign n10689 = ~n1227 & n1742 ;
  assign n10690 = ~n7334 & ~n10689 ;
  assign n10691 = n8331 & ~n10690 ;
  assign n10692 = n2458 & n8283 ;
  assign n10693 = n884 & n3225 ;
  assign n10694 = ~n10692 & ~n10693 ;
  assign n10695 = x1 & ~n10694 ;
  assign n10696 = ~n17 & ~n10648 ;
  assign n10697 = n4829 & ~n10696 ;
  assign n10698 = ~x0 & n10697 ;
  assign n10699 = ~n10695 & ~n10698 ;
  assign n10700 = n8808 & ~n10699 ;
  assign n10701 = n363 & n1743 ;
  assign n10702 = n673 & ~n2633 ;
  assign n10703 = ~n1002 & n6003 ;
  assign n10704 = ~n10702 & n10703 ;
  assign n10705 = n20 & n10412 ;
  assign n10706 = n1742 & n10705 ;
  assign n10707 = ~n10704 & ~n10706 ;
  assign n10708 = ~n10701 & n10707 ;
  assign n10709 = ~n10700 & n10708 ;
  assign n10710 = ~n10691 & n10709 ;
  assign n10711 = x5 & ~n10710 ;
  assign n10712 = n673 & n1742 ;
  assign n10713 = ~n7307 & ~n10712 ;
  assign n10714 = x5 ^ x2 ;
  assign n10715 = n10627 ^ n6418 ;
  assign n10716 = ~n10714 & ~n10715 ;
  assign n10717 = n10716 ^ n10714 ;
  assign n10718 = x7 ^ x5 ;
  assign n10719 = n10718 ^ n10716 ;
  assign n10720 = ~n10627 & n10719 ;
  assign n10721 = n10720 ^ n10627 ;
  assign n10722 = n10721 ^ n6418 ;
  assign n10723 = ~n10717 & ~n10722 ;
  assign n10724 = ~n10713 & n10723 ;
  assign n10725 = ~n10711 & ~n10724 ;
  assign n10726 = ~n10688 & n10725 ;
  assign n10727 = n2701 & ~n10726 ;
  assign n10728 = n712 & n10488 ;
  assign n10729 = n4987 & n9668 ;
  assign n10730 = ~n10728 & ~n10729 ;
  assign n10731 = n7291 & ~n10730 ;
  assign n10732 = n44 & n1630 ;
  assign n10733 = n1034 & n10732 ;
  assign n10734 = ~n2600 & n10733 ;
  assign n10735 = ~n10731 & ~n10734 ;
  assign n10736 = ~n10727 & n10735 ;
  assign n10820 = n10819 ^ n10736 ;
  assign n10821 = n10820 ^ n10736 ;
  assign n10738 = n6574 & n10737 ;
  assign n10739 = x0 & n142 ;
  assign n10740 = n740 & ~n4340 ;
  assign n10741 = ~n10739 & ~n10740 ;
  assign n10742 = n2901 & ~n10741 ;
  assign n10743 = n261 & n6824 ;
  assign n10744 = n232 & n10743 ;
  assign n10745 = ~n10742 & ~n10744 ;
  assign n10746 = ~n10738 & n10745 ;
  assign n10747 = n828 & ~n10746 ;
  assign n10748 = n1400 & n7718 ;
  assign n10749 = ~n3261 & ~n10748 ;
  assign n10750 = n3963 & ~n10749 ;
  assign n10751 = n2036 & n8685 ;
  assign n10752 = ~n10750 & ~n10751 ;
  assign n10753 = ~n10747 & n10752 ;
  assign n10754 = n2701 & ~n10753 ;
  assign n10755 = n127 & n1683 ;
  assign n10756 = ~n1743 & ~n10755 ;
  assign n10757 = ~n8619 & ~n10756 ;
  assign n10758 = n1377 & n2850 ;
  assign n10759 = n4656 & n10758 ;
  assign n10760 = ~n10757 & ~n10759 ;
  assign n10761 = n2901 & ~n10760 ;
  assign n10762 = n58 & n2811 ;
  assign n10763 = ~x7 & n929 ;
  assign n10764 = ~n10762 & ~n10763 ;
  assign n10765 = n739 & n1382 ;
  assign n10766 = ~n10764 & n10765 ;
  assign n10767 = ~n10761 & ~n10766 ;
  assign n10768 = ~n10754 & n10767 ;
  assign n10769 = x14 & ~n10768 ;
  assign n10770 = n10769 ^ n10736 ;
  assign n10771 = n10770 ^ n10736 ;
  assign n10822 = n10821 ^ n10771 ;
  assign n10823 = n7450 ^ x7 ;
  assign n10824 = n10823 ^ n7450 ;
  assign n10825 = n10824 ^ n1641 ;
  assign n10826 = ~n60 & ~n1954 ;
  assign n10827 = ~n1295 & ~n10826 ;
  assign n10828 = ~n8809 & n10827 ;
  assign n10829 = n10828 ^ n718 ;
  assign n10830 = ~n7412 & n10829 ;
  assign n10831 = n10830 ^ n718 ;
  assign n10832 = n126 & n9563 ;
  assign n10833 = n10832 ^ n10831 ;
  assign n10834 = ~n10831 & n10833 ;
  assign n10835 = n10834 ^ n7450 ;
  assign n10836 = n10835 ^ n10831 ;
  assign n10837 = ~n10825 & n10836 ;
  assign n10838 = n10837 ^ n10834 ;
  assign n10839 = n10838 ^ n10831 ;
  assign n10840 = n1641 & ~n10839 ;
  assign n10841 = n10840 ^ n1641 ;
  assign n10842 = ~n24 & n7412 ;
  assign n10843 = ~n2678 & n7041 ;
  assign n10844 = ~n10842 & ~n10843 ;
  assign n10845 = n1702 & ~n10844 ;
  assign n10846 = ~n3960 & n10648 ;
  assign n10847 = ~n8204 & ~n10846 ;
  assign n10848 = ~n160 & ~n10847 ;
  assign n10849 = n1034 & ~n7181 ;
  assign n10850 = n3105 & n10849 ;
  assign n10851 = n3196 & n6295 ;
  assign n10852 = ~n10477 & ~n10851 ;
  assign n10853 = ~n10850 & n10852 ;
  assign n10854 = ~n10848 & n10853 ;
  assign n10855 = ~x6 & ~n10854 ;
  assign n10856 = ~n2902 & n6905 ;
  assign n10857 = ~n1327 & ~n1641 ;
  assign n10858 = n10856 & n10857 ;
  assign n10859 = ~n160 & n2881 ;
  assign n10860 = n828 & n10859 ;
  assign n10861 = ~n10858 & ~n10860 ;
  assign n10862 = ~n10855 & n10861 ;
  assign n10863 = n10862 ^ x0 ;
  assign n10864 = n10863 ^ n10862 ;
  assign n10865 = n10864 ^ n10845 ;
  assign n10866 = ~n2356 & ~n10781 ;
  assign n10867 = n2806 & ~n10866 ;
  assign n10868 = ~n673 & ~n9794 ;
  assign n10869 = ~n7278 & ~n10868 ;
  assign n10870 = n2881 & ~n10869 ;
  assign n10871 = ~n10601 & ~n10870 ;
  assign n10872 = ~n10867 & n10871 ;
  assign n10873 = n10872 ^ x5 ;
  assign n10874 = ~n10872 & n10873 ;
  assign n10875 = n10874 ^ n10862 ;
  assign n10876 = n10875 ^ n10872 ;
  assign n10877 = n10865 & n10876 ;
  assign n10878 = n10877 ^ n10874 ;
  assign n10879 = n10878 ^ n10872 ;
  assign n10880 = ~n10845 & ~n10879 ;
  assign n10881 = n10880 ^ n10845 ;
  assign n10882 = ~n10841 & ~n10881 ;
  assign n10883 = n352 & ~n10882 ;
  assign n10884 = n10883 ^ n10736 ;
  assign n10885 = n10884 ^ n10736 ;
  assign n10886 = n10885 ^ n10821 ;
  assign n10887 = n10821 & ~n10886 ;
  assign n10888 = n10887 ^ n10821 ;
  assign n10889 = ~n10822 & n10888 ;
  assign n10890 = n10889 ^ n10887 ;
  assign n10891 = n10890 ^ n10736 ;
  assign n10892 = n10891 ^ n10821 ;
  assign n10893 = x3 & n10892 ;
  assign n10894 = n10893 ^ n10736 ;
  assign n10895 = n10673 & n10894 ;
  assign n10896 = ~n10382 & ~n10895 ;
  assign n10897 = ~n263 & n10896 ;
  assign n10898 = n10381 & ~n10897 ;
  assign n10899 = n9597 & n10898 ;
  assign n10900 = ~x8 & ~n7163 ;
  assign n10901 = n2831 & n7352 ;
  assign n10902 = ~n10900 & n10901 ;
  assign n10903 = n151 & n1282 ;
  assign n10904 = n6974 & n10903 ;
  assign n10905 = n2608 ^ n124 ;
  assign n10906 = x13 & n3031 ;
  assign n10907 = n10906 ^ n2608 ;
  assign n10908 = n10907 ^ n10906 ;
  assign n10909 = n10908 ^ n10905 ;
  assign n10910 = n1407 ^ n718 ;
  assign n10911 = n1407 & n10910 ;
  assign n10912 = n10911 ^ n10906 ;
  assign n10913 = n10912 ^ n1407 ;
  assign n10914 = n10909 & ~n10913 ;
  assign n10915 = n10914 ^ n10911 ;
  assign n10916 = n10915 ^ n1407 ;
  assign n10917 = n10905 & n10916 ;
  assign n10918 = n10917 ^ n124 ;
  assign n10919 = n462 & n10918 ;
  assign n10920 = ~n10904 & ~n10919 ;
  assign n10921 = n846 & ~n4098 ;
  assign n10922 = n3230 & n5698 ;
  assign n10923 = ~n10921 & ~n10922 ;
  assign n10926 = n10923 ^ n4832 ;
  assign n10927 = n10926 ^ n10923 ;
  assign n10924 = n10923 ^ n311 ;
  assign n10925 = n10924 ^ n10923 ;
  assign n10928 = n10927 ^ n10925 ;
  assign n10929 = n10923 ^ x3 ;
  assign n10930 = n10929 ^ n10923 ;
  assign n10931 = n10930 ^ n10927 ;
  assign n10932 = n10927 & n10931 ;
  assign n10933 = n10932 ^ n10927 ;
  assign n10934 = n10928 & n10933 ;
  assign n10935 = n10934 ^ n10932 ;
  assign n10936 = n10935 ^ n10923 ;
  assign n10937 = n10936 ^ n10927 ;
  assign n10938 = ~x8 & ~n10937 ;
  assign n10939 = n10938 ^ n10923 ;
  assign n10940 = n6918 & ~n10939 ;
  assign n10941 = n328 & n3094 ;
  assign n10942 = n430 & n10941 ;
  assign n10953 = n750 & ~n1227 ;
  assign n10954 = n2959 & ~n10953 ;
  assign n10943 = n311 & n2535 ;
  assign n10944 = ~n24 & n2669 ;
  assign n10945 = ~n2608 & ~n10944 ;
  assign n10946 = ~n10943 & n10945 ;
  assign n10947 = n1117 & ~n10946 ;
  assign n10948 = ~x3 & n3031 ;
  assign n10949 = ~n1327 & n3287 ;
  assign n10950 = n366 & n10949 ;
  assign n10951 = ~n10948 & ~n10950 ;
  assign n10952 = ~n10947 & n10951 ;
  assign n10955 = n10954 ^ n10952 ;
  assign n10956 = x1 & ~n10955 ;
  assign n10957 = n10956 ^ n10954 ;
  assign n10958 = ~n10942 & ~n10957 ;
  assign n10959 = ~n10940 & n10958 ;
  assign n10960 = n10959 ^ x11 ;
  assign n10961 = n10960 ^ n10959 ;
  assign n10962 = n1282 & n2624 ;
  assign n10963 = n3187 & ~n7105 ;
  assign n10964 = ~n10962 & ~n10963 ;
  assign n10965 = n38 & ~n10964 ;
  assign n10966 = n828 & n2608 ;
  assign n10967 = ~n9748 & n10966 ;
  assign n10968 = n348 & n10967 ;
  assign n10969 = n690 & n1665 ;
  assign n10970 = n2955 & n10969 ;
  assign n10971 = ~n2624 & ~n9501 ;
  assign n10972 = n5590 & ~n10971 ;
  assign n10973 = ~n10970 & ~n10972 ;
  assign n10974 = ~n10968 & n10973 ;
  assign n10975 = ~n10965 & n10974 ;
  assign n10976 = n10975 ^ n10959 ;
  assign n10977 = ~n10961 & n10976 ;
  assign n10978 = n10977 ^ n10959 ;
  assign n10979 = n10920 & n10978 ;
  assign n10980 = ~x9 & ~n10979 ;
  assign n10981 = ~n3009 & ~n5062 ;
  assign n10982 = ~n230 & ~n10981 ;
  assign n10983 = n10982 ^ x12 ;
  assign n10984 = n10983 ^ n10982 ;
  assign n10985 = n10982 ^ n151 ;
  assign n10986 = n10985 ^ n10982 ;
  assign n10987 = ~n10984 & n10986 ;
  assign n10988 = n10987 ^ n10982 ;
  assign n10989 = x1 & n10988 ;
  assign n10990 = n10989 ^ n10982 ;
  assign n10991 = n9501 & n10990 ;
  assign n10992 = n230 & n828 ;
  assign n10993 = ~n1234 & ~n10992 ;
  assign n10994 = n2608 & ~n10993 ;
  assign n10995 = n2535 & ~n5231 ;
  assign n10996 = n730 & n10995 ;
  assign n10997 = ~n10994 & ~n10996 ;
  assign n10998 = n370 & ~n10997 ;
  assign n10999 = ~n10991 & ~n10998 ;
  assign n11000 = ~x3 & ~n10999 ;
  assign n11001 = ~x1 & n1243 ;
  assign n11002 = n106 & n2291 ;
  assign n11003 = ~n1898 & ~n11002 ;
  assign n11004 = n7664 & ~n11003 ;
  assign n11005 = ~n11001 & n11004 ;
  assign n11006 = n1226 & n5976 ;
  assign n11007 = ~n2466 & ~n3030 ;
  assign n11008 = n605 & n11007 ;
  assign n11009 = ~n5062 & ~n11008 ;
  assign n11010 = ~x1 & ~n11009 ;
  assign n11011 = ~n1247 & ~n11010 ;
  assign n11012 = ~n11006 & n11011 ;
  assign n11013 = n3187 & ~n11012 ;
  assign n11014 = n492 & n11013 ;
  assign n11015 = ~n11005 & ~n11014 ;
  assign n11016 = ~n11000 & n11015 ;
  assign n11017 = ~n10980 & n11016 ;
  assign n11018 = n11017 ^ x2 ;
  assign n11019 = n11018 ^ n11017 ;
  assign n11020 = n11019 ^ n10902 ;
  assign n11021 = ~n1169 & ~n1565 ;
  assign n11022 = n10992 & ~n11021 ;
  assign n11023 = ~n442 & n11022 ;
  assign n11024 = x1 & ~n5141 ;
  assign n11025 = n206 & n1270 ;
  assign n11026 = ~n1117 & ~n11025 ;
  assign n11027 = ~n11024 & n11026 ;
  assign n11028 = n2154 & ~n11027 ;
  assign n11029 = n442 & n1605 ;
  assign n11030 = ~x1 & n4794 ;
  assign n11031 = ~n11029 & ~n11030 ;
  assign n11032 = ~n11028 & n11031 ;
  assign n11033 = n105 & ~n11032 ;
  assign n11034 = n4612 & ~n5537 ;
  assign n11035 = n462 & n1440 ;
  assign n11036 = ~n530 & ~n633 ;
  assign n11037 = ~n870 & n11036 ;
  assign n11038 = n11035 & ~n11037 ;
  assign n11039 = ~n11034 & ~n11038 ;
  assign n11040 = x12 & ~n11039 ;
  assign n11041 = ~n11033 & ~n11040 ;
  assign n11042 = ~n11023 & n11041 ;
  assign n11043 = n11042 ^ n2608 ;
  assign n11044 = n2608 & ~n11043 ;
  assign n11045 = n11044 ^ n11017 ;
  assign n11046 = n11045 ^ n2608 ;
  assign n11047 = n11020 & ~n11046 ;
  assign n11048 = n11047 ^ n11044 ;
  assign n11049 = n11048 ^ n2608 ;
  assign n11050 = ~n10902 & n11049 ;
  assign n11051 = n11050 ^ n10902 ;
  assign n11052 = n489 & n11051 ;
  assign n11053 = n2785 & n8822 ;
  assign n11054 = n1514 & n2608 ;
  assign n11055 = n6039 & n11054 ;
  assign n11056 = ~n11053 & ~n11055 ;
  assign n11057 = n462 & ~n11056 ;
  assign n11058 = n7631 & n8822 ;
  assign n11059 = n11058 ^ x13 ;
  assign n11060 = n11059 ^ n11058 ;
  assign n11061 = n11058 ^ n11054 ;
  assign n11062 = n11061 ^ n11058 ;
  assign n11063 = ~n11060 & n11062 ;
  assign n11064 = n11063 ^ n11058 ;
  assign n11065 = ~x12 & n11064 ;
  assign n11066 = n11065 ^ n11058 ;
  assign n11067 = n5725 & n11066 ;
  assign n11068 = ~n11057 & ~n11067 ;
  assign n11069 = n175 & ~n11068 ;
  assign n11070 = n162 & n2995 ;
  assign n11071 = n1405 & n11070 ;
  assign n11072 = n1494 & n2910 ;
  assign n11073 = n4565 & n11072 ;
  assign n11074 = n3146 & n11073 ;
  assign n11075 = ~n11071 & ~n11074 ;
  assign n11076 = ~n11069 & n11075 ;
  assign n11077 = x14 & ~n11076 ;
  assign n11078 = n1265 & n2466 ;
  assign n11079 = n1869 & ~n11078 ;
  assign n11080 = x8 ^ x1 ;
  assign n11081 = n284 & n11080 ;
  assign n11082 = ~n11079 & ~n11081 ;
  assign n11083 = n2608 & ~n11082 ;
  assign n11084 = ~x11 & n718 ;
  assign n11085 = n1117 & n11084 ;
  assign n11086 = n5998 & n11007 ;
  assign n11087 = ~n2527 & ~n11086 ;
  assign n11088 = n248 & ~n1440 ;
  assign n11089 = ~n11087 & n11088 ;
  assign n11090 = ~n11085 & ~n11089 ;
  assign n11091 = ~n6528 & n11090 ;
  assign n11092 = n1169 & ~n11091 ;
  assign n11093 = n124 & n10087 ;
  assign n11094 = n456 & n623 ;
  assign n11095 = n230 & n1353 ;
  assign n11096 = ~n11094 & ~n11095 ;
  assign n11097 = ~n200 & n11096 ;
  assign n11098 = n55 & ~n11097 ;
  assign n11099 = ~n2436 & ~n11098 ;
  assign n11100 = n1364 & ~n11099 ;
  assign n11101 = ~n11093 & ~n11100 ;
  assign n11102 = n395 & n1356 ;
  assign n11103 = n442 & n2527 ;
  assign n11104 = ~n718 & n7595 ;
  assign n11105 = n11103 & ~n11104 ;
  assign n11106 = n11105 ^ x9 ;
  assign n11107 = n11106 ^ n11105 ;
  assign n11108 = n11107 ^ n11102 ;
  assign n11109 = n1117 & ~n1243 ;
  assign n11110 = ~x12 & ~n4087 ;
  assign n11111 = x8 & n6020 ;
  assign n11112 = ~n11110 & n11111 ;
  assign n11113 = ~n11109 & ~n11112 ;
  assign n11114 = n11113 ^ x1 ;
  assign n11115 = ~n11113 & ~n11114 ;
  assign n11116 = n11115 ^ n11105 ;
  assign n11117 = n11116 ^ n11113 ;
  assign n11118 = n11108 & ~n11117 ;
  assign n11119 = n11118 ^ n11115 ;
  assign n11120 = n11119 ^ n11113 ;
  assign n11121 = ~n11102 & ~n11120 ;
  assign n11122 = n11121 ^ n11102 ;
  assign n11123 = n11101 & ~n11122 ;
  assign n11124 = ~n11092 & n11123 ;
  assign n11125 = n2535 & ~n11124 ;
  assign n11126 = ~n11083 & ~n11125 ;
  assign n11127 = x2 & ~n11126 ;
  assign n11128 = x6 & n1841 ;
  assign n11129 = ~n151 & n3031 ;
  assign n11130 = ~n10966 & ~n11129 ;
  assign n11131 = ~n11128 & n11130 ;
  assign n11132 = n2083 & ~n11131 ;
  assign n11133 = ~n151 & ~n1353 ;
  assign n11134 = ~x12 & n3808 ;
  assign n11135 = ~n11133 & n11134 ;
  assign n11136 = n633 & n2669 ;
  assign n11137 = n1605 & n2535 ;
  assign n11138 = ~n1704 & n2624 ;
  assign n11139 = ~n11137 & ~n11138 ;
  assign n11140 = n76 & ~n11139 ;
  assign n11141 = ~n11136 & ~n11140 ;
  assign n11142 = ~n11135 & n11141 ;
  assign n11143 = n348 & ~n11142 ;
  assign n11144 = n263 & n2535 ;
  assign n11145 = n7201 & n11144 ;
  assign n11146 = n55 & n11145 ;
  assign n11147 = n2374 & n11072 ;
  assign n11148 = n263 & ~n1327 ;
  assign n11149 = n38 & n2608 ;
  assign n11150 = n11148 & n11149 ;
  assign n11151 = ~n11147 & ~n11150 ;
  assign n11152 = n270 & n10962 ;
  assign n11153 = n11151 & ~n11152 ;
  assign n11154 = ~n11146 & n11153 ;
  assign n11155 = n76 & n206 ;
  assign n11156 = ~n1287 & ~n11155 ;
  assign n11157 = n10921 & ~n11156 ;
  assign n11158 = n2535 & n11157 ;
  assign n11159 = n11154 & ~n11158 ;
  assign n11160 = ~n11143 & n11159 ;
  assign n11161 = ~n11132 & n11160 ;
  assign n11162 = n1524 & ~n11161 ;
  assign n11163 = n1807 & n7041 ;
  assign n11164 = n366 & n11163 ;
  assign n11165 = ~n11162 & ~n11164 ;
  assign n11166 = ~n11127 & n11165 ;
  assign n11167 = n371 & ~n11166 ;
  assign n11168 = ~n11077 & ~n11167 ;
  assign n11169 = n11009 & ~n11084 ;
  assign n11170 = ~x0 & ~n11169 ;
  assign n11171 = n1353 & n2810 ;
  assign n11172 = ~n11170 & ~n11171 ;
  assign n11173 = n3564 & ~n11172 ;
  assign n11174 = n2973 & ~n7481 ;
  assign n11175 = n1363 & n11174 ;
  assign n11176 = ~n11173 & ~n11175 ;
  assign n11177 = n466 & ~n11176 ;
  assign n11178 = n1423 & n3735 ;
  assign n11179 = n3295 & n11178 ;
  assign n11180 = n364 & ~n869 ;
  assign n11181 = ~n5095 & ~n11180 ;
  assign n11182 = n799 & n8838 ;
  assign n11183 = ~n11181 & n11182 ;
  assign n11184 = ~n623 & n7612 ;
  assign n11185 = n828 & n3187 ;
  assign n11186 = n2535 & n5838 ;
  assign n11187 = ~n11185 & ~n11186 ;
  assign n11188 = ~n11184 & ~n11187 ;
  assign n11189 = x11 & ~n1977 ;
  assign n11190 = n2608 & ~n11189 ;
  assign n11191 = ~n718 & ~n2036 ;
  assign n11192 = ~n1241 & n11191 ;
  assign n11193 = n2917 & ~n11192 ;
  assign n11194 = ~n11190 & ~n11193 ;
  assign n11195 = n465 & ~n11194 ;
  assign n11196 = ~n11188 & ~n11195 ;
  assign n11197 = n58 & ~n11196 ;
  assign n11198 = ~n11183 & ~n11197 ;
  assign n11199 = ~n11179 & n11198 ;
  assign n11200 = ~n11177 & n11199 ;
  assign n11201 = ~x9 & ~n11200 ;
  assign n11202 = ~n76 & ~n5698 ;
  assign n11203 = ~n2539 & ~n11202 ;
  assign n11204 = n874 & n2535 ;
  assign n11205 = ~n2466 & n11204 ;
  assign n11206 = ~n11203 & ~n11205 ;
  assign n11207 = n845 & ~n11206 ;
  assign n11208 = n4287 & n10247 ;
  assign n11209 = ~x4 & ~n4179 ;
  assign n11210 = ~n524 & n11209 ;
  assign n11211 = n2702 & ~n11210 ;
  assign n11212 = x0 & n11211 ;
  assign n11213 = ~n11208 & ~n11212 ;
  assign n11214 = ~n11207 & n11213 ;
  assign n11215 = n11214 ^ x2 ;
  assign n11216 = n11215 ^ n11214 ;
  assign n11217 = n1242 & n7103 ;
  assign n11218 = n11217 ^ n11214 ;
  assign n11219 = ~n11216 & ~n11218 ;
  assign n11220 = n11219 ^ n11214 ;
  assign n11221 = n263 & ~n11220 ;
  assign n11222 = ~n11201 & ~n11221 ;
  assign n11223 = n4333 & ~n11222 ;
  assign n11224 = ~n395 & n11128 ;
  assign n11225 = n56 & n58 ;
  assign n11226 = n11224 & n11225 ;
  assign n11227 = ~n11223 & ~n11226 ;
  assign n11228 = n11168 & n11227 ;
  assign n11311 = n798 & ~n4672 ;
  assign n11312 = n11311 ^ n6418 ;
  assign n11313 = n11312 ^ x2 ;
  assign n11314 = n11313 ^ n11312 ;
  assign n11315 = n11312 ^ n266 ;
  assign n11316 = n11315 ^ n6418 ;
  assign n11317 = ~n11314 & ~n11316 ;
  assign n11318 = n11317 ^ n266 ;
  assign n11319 = ~n266 & ~n275 ;
  assign n11320 = n11319 ^ n6418 ;
  assign n11321 = ~n11318 & ~n11320 ;
  assign n11322 = n11321 ^ n11319 ;
  assign n11323 = ~n6418 & n11322 ;
  assign n11324 = n11323 ^ n11317 ;
  assign n11325 = n11324 ^ x0 ;
  assign n11326 = n11325 ^ n266 ;
  assign n11327 = n127 & n11326 ;
  assign n11328 = n176 & n5180 ;
  assign n11329 = n442 & n11328 ;
  assign n11330 = ~n11327 & ~n11329 ;
  assign n11331 = n3031 & ~n11330 ;
  assign n11332 = ~x12 & ~n74 ;
  assign n11333 = ~n1038 & n11332 ;
  assign n11334 = ~n596 & n11333 ;
  assign n11335 = ~n3305 & n11334 ;
  assign n11336 = n1954 & n5175 ;
  assign n11337 = ~n11335 & ~n11336 ;
  assign n11338 = n2831 & ~n11337 ;
  assign n11339 = ~n1377 & ~n10739 ;
  assign n11340 = n11339 ^ x2 ;
  assign n11341 = n11340 ^ n11339 ;
  assign n11342 = n11339 ^ x1 ;
  assign n11343 = n11342 ^ n11339 ;
  assign n11344 = n11341 & ~n11343 ;
  assign n11345 = n11344 ^ n11339 ;
  assign n11346 = x13 & ~n11345 ;
  assign n11347 = n11346 ^ n11339 ;
  assign n11348 = n2358 & ~n11347 ;
  assign n11349 = ~n74 & ~n10573 ;
  assign n11350 = n1667 & ~n11349 ;
  assign n11351 = ~n1741 & ~n11350 ;
  assign n11352 = ~n11348 & n11351 ;
  assign n11353 = n265 & ~n11352 ;
  assign n11354 = n263 & n964 ;
  assign n11355 = n1743 & n11354 ;
  assign n11356 = ~n11353 & ~n11355 ;
  assign n11357 = n2608 & ~n11356 ;
  assign n11358 = x4 & n2686 ;
  assign n11359 = n9980 & n11358 ;
  assign n11360 = ~n1095 & ~n5231 ;
  assign n11361 = n11359 & n11360 ;
  assign n11362 = n11185 ^ x2 ;
  assign n11363 = n11362 ^ n11185 ;
  assign n11364 = n11363 ^ n11361 ;
  assign n11365 = n3569 ^ x9 ;
  assign n11366 = ~x9 & ~n11365 ;
  assign n11367 = n11366 ^ n11185 ;
  assign n11368 = n11367 ^ x9 ;
  assign n11369 = n11364 & ~n11368 ;
  assign n11370 = n11369 ^ n11366 ;
  assign n11371 = n11370 ^ x9 ;
  assign n11372 = ~n11361 & ~n11371 ;
  assign n11373 = n11372 ^ n11361 ;
  assign n11374 = n261 & n11373 ;
  assign n11375 = n1476 & n2910 ;
  assign n11376 = ~n3428 & ~n11375 ;
  assign n11377 = n4751 & ~n11376 ;
  assign n11378 = ~n11374 & ~n11377 ;
  assign n11379 = ~x3 & ~n11378 ;
  assign n11380 = n1742 & n2911 ;
  assign n11381 = n1382 & n11375 ;
  assign n11382 = n2182 & n3186 ;
  assign n11383 = n8341 & n11382 ;
  assign n11384 = ~n11381 & ~n11383 ;
  assign n11385 = ~x3 & ~n11384 ;
  assign n11386 = n55 & ~n3305 ;
  assign n11387 = ~x2 & ~n3094 ;
  assign n11388 = ~n3327 & ~n11387 ;
  assign n11389 = n11386 & n11388 ;
  assign n11390 = ~n11385 & ~n11389 ;
  assign n11391 = ~n11380 & n11390 ;
  assign n11392 = n530 & ~n11391 ;
  assign n11393 = n3295 & n6195 ;
  assign n11394 = n1756 & n11393 ;
  assign n11395 = n1275 & n2535 ;
  assign n11396 = n2608 & n5025 ;
  assign n11397 = ~n11395 & ~n11396 ;
  assign n11398 = ~n11137 & n11397 ;
  assign n11399 = ~n70 & ~n11398 ;
  assign n11400 = ~n1685 & ~n1686 ;
  assign n11401 = n1581 & n5013 ;
  assign n11402 = ~n11400 & n11401 ;
  assign n11403 = n2850 & n11402 ;
  assign n11404 = ~n11399 & ~n11403 ;
  assign n11405 = ~n11394 & n11404 ;
  assign n11406 = ~n11392 & n11405 ;
  assign n11407 = x15 & ~n11406 ;
  assign n11408 = ~n11379 & ~n11407 ;
  assign n11409 = ~n11357 & n11408 ;
  assign n11410 = ~n11338 & n11409 ;
  assign n11411 = n623 & ~n11410 ;
  assign n11412 = ~n11331 & ~n11411 ;
  assign n11413 = n2374 & n11054 ;
  assign n11414 = ~n4881 & n6436 ;
  assign n11415 = ~x12 & n123 ;
  assign n11416 = ~n11414 & ~n11415 ;
  assign n11417 = n2535 & ~n11416 ;
  assign n11418 = n7431 & n10142 ;
  assign n11419 = ~n11417 & ~n11418 ;
  assign n11420 = n370 & ~n11419 ;
  assign n11421 = n1282 ^ x9 ;
  assign n11422 = n11421 ^ n1282 ;
  assign n11423 = n11191 ^ n1282 ;
  assign n11424 = n11422 & ~n11423 ;
  assign n11425 = n11424 ^ n1282 ;
  assign n11426 = n2535 & n11425 ;
  assign n11427 = ~n11358 & ~n11426 ;
  assign n11428 = n5929 & ~n11427 ;
  assign n11429 = ~n3031 & ~n10966 ;
  assign n11430 = n284 & ~n11429 ;
  assign n11431 = n718 & n2831 ;
  assign n11432 = n1364 & n11431 ;
  assign n11433 = ~n11430 & ~n11432 ;
  assign n11434 = n74 & ~n11433 ;
  assign n11435 = ~n11428 & ~n11434 ;
  assign n11436 = ~n11420 & n11435 ;
  assign n11437 = ~n11413 & n11436 ;
  assign n11438 = n1217 & ~n11437 ;
  assign n11439 = n284 & n2754 ;
  assign n11440 = n3530 & n11439 ;
  assign n11441 = n141 & n11440 ;
  assign n11442 = ~n1382 & ~n2608 ;
  assign n11443 = ~n1349 & ~n2535 ;
  assign n11444 = n6562 & ~n11443 ;
  assign n11445 = ~n11442 & n11444 ;
  assign n11446 = n178 & n2668 ;
  assign n11447 = n6484 & n11446 ;
  assign n11448 = ~n11445 & ~n11447 ;
  assign n11449 = n579 & ~n11448 ;
  assign n11450 = n442 & n530 ;
  assign n11451 = ~x13 & n5193 ;
  assign n11452 = ~n11450 & ~n11451 ;
  assign n11453 = n3287 & n8863 ;
  assign n11454 = n11453 ^ x0 ;
  assign n11455 = n11454 ^ n11453 ;
  assign n11456 = n11453 ^ n3566 ;
  assign n11457 = n11456 ^ n11453 ;
  assign n11458 = n11455 & ~n11457 ;
  assign n11459 = n11458 ^ n11453 ;
  assign n11460 = x12 & n11459 ;
  assign n11461 = n11460 ^ n11453 ;
  assign n11462 = ~n11452 & n11461 ;
  assign n11463 = ~n11449 & ~n11462 ;
  assign n11464 = ~n11441 & n11463 ;
  assign n11465 = n1270 & ~n11464 ;
  assign n11466 = n3094 & ~n11036 ;
  assign n11467 = n2535 & n5759 ;
  assign n11468 = ~n11466 & ~n11467 ;
  assign n11469 = n38 & ~n11468 ;
  assign n11470 = n396 & ~n673 ;
  assign n11471 = ~n2326 & n11470 ;
  assign n11472 = ~n9860 & ~n11471 ;
  assign n11473 = n3094 & ~n11472 ;
  assign n11474 = n6993 & n9501 ;
  assign n11475 = ~n11473 & ~n11474 ;
  assign n11476 = ~n11469 & n11475 ;
  assign n11477 = n2608 ^ x9 ;
  assign n11478 = n11477 ^ n348 ;
  assign n11479 = n10944 ^ n6021 ;
  assign n11480 = x9 & ~n11479 ;
  assign n11481 = n11480 ^ n6021 ;
  assign n11482 = n11478 & n11481 ;
  assign n11483 = n11482 ^ n11480 ;
  assign n11484 = n11483 ^ n6021 ;
  assign n11485 = n11484 ^ x9 ;
  assign n11486 = n348 & n11485 ;
  assign n11487 = n11476 & ~n11486 ;
  assign n11488 = n988 & ~n11487 ;
  assign n11489 = ~n11465 & ~n11488 ;
  assign n11490 = n282 & n333 ;
  assign n11491 = n3031 & n11490 ;
  assign n11492 = n2083 & ~n11191 ;
  assign n11493 = x9 & n55 ;
  assign n11494 = ~n7481 & n11493 ;
  assign n11495 = ~n11492 & ~n11494 ;
  assign n11496 = n9157 & ~n11495 ;
  assign n11497 = ~x2 & n11496 ;
  assign n11498 = ~n11491 & ~n11497 ;
  assign n11499 = ~n5143 & ~n9024 ;
  assign n11500 = ~n3566 & ~n11499 ;
  assign n11501 = ~n4672 & n11500 ;
  assign n11502 = n310 & n3569 ;
  assign n11503 = n175 & n3295 ;
  assign n11504 = ~n19 & n11503 ;
  assign n11505 = ~n11502 & ~n11504 ;
  assign n11506 = n6986 & ~n11505 ;
  assign n11507 = n57 & n2538 ;
  assign n11508 = n306 & n2535 ;
  assign n11509 = ~n8952 & n11508 ;
  assign n11510 = ~n11507 & ~n11509 ;
  assign n11511 = ~n267 & ~n11510 ;
  assign n11512 = n263 & n11446 ;
  assign n11513 = n1756 & n6916 ;
  assign n11514 = ~n11512 & ~n11513 ;
  assign n11515 = n262 & n874 ;
  assign n11516 = n45 & n65 ;
  assign n11517 = ~n11515 & ~n11516 ;
  assign n11518 = ~n11514 & ~n11517 ;
  assign n11519 = ~n11511 & ~n11518 ;
  assign n11520 = ~n11506 & n11519 ;
  assign n11521 = ~n11501 & n11520 ;
  assign n11522 = n311 & ~n11521 ;
  assign n11523 = n11498 & ~n11522 ;
  assign n11524 = n11489 & n11523 ;
  assign n11525 = ~n11438 & n11524 ;
  assign n11526 = n11525 ^ n2608 ;
  assign n11527 = n11526 ^ x11 ;
  assign n11569 = n11527 ^ n11526 ;
  assign n11528 = ~n1146 & n2083 ;
  assign n11529 = n492 & n11332 ;
  assign n11530 = ~n11528 & ~n11529 ;
  assign n11531 = n718 & ~n11530 ;
  assign n11532 = n404 & ~n1665 ;
  assign n11533 = n205 & n11532 ;
  assign n11534 = n5721 & n9925 ;
  assign n11535 = n332 & n1665 ;
  assign n11536 = ~n1038 & n11535 ;
  assign n11537 = ~n11534 & ~n11536 ;
  assign n11538 = ~n757 & n6099 ;
  assign n11539 = ~n1317 & n11538 ;
  assign n11540 = n11537 & ~n11539 ;
  assign n11541 = ~n11533 & n11540 ;
  assign n11542 = ~n11531 & n11541 ;
  assign n11543 = x0 & ~n11542 ;
  assign n11544 = n123 & n6958 ;
  assign n11545 = n1263 & ~n9926 ;
  assign n11546 = n5193 & ~n8952 ;
  assign n11547 = ~n11450 & ~n11546 ;
  assign n11548 = ~n741 & ~n11547 ;
  assign n11549 = ~n11545 & ~n11548 ;
  assign n11550 = x14 & ~n11549 ;
  assign n11551 = ~n11544 & ~n11550 ;
  assign n11552 = ~n11543 & n11551 ;
  assign n11553 = n406 & ~n11552 ;
  assign n11554 = n1251 & n6574 ;
  assign n11555 = ~n1704 & n5512 ;
  assign n11556 = n492 & n7277 ;
  assign n11557 = ~n11555 & ~n11556 ;
  assign n11558 = ~n5193 & n11557 ;
  assign n11559 = n2913 & ~n11558 ;
  assign n11560 = ~x8 & n11559 ;
  assign n11561 = ~n11554 & ~n11560 ;
  assign n11562 = ~n11553 & n11561 ;
  assign n11563 = n11562 ^ n11527 ;
  assign n11564 = n11563 ^ n11526 ;
  assign n11565 = n11527 ^ n11525 ;
  assign n11566 = n11565 ^ n11562 ;
  assign n11567 = n11566 ^ n11564 ;
  assign n11568 = ~n11564 & ~n11567 ;
  assign n11570 = n11569 ^ n11568 ;
  assign n11571 = n11570 ^ n11564 ;
  assign n11572 = n74 & n7783 ;
  assign n11573 = x8 & n11572 ;
  assign n11574 = n333 & n11148 ;
  assign n11575 = n264 & n306 ;
  assign n11576 = ~n11574 & ~n11575 ;
  assign n11577 = ~n1627 & n9677 ;
  assign n11578 = n1374 & n11577 ;
  assign n11579 = n1275 & ~n9623 ;
  assign n11580 = ~n11578 & ~n11579 ;
  assign n11581 = n11576 & n11580 ;
  assign n11582 = ~n11573 & n11581 ;
  assign n11583 = n11582 ^ n11526 ;
  assign n11584 = n11568 ^ n11564 ;
  assign n11585 = ~n11583 & ~n11584 ;
  assign n11586 = n11585 ^ n11526 ;
  assign n11587 = n11571 & ~n11586 ;
  assign n11588 = n11587 ^ n11526 ;
  assign n11589 = n11588 ^ n2608 ;
  assign n11590 = n11589 ^ n11526 ;
  assign n11591 = n11412 & ~n11590 ;
  assign n11229 = x3 & n2535 ;
  assign n11230 = n10903 & n11229 ;
  assign n11231 = n846 & n3687 ;
  assign n11232 = ~n11230 & ~n11231 ;
  assign n11233 = ~n370 & ~n11232 ;
  assign n11234 = n1263 & n1353 ;
  assign n11235 = ~n1977 & ~n11234 ;
  assign n11236 = n3002 & ~n11235 ;
  assign n11237 = x3 & ~n1327 ;
  assign n11238 = n3808 & n11237 ;
  assign n11239 = ~n11236 & ~n11238 ;
  assign n11240 = n214 & ~n11239 ;
  assign n11241 = n7806 & n10943 ;
  assign n11242 = n370 & n10943 ;
  assign n11243 = ~n633 & ~n1270 ;
  assign n11244 = n7393 & ~n11243 ;
  assign n11245 = ~n1038 & n11244 ;
  assign n11246 = ~n11242 & ~n11245 ;
  assign n11247 = n2608 ^ x13 ;
  assign n11248 = n11247 ^ n396 ;
  assign n11249 = n10943 ^ x14 ;
  assign n11250 = x13 & ~n11249 ;
  assign n11251 = n11250 ^ x14 ;
  assign n11252 = n11248 & n11251 ;
  assign n11253 = n11252 ^ n11250 ;
  assign n11254 = n11253 ^ x14 ;
  assign n11255 = n11254 ^ x13 ;
  assign n11256 = n396 & n11255 ;
  assign n11257 = n11246 & ~n11256 ;
  assign n11258 = ~x12 & ~n11257 ;
  assign n11259 = ~n11241 & ~n11258 ;
  assign n11260 = n162 & ~n11259 ;
  assign n11261 = n650 & n1627 ;
  assign n11262 = n11144 & n11261 ;
  assign n11263 = ~n311 & ~n2154 ;
  assign n11264 = ~n24 & ~n370 ;
  assign n11265 = ~n11263 & n11264 ;
  assign n11266 = ~x6 & n11265 ;
  assign n11267 = ~x4 & ~n11266 ;
  assign n11268 = n1117 & ~n2575 ;
  assign n11269 = ~n1364 & n11268 ;
  assign n11270 = ~n19 & n11269 ;
  assign n11271 = ~n1169 & n11270 ;
  assign n11272 = ~n11267 & n11271 ;
  assign n11273 = n7023 & n9817 ;
  assign n11274 = ~n11272 & ~n11273 ;
  assign n11275 = ~n11262 & n11274 ;
  assign n11276 = ~n11260 & n11275 ;
  assign n11277 = ~n11240 & n11276 ;
  assign n11278 = x11 & ~n11277 ;
  assign n11279 = ~n11233 & ~n11278 ;
  assign n11280 = n20 & ~n11279 ;
  assign n11281 = ~n2824 & ~n5129 ;
  assign n11282 = n11054 & ~n11281 ;
  assign n11283 = ~n11053 & ~n11282 ;
  assign n11284 = n1264 & ~n11283 ;
  assign n11285 = n690 & n11284 ;
  assign n11286 = ~n11280 & ~n11285 ;
  assign n11287 = n1214 & n5013 ;
  assign n11288 = x12 ^ x1 ;
  assign n11289 = n11288 ^ x12 ;
  assign n11290 = n4832 ^ x12 ;
  assign n11291 = ~n11289 & ~n11290 ;
  assign n11292 = n11291 ^ x12 ;
  assign n11293 = n275 & ~n11292 ;
  assign n11294 = ~n11287 & ~n11293 ;
  assign n11295 = n6992 & ~n11294 ;
  assign n11296 = n1869 & n4656 ;
  assign n11297 = ~n11029 & ~n11296 ;
  assign n11298 = ~x13 & ~n11297 ;
  assign n11299 = n56 & n5129 ;
  assign n11300 = n265 & n11299 ;
  assign n11301 = ~n9830 & ~n11024 ;
  assign n11302 = n870 & ~n1665 ;
  assign n11303 = ~n11301 & n11302 ;
  assign n11304 = ~n11300 & ~n11303 ;
  assign n11305 = ~n11298 & n11304 ;
  assign n11306 = n2608 & ~n11305 ;
  assign n11307 = ~n11295 & ~n11306 ;
  assign n11308 = n623 & ~n11307 ;
  assign n11309 = n928 & n11308 ;
  assign n11310 = n11286 & ~n11309 ;
  assign n11592 = n11591 ^ n11310 ;
  assign n11593 = x10 & n11592 ;
  assign n11594 = n11593 ^ n11591 ;
  assign n11595 = n11228 & n11594 ;
  assign n11596 = ~n11052 & n11595 ;
  assign n11597 = ~n2902 & ~n11596 ;
  assign n11598 = n10899 & ~n11597 ;
  assign n11599 = ~n7980 & n11598 ;
  assign n11600 = ~n6904 & n11599 ;
  assign n11601 = n5784 & n11600 ;
  assign y0 = ~n11601 ;
endmodule
