module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 ;
  output y0 ;
  wire n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 ;
  assign n31 = ~x6 & ~x7 ;
  assign n32 = ~x22 & ~x23 ;
  assign n33 = ~x28 & ~x29 ;
  assign n34 = ~x27 & ~n33 ;
  assign n35 = ~x26 & ~n34 ;
  assign n36 = ~x24 & ~x25 ;
  assign n37 = ~n35 & n36 ;
  assign n38 = n32 & ~n37 ;
  assign n39 = ~x20 & ~x21 ;
  assign n40 = ~n38 & n39 ;
  assign n41 = ~x19 & ~n40 ;
  assign n42 = ~x18 & ~n41 ;
  assign n43 = ~x16 & ~x17 ;
  assign n44 = ~n42 & n43 ;
  assign n45 = ~x15 & ~n44 ;
  assign n46 = ~x14 & ~n45 ;
  assign n47 = ~x12 & ~x13 ;
  assign n48 = ~n46 & n47 ;
  assign n49 = ~x11 & ~n48 ;
  assign n50 = ~x10 & ~n49 ;
  assign n51 = ~x8 & ~x9 ;
  assign n52 = ~n50 & n51 ;
  assign n53 = n31 & ~n52 ;
  assign n54 = ~x4 & ~x5 ;
  assign n55 = ~n53 & n54 ;
  assign n56 = ~x3 & ~n55 ;
  assign n57 = ~x2 & ~n56 ;
  assign n58 = ~x0 & ~n57 ;
  assign n59 = ~x1 & n58 ;
  assign y0 = ~n59 ;
endmodule
