// Benchmark "./pla/exam.pla_dbb_orig_8NonExact" written by ABC on Fri Nov 20 10:21:17 2020

module \./pla/exam.pla_dbb_orig_8NonExact  ( 
    x0,
    z0  );
  input  x0;
  output z0;
  assign z0 = 1'b1;
endmodule


